module fake_jpeg_26709_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_18;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_22),
.A2(n_1),
.B(n_2),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_25),
.Y(n_50)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_50),
.B1(n_36),
.B2(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_15),
.B1(n_21),
.B2(n_27),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_15),
.B1(n_21),
.B2(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_51),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_57),
.A2(n_72),
.B1(n_69),
.B2(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_71),
.B1(n_75),
.B2(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_61),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_32),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_32),
.C(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_36),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_77),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_40),
.A2(n_37),
.B1(n_39),
.B2(n_20),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_46),
.A2(n_16),
.B1(n_30),
.B2(n_17),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_74),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_44),
.A2(n_37),
.B1(n_39),
.B2(n_53),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_39),
.B1(n_20),
.B2(n_16),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g79 ( 
.A(n_46),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_20),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_17),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_55),
.Y(n_128)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_87),
.B(n_90),
.Y(n_116)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_54),
.B1(n_22),
.B2(n_32),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_95),
.B1(n_57),
.B2(n_77),
.Y(n_113)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_100),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_32),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_61),
.B(n_30),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_105),
.B(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_59),
.B1(n_65),
.B2(n_67),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_129),
.B1(n_114),
.B2(n_128),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_108),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_114),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_71),
.B1(n_64),
.B2(n_75),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_118),
.B1(n_83),
.B2(n_96),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_92),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_128),
.B1(n_98),
.B2(n_25),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_64),
.B1(n_78),
.B2(n_76),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_85),
.B(n_62),
.C(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_130),
.B(n_91),
.Y(n_146)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_32),
.C(n_60),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_123),
.C(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_55),
.C(n_81),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_29),
.Y(n_127)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_69),
.B1(n_73),
.B2(n_20),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_25),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_25),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_92),
.B1(n_99),
.B2(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_137),
.B1(n_140),
.B2(n_148),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_147),
.B1(n_155),
.B2(n_118),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_112),
.A2(n_87),
.B1(n_90),
.B2(n_88),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_84),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_88),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_150),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_125),
.B(n_117),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_150),
.B(n_10),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_91),
.B1(n_83),
.B2(n_82),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_82),
.B1(n_106),
.B2(n_98),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_151),
.B1(n_158),
.B2(n_18),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_89),
.B(n_19),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_98),
.B1(n_31),
.B2(n_29),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_19),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_25),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_156),
.C(n_123),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_111),
.A2(n_31),
.B1(n_29),
.B2(n_26),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_31),
.C(n_26),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_18),
.B1(n_19),
.B2(n_4),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_167),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_162),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_166),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_131),
.C(n_121),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_144),
.C(n_154),
.Y(n_194)
);

XNOR2x2_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_152),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_18),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_174),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_10),
.C(n_5),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_178),
.B1(n_136),
.B2(n_143),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_179),
.B(n_181),
.Y(n_191)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_143),
.Y(n_181)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_136),
.B1(n_140),
.B2(n_153),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_124),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_195),
.C(n_199),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_164),
.C(n_160),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_146),
.B(n_158),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_1),
.B(n_6),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_157),
.C(n_135),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_173),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_207),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_183),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_202),
.Y(n_218)
);

AOI322xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_159),
.A3(n_170),
.B1(n_174),
.B2(n_171),
.C1(n_166),
.C2(n_180),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_178),
.C(n_181),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_210),
.Y(n_221)
);

XNOR2x2_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_11),
.Y(n_206)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_211),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_124),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_124),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_11),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_9),
.C(n_6),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_211),
.C(n_191),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_189),
.B1(n_188),
.B2(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_190),
.B1(n_185),
.B2(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_219),
.Y(n_235)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_208),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_196),
.Y(n_231)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_218),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_233),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_221),
.B(n_207),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_212),
.C(n_223),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_231),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_191),
.B(n_206),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_224),
.B(n_222),
.Y(n_236)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_212),
.CI(n_211),
.CON(n_233),
.SN(n_233)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_234),
.B(n_6),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_223),
.C(n_219),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g239 ( 
.A1(n_233),
.A2(n_224),
.B(n_226),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_239),
.A2(n_242),
.B(n_11),
.Y(n_244)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_215),
.Y(n_242)
);

AOI322xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_1),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_224),
.C2(n_220),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_8),
.B(n_9),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_247),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_242),
.B(n_8),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_7),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_252),
.B(n_250),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_254),
.A2(n_253),
.B1(n_251),
.B2(n_14),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_12),
.Y(n_256)
);


endmodule