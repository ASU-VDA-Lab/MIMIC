module fake_jpeg_25662_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_10),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_42),
.Y(n_52)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_22),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_48),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_20),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_50),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_15),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_27),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_74),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_26),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_26),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_70),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_41),
.A2(n_29),
.B1(n_17),
.B2(n_22),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_23),
.B1(n_19),
.B2(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_28),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_29),
.B1(n_17),
.B2(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_73),
.B1(n_77),
.B2(n_18),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_29),
.B1(n_17),
.B2(n_16),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_28),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_79),
.B(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_16),
.B1(n_34),
.B2(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_34),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_86),
.A2(n_53),
.B1(n_81),
.B2(n_74),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_87),
.B(n_99),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_97),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_57),
.A2(n_33),
.B1(n_24),
.B2(n_31),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_54),
.A2(n_31),
.B(n_18),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_33),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_33),
.B1(n_24),
.B2(n_3),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_53),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_63),
.B1(n_60),
.B2(n_59),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_4),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_4),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_63),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_111),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_84),
.B1(n_101),
.B2(n_90),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_124),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_80),
.B1(n_60),
.B2(n_67),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_110),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_11),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_126),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_80),
.B1(n_63),
.B2(n_5),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_12),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_130),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_5),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_133),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_13),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_107),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_13),
.B1(n_99),
.B2(n_88),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_126),
.Y(n_157)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_104),
.Y(n_156)
);

OR2x6_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_91),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_137),
.A2(n_98),
.B(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_148),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_129),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_143),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_95),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_97),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_151),
.A2(n_153),
.B(n_155),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_137),
.A2(n_108),
.B1(n_103),
.B2(n_90),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_103),
.B(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_126),
.B(n_115),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_128),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_157),
.A2(n_116),
.A3(n_121),
.B1(n_135),
.B2(n_118),
.C1(n_134),
.C2(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_175),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_149),
.B(n_121),
.C(n_116),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_166),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_158),
.C(n_154),
.Y(n_166)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_152),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_172),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_133),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_120),
.B(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_136),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_181),
.Y(n_191)
);

AND5x1_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_157),
.C(n_150),
.D(n_159),
.E(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_183),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_150),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_176),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_184),
.Y(n_197)
);

OAI22x1_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_150),
.B1(n_146),
.B2(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_169),
.B1(n_163),
.B2(n_171),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_140),
.B1(n_148),
.B2(n_130),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_163),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_173),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_196),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_173),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_166),
.C(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_200),
.A2(n_188),
.B1(n_180),
.B2(n_181),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_203),
.B1(n_207),
.B2(n_170),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_191),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_202),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_194),
.A2(n_183),
.B1(n_195),
.B2(n_186),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_145),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_187),
.B1(n_185),
.B2(n_189),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_213),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_208),
.C(n_193),
.Y(n_216)
);

NAND4xp25_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_177),
.C(n_180),
.D(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_160),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_217),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_210),
.B(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_215),
.B(n_201),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_219),
.B(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

AOI321xp33_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_216),
.A3(n_223),
.B1(n_165),
.B2(n_204),
.C(n_212),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_204),
.Y(n_227)
);


endmodule