module fake_jpeg_19773_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_62),
.Y(n_77)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_50),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_64),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_32),
.B1(n_27),
.B2(n_41),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_70),
.B1(n_92),
.B2(n_43),
.Y(n_104)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_71),
.Y(n_110)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_18),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_32),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_79),
.B1(n_85),
.B2(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_26),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_89),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_35),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_95),
.Y(n_117)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_37),
.B1(n_40),
.B2(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_52),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_27),
.B1(n_33),
.B2(n_38),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_52),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_40),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_93),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_74),
.B1(n_84),
.B2(n_39),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_43),
.B1(n_38),
.B2(n_48),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_86),
.B1(n_70),
.B2(n_48),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_112),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_38),
.B(n_56),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_52),
.B(n_44),
.Y(n_154)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_75),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_43),
.B1(n_39),
.B2(n_36),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_123),
.B1(n_60),
.B2(n_83),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_39),
.B1(n_36),
.B2(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_88),
.Y(n_129)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_133),
.B1(n_137),
.B2(n_150),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_152),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_134),
.B1(n_141),
.B2(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_112),
.B1(n_100),
.B2(n_114),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_83),
.B1(n_36),
.B2(n_87),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_26),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_121),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_107),
.B1(n_116),
.B2(n_86),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_93),
.B1(n_90),
.B2(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_52),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_143),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_96),
.A2(n_0),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_154),
.B(n_122),
.Y(n_178)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_44),
.B1(n_42),
.B2(n_52),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_99),
.B(n_69),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_102),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_44),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_161),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_150),
.B1(n_153),
.B2(n_149),
.Y(n_189)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_176),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_106),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_101),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_187),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_116),
.C(n_101),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_80),
.C(n_44),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_106),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_168),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_173),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_154),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_110),
.B1(n_115),
.B2(n_124),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_171),
.B1(n_42),
.B2(n_20),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_127),
.B1(n_136),
.B2(n_137),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_125),
.B(n_122),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_178),
.B(n_185),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_110),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_186),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_183),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_98),
.B(n_102),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_103),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_20),
.A3(n_42),
.B1(n_44),
.B2(n_26),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_194),
.B1(n_203),
.B2(n_177),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_184),
.A2(n_138),
.B1(n_120),
.B2(n_113),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_190),
.A2(n_200),
.B1(n_185),
.B2(n_183),
.Y(n_227)
);

XNOR2x1_ASAP7_75t_L g191 ( 
.A(n_161),
.B(n_138),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_191),
.A2(n_164),
.B1(n_180),
.B2(n_178),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_195),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_163),
.A2(n_120),
.B1(n_67),
.B2(n_63),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_168),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_42),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_157),
.A2(n_29),
.B1(n_22),
.B2(n_16),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_17),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_217),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_0),
.B(n_1),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_210),
.A2(n_31),
.B(n_2),
.Y(n_241)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_213),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_103),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_80),
.B1(n_28),
.B2(n_24),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_80),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_24),
.Y(n_243)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_229),
.C(n_211),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_206),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_179),
.B1(n_172),
.B2(n_159),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_227),
.B1(n_231),
.B2(n_236),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_180),
.B1(n_171),
.B2(n_176),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_225),
.A2(n_197),
.B1(n_219),
.B2(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_155),
.C(n_165),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_187),
.B(n_2),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_233),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_198),
.A2(n_29),
.B1(n_22),
.B2(n_34),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_191),
.A2(n_31),
.B(n_30),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_200),
.A2(n_34),
.B1(n_28),
.B2(n_24),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_194),
.B1(n_196),
.B2(n_203),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_188),
.B1(n_208),
.B2(n_209),
.Y(n_254)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_196),
.A2(n_45),
.B1(n_80),
.B2(n_28),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_241),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_0),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_246),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_214),
.C(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_248),
.B(n_251),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_218),
.C(n_204),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_225),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_240),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_224),
.A2(n_212),
.B1(n_202),
.B2(n_205),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_239),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_262),
.B(n_265),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_216),
.C(n_45),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_45),
.C(n_10),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_9),
.C(n_14),
.Y(n_263)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_9),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_264),
.A2(n_241),
.B1(n_232),
.B2(n_223),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_9),
.B(n_14),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_231),
.B1(n_236),
.B2(n_235),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_275),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_230),
.B1(n_237),
.B2(n_244),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_234),
.B(n_226),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_234),
.B(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_250),
.A2(n_223),
.B1(n_240),
.B2(n_11),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_240),
.B1(n_15),
.B2(n_13),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_279),
.A2(n_263),
.B1(n_11),
.B2(n_12),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_245),
.B1(n_253),
.B2(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_295),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_286),
.A2(n_275),
.B1(n_270),
.B2(n_274),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_251),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_293),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_246),
.C(n_248),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_13),
.C(n_6),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_267),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_15),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_15),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_276),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_293),
.Y(n_306)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_12),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_268),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_280),
.C(n_279),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_12),
.B(n_11),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_306),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_287),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_297),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_309),
.A2(n_13),
.B(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_2),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_290),
.B(n_289),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_314),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_319),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_284),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_310),
.B(n_303),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_299),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_SL g324 ( 
.A(n_311),
.B(n_300),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_299),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_323),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_315),
.Y(n_327)
);

AO221x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_325),
.B1(n_314),
.B2(n_320),
.C(n_296),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_307),
.B(n_7),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_6),
.C(n_7),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_6),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_8),
.B1(n_262),
.B2(n_258),
.Y(n_334)
);


endmodule