module fake_jpeg_3756_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx11_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_7),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_21),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_1),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_3),
.C(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_18),
.B(n_5),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_23),
.B1(n_17),
.B2(n_13),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_9),
.B1(n_15),
.B2(n_12),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_13),
.B1(n_14),
.B2(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_31),
.B1(n_19),
.B2(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_9),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_14),
.B1(n_8),
.B2(n_16),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_38),
.B(n_39),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_23),
.B1(n_27),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_36),
.B1(n_37),
.B2(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_12),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_20),
.B1(n_6),
.B2(n_5),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_28),
.B(n_24),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_44),
.B(n_40),
.Y(n_47)
);

BUFx24_ASAP7_75t_SL g46 ( 
.A(n_42),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_26),
.B(n_20),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_43),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_42),
.Y(n_51)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_52),
.A3(n_36),
.B1(n_37),
.B2(n_45),
.C1(n_30),
.C2(n_6),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_46),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_52),
.B(n_30),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_30),
.Y(n_55)
);


endmodule