module fake_jpeg_27628_n_250 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_16),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_40),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_22),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_18),
.B1(n_23),
.B2(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_18),
.B1(n_21),
.B2(n_27),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_18),
.B1(n_27),
.B2(n_31),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_21),
.B1(n_33),
.B2(n_17),
.Y(n_54)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_34),
.Y(n_59)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_15),
.C(n_14),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_62),
.B(n_64),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_34),
.B1(n_31),
.B2(n_20),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_66),
.B1(n_68),
.B2(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_59),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_71),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_61),
.A2(n_20),
.B1(n_19),
.B2(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_29),
.B1(n_26),
.B2(n_24),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_36),
.B1(n_42),
.B2(n_24),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_92),
.Y(n_94)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_77),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_25),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_29),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_28),
.C(n_33),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_25),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_42),
.Y(n_81)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_88),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_24),
.B1(n_28),
.B2(n_33),
.Y(n_82)
);

NOR2x1_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_24),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_86),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_28),
.Y(n_86)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_24),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_88),
.A2(n_52),
.B1(n_55),
.B2(n_51),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_73),
.B1(n_87),
.B2(n_76),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_78),
.A2(n_0),
.B(n_1),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_1),
.B(n_2),
.Y(n_138)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_108),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_55),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_79),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_104),
.B(n_105),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_89),
.A2(n_55),
.B1(n_33),
.B2(n_17),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_144)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_65),
.B(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_116),
.B(n_117),
.Y(n_143)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_14),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_131),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_78),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_129),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_125),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_104),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_145),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_94),
.A2(n_92),
.B1(n_93),
.B2(n_90),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_137),
.B1(n_142),
.B2(n_107),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_95),
.B(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_134),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_69),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_91),
.B(n_72),
.C(n_71),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_140),
.B(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_144),
.B1(n_108),
.B2(n_101),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_97),
.A2(n_70),
.B1(n_73),
.B2(n_83),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_141),
.B(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_83),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_146),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_1),
.B(n_2),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_17),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_4),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_117),
.B1(n_100),
.B2(n_98),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_157),
.B1(n_167),
.B2(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_136),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_155),
.B1(n_159),
.B2(n_144),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_163),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_145),
.A2(n_96),
.B1(n_107),
.B2(n_8),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_121),
.A2(n_96),
.B(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_161),
.Y(n_188)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_168),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_7),
.C(n_9),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_138),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_143),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_133),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_10),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_141),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_11),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_171),
.A2(n_172),
.B1(n_177),
.B2(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_132),
.B1(n_130),
.B2(n_123),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_179),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_160),
.B(n_123),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_168),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_132),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_177),
.A2(n_159),
.B(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_180),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_135),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_132),
.B1(n_130),
.B2(n_12),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_190),
.B1(n_164),
.B2(n_158),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_12),
.B1(n_132),
.B2(n_148),
.Y(n_190)
);

OA21x2_ASAP7_75t_SL g191 ( 
.A1(n_186),
.A2(n_160),
.B(n_166),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_193),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_197),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_213)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_184),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.C(n_174),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_147),
.C(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_196),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_177),
.B1(n_190),
.B2(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_203),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g210 ( 
.A(n_200),
.B(n_147),
.CI(n_182),
.CON(n_210),
.SN(n_210)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_211),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_164),
.C(n_167),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_216),
.C(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_188),
.C(n_169),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_218),
.B(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_222),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_226),
.Y(n_234)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_202),
.C(n_201),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_185),
.B1(n_204),
.B2(n_217),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_198),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_206),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_212),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_233),
.B1(n_210),
.B2(n_225),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_170),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_215),
.B1(n_197),
.B2(n_222),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_212),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_231),
.A2(n_220),
.B(n_216),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_238),
.B(n_239),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_237),
.B(n_240),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_210),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_240),
.A2(n_234),
.B1(n_225),
.B2(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_244),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_245),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_243),
.C(n_211),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_228),
.Y(n_250)
);


endmodule