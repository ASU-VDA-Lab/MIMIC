module fake_jpeg_16387_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx12_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_27),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_18),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_2),
.B(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_1),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_9),
.B(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_15),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_30),
.B(n_41),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_20),
.A2(n_12),
.B1(n_17),
.B2(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_12),
.B1(n_21),
.B2(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_10),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_43),
.A2(n_44),
.B1(n_51),
.B2(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_26),
.B1(n_14),
.B2(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_49),
.A2(n_33),
.B1(n_31),
.B2(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_14),
.B1(n_24),
.B2(n_7),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_35),
.C(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_42),
.Y(n_59)
);

AO22x1_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_45),
.B1(n_43),
.B2(n_51),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_54),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_58),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_62),
.Y(n_65)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

AO221x1_ASAP7_75t_L g66 ( 
.A1(n_61),
.A2(n_64),
.B1(n_46),
.B2(n_48),
.C(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_47),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_58),
.C(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_68),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_67),
.B(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.C(n_69),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_65),
.C(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_53),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_57),
.Y(n_75)
);


endmodule