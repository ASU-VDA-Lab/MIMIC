module fake_netlist_6_4893_n_1785 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1785);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1785;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_71),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_53),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_43),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_117),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_0),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_26),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_7),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_40),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_23),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_10),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_25),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_37),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_6),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_54),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_41),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_87),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_140),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_86),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_63),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_51),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_60),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_68),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_15),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_75),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_31),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_130),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_21),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_70),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_2),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_94),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_156),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_72),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_77),
.Y(n_217)
);

BUFx8_ASAP7_75t_SL g218 ( 
.A(n_149),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_18),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_93),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_42),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_139),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_74),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_30),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_107),
.Y(n_229)
);

BUFx8_ASAP7_75t_SL g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_62),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_80),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_79),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_106),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_105),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_114),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_122),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_151),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_43),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_50),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_59),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_99),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_119),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_143),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_46),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_58),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_108),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_85),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_88),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_39),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_49),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_12),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_103),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_16),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_44),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_33),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_154),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_25),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_23),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_100),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_89),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_135),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_116),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_50),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_112),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_133),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_155),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_55),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_37),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_91),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_73),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_64),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_27),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_47),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_66),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_96),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_57),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_32),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_41),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_138),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_46),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_128),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_8),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_160),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_52),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_78),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_141),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_49),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_36),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_81),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_113),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_158),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_5),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_126),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_162),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_134),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_10),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_28),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_33),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_164),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_27),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_101),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_24),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_38),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_31),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_61),
.Y(n_320)
);

BUFx10_ASAP7_75t_L g321 ( 
.A(n_51),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_32),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_13),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_137),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_157),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_123),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_47),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_84),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_40),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_4),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_97),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_21),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_18),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_44),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_29),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_13),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_3),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_163),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_102),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_292),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_262),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_218),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_192),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_195),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_274),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_226),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_230),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_337),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_247),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_247),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_292),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_206),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

BUFx6f_ASAP7_75t_SL g362 ( 
.A(n_208),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_259),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_256),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_259),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_223),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_214),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_259),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_259),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_211),
.Y(n_370)
);

INVxp33_ASAP7_75t_L g371 ( 
.A(n_196),
.Y(n_371)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_256),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_259),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_266),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_266),
.Y(n_375)
);

INVx4_ASAP7_75t_R g376 ( 
.A(n_282),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_216),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_217),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_220),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_266),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_266),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_266),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_176),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_176),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_221),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_222),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_250),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_173),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_321),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_282),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_250),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_231),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_201),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_232),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_173),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_227),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_227),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_207),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_237),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_209),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_240),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_293),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_219),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_224),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_244),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_258),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_208),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_293),
.Y(n_412)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_264),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_281),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_208),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_177),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_287),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_245),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_295),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_171),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_297),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_246),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_248),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_177),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_299),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_307),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_311),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_175),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_341),
.A2(n_346),
.B(n_343),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_365),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_354),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_360),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_395),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g438 ( 
.A(n_424),
.Y(n_438)
);

NAND2x1p5_ASAP7_75t_L g439 ( 
.A(n_341),
.B(n_187),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_359),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_187),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_365),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_169),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_370),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_395),
.B(n_201),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g452 ( 
.A(n_411),
.B(n_236),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_377),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_343),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_406),
.Y(n_456)
);

OA21x2_ASAP7_75t_L g457 ( 
.A1(n_346),
.A2(n_323),
.B(n_319),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_353),
.B(n_236),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_350),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_356),
.B(n_169),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_350),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_372),
.B(n_390),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_357),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_342),
.A2(n_178),
.B1(n_257),
.B2(n_205),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_373),
.B(n_242),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_357),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_172),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_374),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_R g476 ( 
.A(n_344),
.B(n_249),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_380),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_385),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_358),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_402),
.B(n_313),
.C(n_203),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_381),
.B(n_172),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_406),
.B(n_242),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_358),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_411),
.A2(n_312),
.B1(n_317),
.B2(n_243),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_383),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_349),
.B(n_252),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_384),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_347),
.A2(n_198),
.B1(n_188),
.B2(n_338),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_424),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_364),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_364),
.B(n_284),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_355),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_400),
.B(n_174),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_409),
.B(n_284),
.Y(n_503)
);

BUFx8_ASAP7_75t_L g504 ( 
.A(n_362),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_422),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_441),
.A2(n_348),
.B1(n_313),
.B2(n_398),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_441),
.A2(n_458),
.B1(n_431),
.B2(n_457),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_455),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_455),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_462),
.B(n_416),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_461),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_461),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_462),
.B(n_378),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_458),
.B(n_400),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_465),
.B(n_451),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_470),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_470),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_435),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_452),
.B(n_415),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_461),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_496),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_451),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_470),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_463),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_451),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_441),
.A2(n_333),
.B1(n_324),
.B2(n_404),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_458),
.B(n_401),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_435),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_440),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_452),
.B(n_415),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_463),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_440),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_480),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_440),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_452),
.A2(n_397),
.B1(n_423),
.B2(n_418),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_467),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_471),
.B(n_379),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_L g545 ( 
.A(n_439),
.B(n_201),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_480),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_476),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_465),
.B(n_170),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_444),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_431),
.A2(n_324),
.B1(n_413),
.B2(n_371),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_456),
.B(n_213),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_L g552 ( 
.A1(n_495),
.A2(n_180),
.B1(n_275),
.B2(n_269),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_470),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_471),
.B(n_386),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_456),
.B(n_309),
.Y(n_555)
);

OAI21xp33_ASAP7_75t_SL g556 ( 
.A1(n_484),
.A2(n_392),
.B(n_391),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_455),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_361),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_470),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_506),
.B(n_403),
.Y(n_562)
);

INVx8_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_466),
.Y(n_564)
);

CKINVDCx6p67_ASAP7_75t_R g565 ( 
.A(n_460),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_449),
.B(n_405),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_456),
.B(n_339),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_480),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_484),
.B(n_401),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_484),
.B(n_421),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_466),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_431),
.A2(n_241),
.B1(n_294),
.B2(n_201),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_466),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_466),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_492),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_439),
.B(n_253),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_454),
.B(n_351),
.Y(n_578)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_486),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_499),
.B(n_421),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_444),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_479),
.B(n_367),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

INVx4_ASAP7_75t_L g584 ( 
.A(n_486),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_429),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_493),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_493),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_499),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_486),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_497),
.B(n_504),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_497),
.B(n_389),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_493),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_430),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_493),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_495),
.A2(n_212),
.B1(n_234),
.B2(n_228),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_486),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_446),
.B(n_362),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_486),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_439),
.B(n_254),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_486),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_433),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_431),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_431),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_493),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_491),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_439),
.B(n_255),
.Y(n_610)
);

NAND2xp33_ASAP7_75t_L g611 ( 
.A(n_450),
.B(n_201),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_446),
.A2(n_362),
.B1(n_345),
.B2(n_366),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_499),
.B(n_425),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_430),
.Y(n_615)
);

BUFx6f_ASAP7_75t_SL g616 ( 
.A(n_499),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_434),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_433),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_437),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_437),
.Y(n_620)
);

OAI22x1_ASAP7_75t_L g621 ( 
.A1(n_467),
.A2(n_179),
.B1(n_181),
.B2(n_183),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_434),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_501),
.B(n_425),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_442),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_460),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_482),
.B(n_437),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_501),
.Y(n_627)
);

CKINVDCx6p67_ASAP7_75t_R g628 ( 
.A(n_500),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_442),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_445),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_504),
.B(n_271),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_437),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_469),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_445),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_482),
.B(n_261),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_491),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_490),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_453),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_457),
.A2(n_241),
.B1(n_294),
.B2(n_427),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_498),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_453),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_498),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_481),
.A2(n_239),
.B1(n_210),
.B2(n_202),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_498),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_443),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_459),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_459),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_504),
.B(n_271),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_443),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_443),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_464),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_450),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_443),
.B(n_270),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_450),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_464),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_447),
.B(n_273),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_468),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_606),
.B(n_438),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_606),
.B(n_241),
.Y(n_660)
);

AND2x4_ASAP7_75t_SL g661 ( 
.A(n_583),
.B(n_271),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_627),
.B(n_457),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_512),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_627),
.B(n_457),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_623),
.B(n_457),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_623),
.B(n_519),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_514),
.B(n_490),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_548),
.B(n_481),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_573),
.B(n_469),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_606),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_517),
.B(n_504),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_606),
.B(n_469),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_513),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_618),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_606),
.B(n_241),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_513),
.Y(n_676)
);

OAI221xp5_ASAP7_75t_L g677 ( 
.A1(n_532),
.A2(n_285),
.B1(n_182),
.B2(n_189),
.C(n_193),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_607),
.B(n_468),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_544),
.B(n_174),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_508),
.A2(n_503),
.B1(n_294),
.B2(n_241),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_607),
.B(n_472),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_521),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_618),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_607),
.B(n_550),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_607),
.B(n_472),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_518),
.B(n_407),
.Y(n_688)
);

AO221x1_ASAP7_75t_L g689 ( 
.A1(n_552),
.A2(n_294),
.B1(n_260),
.B2(n_251),
.C(n_238),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_614),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_607),
.B(n_294),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_626),
.A2(n_448),
.B(n_447),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_614),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_523),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_554),
.B(n_190),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_547),
.B(n_190),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_507),
.B(n_267),
.C(n_263),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_618),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_640),
.B(n_277),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_580),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_635),
.B(n_473),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_534),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_580),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_613),
.B(n_633),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_473),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_527),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_654),
.A2(n_448),
.B(n_447),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_613),
.B(n_199),
.Y(n_709)
);

OAI22xp33_ASAP7_75t_L g710 ( 
.A1(n_558),
.A2(n_322),
.B1(n_198),
.B2(n_188),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_571),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_657),
.A2(n_448),
.B(n_447),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_531),
.B(n_474),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_528),
.B(n_408),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_613),
.B(n_633),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

BUFx8_ASAP7_75t_L g718 ( 
.A(n_616),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_613),
.B(n_200),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_527),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_570),
.B(n_474),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_534),
.A2(n_503),
.B1(n_265),
.B2(n_235),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_547),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_556),
.A2(n_276),
.B(n_204),
.C(n_215),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_535),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_570),
.A2(n_545),
.B1(n_621),
.B2(n_637),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_563),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_585),
.B(n_475),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_585),
.B(n_475),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_633),
.B(n_225),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_591),
.B(n_477),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_577),
.B(n_278),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_524),
.A2(n_279),
.B1(n_280),
.B2(n_283),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_633),
.B(n_229),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_595),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_615),
.B(n_477),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_615),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_617),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_537),
.B(n_191),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_592),
.B(n_191),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_605),
.B(n_410),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_526),
.B(n_410),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_563),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_628),
.B(n_414),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_535),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_SL g747 ( 
.A(n_631),
.B(n_179),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_563),
.B(n_414),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_617),
.B(n_478),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_622),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_528),
.Y(n_751)
);

NAND2xp33_ASAP7_75t_L g752 ( 
.A(n_602),
.B(n_296),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_633),
.B(n_233),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_624),
.B(n_478),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_624),
.B(n_417),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_551),
.B(n_194),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_629),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_600),
.A2(n_272),
.B(n_288),
.C(n_289),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_536),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_616),
.A2(n_304),
.B1(n_306),
.B2(n_308),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_588),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_655),
.B(n_298),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_545),
.A2(n_503),
.B(n_483),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_536),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_629),
.Y(n_765)
);

AND2x2_ASAP7_75t_SL g766 ( 
.A(n_611),
.B(n_300),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_630),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_616),
.A2(n_503),
.B1(n_326),
.B2(n_325),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_555),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_630),
.B(n_483),
.Y(n_770)
);

AO21x2_ASAP7_75t_L g771 ( 
.A1(n_610),
.A2(n_316),
.B(n_331),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_542),
.A2(n_301),
.B1(n_314),
.B2(n_305),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_567),
.B(n_194),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_634),
.B(n_485),
.Y(n_774)
);

BUFx3_ASAP7_75t_L g775 ( 
.A(n_583),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_634),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_588),
.A2(n_328),
.B1(n_310),
.B2(n_320),
.Y(n_777)
);

INVx8_ASAP7_75t_L g778 ( 
.A(n_653),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_562),
.B(n_417),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_576),
.B(n_489),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_638),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_539),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_625),
.B(n_419),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_638),
.B(n_419),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_642),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_642),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_647),
.B(n_485),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_655),
.B(n_197),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_647),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_SL g790 ( 
.A(n_655),
.B(n_197),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_628),
.B(n_426),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_648),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_648),
.B(n_488),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_652),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_652),
.A2(n_340),
.B1(n_328),
.B2(n_326),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_656),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_656),
.B(n_488),
.Y(n_797)
);

INVxp33_ASAP7_75t_L g798 ( 
.A(n_621),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_572),
.B(n_575),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_588),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_598),
.B(n_310),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_575),
.B(n_510),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_541),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_637),
.A2(n_330),
.B1(n_183),
.B2(n_184),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_511),
.B(n_489),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_557),
.B(n_320),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_561),
.B(n_325),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_564),
.B(n_494),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_574),
.B(n_494),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_576),
.B(n_583),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_644),
.B(n_340),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_541),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_612),
.B(n_426),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_649),
.B(n_268),
.Y(n_814)
);

INVx2_ASAP7_75t_SL g815 ( 
.A(n_565),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_SL g816 ( 
.A(n_590),
.B(n_181),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_549),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_619),
.B(n_290),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_565),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_658),
.B(n_502),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_543),
.A2(n_330),
.B1(n_185),
.B2(n_186),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_783),
.Y(n_822)
);

BUFx4f_ASAP7_75t_L g823 ( 
.A(n_716),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_723),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_703),
.B(n_566),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_670),
.B(n_578),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_666),
.B(n_515),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_775),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_701),
.Y(n_829)
);

INVxp33_ASAP7_75t_L g830 ( 
.A(n_742),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_668),
.A2(n_543),
.B1(n_540),
.B2(n_533),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_704),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_685),
.B(n_515),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_670),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_668),
.A2(n_538),
.B1(n_546),
.B2(n_540),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_SL g836 ( 
.A(n_727),
.B(n_653),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_711),
.B(n_582),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_R g838 ( 
.A(n_716),
.B(n_619),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_716),
.B(n_619),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_744),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_791),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_672),
.A2(n_653),
.B(n_560),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_751),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_690),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_811),
.A2(n_538),
.B1(n_568),
.B2(n_525),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_679),
.B(n_620),
.Y(n_846)
);

OR2x6_ASAP7_75t_SL g847 ( 
.A(n_772),
.B(n_184),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_680),
.B(n_516),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_815),
.B(n_427),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_679),
.B(n_620),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_680),
.B(n_516),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_711),
.B(n_620),
.Y(n_852)
);

AND2x6_ASAP7_75t_L g853 ( 
.A(n_670),
.B(n_586),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_660),
.A2(n_560),
.B(n_584),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_743),
.B(n_505),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_693),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_745),
.B(n_505),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_717),
.B(n_525),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_717),
.B(n_632),
.Y(n_859)
);

O2A1O1Ixp5_ASAP7_75t_L g860 ( 
.A1(n_660),
.A2(n_651),
.B(n_650),
.C(n_646),
.Y(n_860)
);

OR2x2_ASAP7_75t_SL g861 ( 
.A(n_698),
.B(n_391),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_751),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_731),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_769),
.A2(n_651),
.B1(n_650),
.B2(n_646),
.Y(n_864)
);

NAND2x1p5_ASAP7_75t_L g865 ( 
.A(n_800),
.B(n_651),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_748),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_667),
.B(n_632),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_662),
.B(n_530),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_811),
.A2(n_530),
.B1(n_533),
.B2(n_546),
.Y(n_869)
);

AND2x4_ASAP7_75t_SL g870 ( 
.A(n_748),
.B(n_290),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_800),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_665),
.A2(n_568),
.B(n_581),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_736),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_718),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_801),
.A2(n_689),
.B1(n_659),
.B2(n_740),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_664),
.B(n_549),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_738),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_663),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_SL g879 ( 
.A1(n_675),
.A2(n_593),
.B(n_587),
.C(n_594),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_702),
.B(n_559),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_739),
.B(n_559),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_800),
.B(n_520),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_751),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_659),
.A2(n_581),
.B1(n_643),
.B2(n_641),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_750),
.B(n_509),
.Y(n_885)
);

NAND3xp33_ASAP7_75t_SL g886 ( 
.A(n_814),
.B(n_338),
.C(n_318),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_757),
.B(n_509),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_765),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_756),
.A2(n_601),
.B1(n_509),
.B2(n_569),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_800),
.B(n_520),
.Y(n_890)
);

BUFx12f_ASAP7_75t_SL g891 ( 
.A(n_748),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_767),
.B(n_553),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_810),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_776),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_714),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_781),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_785),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_756),
.B(n_520),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_786),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_773),
.B(n_520),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_740),
.A2(n_645),
.B1(n_643),
.B2(n_641),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_722),
.A2(n_186),
.B1(n_318),
.B2(n_322),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_741),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_789),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_751),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_792),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_779),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_755),
.B(n_586),
.Y(n_908)
);

INVxp67_ASAP7_75t_SL g909 ( 
.A(n_761),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_794),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_755),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_796),
.B(n_553),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_773),
.B(n_520),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_761),
.Y(n_914)
);

NAND2x1_ASAP7_75t_L g915 ( 
.A(n_673),
.B(n_553),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_696),
.B(n_560),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_674),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_779),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_799),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_780),
.B(n_522),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_820),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_784),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_784),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_676),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_682),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_805),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_688),
.Y(n_927)
);

INVx5_ASAP7_75t_L g928 ( 
.A(n_778),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_813),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_678),
.B(n_569),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_808),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_809),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_681),
.B(n_569),
.Y(n_933)
);

CKINVDCx14_ASAP7_75t_R g934 ( 
.A(n_747),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_802),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_733),
.A2(n_599),
.B1(n_601),
.B2(n_579),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_726),
.B(n_522),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_687),
.B(n_599),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_695),
.B(n_599),
.Y(n_939)
);

AND2x6_ASAP7_75t_L g940 ( 
.A(n_669),
.B(n_814),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_684),
.B(n_392),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_697),
.B(n_579),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_683),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_695),
.B(n_721),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_798),
.B(n_579),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_686),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_752),
.A2(n_601),
.B1(n_596),
.B2(n_584),
.Y(n_947)
);

OR2x4_ASAP7_75t_L g948 ( 
.A(n_741),
.B(n_393),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_699),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_661),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_802),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_806),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_695),
.B(n_645),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_705),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_694),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_695),
.B(n_609),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_SL g957 ( 
.A(n_821),
.B(n_334),
.C(n_336),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_695),
.B(n_609),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_707),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_819),
.Y(n_960)
);

NOR2xp67_ASAP7_75t_L g961 ( 
.A(n_671),
.B(n_587),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_720),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_728),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_729),
.B(n_636),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_732),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_737),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_749),
.B(n_636),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_705),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_715),
.Y(n_969)
);

AND3x1_ASAP7_75t_L g970 ( 
.A(n_804),
.B(n_396),
.C(n_399),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_725),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_816),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_746),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_754),
.B(n_639),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_734),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_806),
.B(n_593),
.Y(n_976)
);

OR2x6_ASAP7_75t_L g977 ( 
.A(n_778),
.B(n_393),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_770),
.Y(n_978)
);

AND2x6_ASAP7_75t_L g979 ( 
.A(n_768),
.B(n_759),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_777),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_774),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_771),
.A2(n_639),
.B1(n_594),
.B2(n_608),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_807),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_787),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_793),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_771),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_764),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_782),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_807),
.A2(n_589),
.B1(n_584),
.B2(n_596),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_726),
.B(n_522),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_760),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_722),
.B(n_522),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_797),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_818),
.B(n_522),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_818),
.B(n_529),
.Y(n_995)
);

AO22x1_ASAP7_75t_L g996 ( 
.A1(n_795),
.A2(n_336),
.B1(n_335),
.B2(n_334),
.Y(n_996)
);

NOR2x1p5_ASAP7_75t_L g997 ( 
.A(n_706),
.B(n_329),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_715),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_SL g999 ( 
.A(n_758),
.B(n_335),
.C(n_332),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_803),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_713),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_963),
.B(n_675),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_825),
.A2(n_788),
.B1(n_700),
.B2(n_719),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_965),
.B(n_691),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_966),
.B(n_691),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_886),
.A2(n_677),
.B1(n_719),
.B2(n_709),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_863),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_944),
.A2(n_778),
.B1(n_788),
.B2(n_762),
.Y(n_1008)
);

AOI21x1_ASAP7_75t_L g1009 ( 
.A1(n_898),
.A2(n_913),
.B(n_900),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_840),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_SL g1011 ( 
.A(n_975),
.B(n_766),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_873),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_978),
.B(n_710),
.Y(n_1013)
);

NOR3xp33_ASAP7_75t_SL g1014 ( 
.A(n_991),
.B(n_821),
.C(n_710),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_SL g1015 ( 
.A(n_893),
.B(n_804),
.C(n_332),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_843),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_944),
.A2(n_762),
.B(n_596),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_822),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_981),
.B(n_812),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_825),
.A2(n_753),
.B1(n_730),
.B2(n_735),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_830),
.B(n_766),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_886),
.A2(n_724),
.B(n_709),
.C(n_753),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_843),
.Y(n_1023)
);

NAND2xp33_ASAP7_75t_SL g1024 ( 
.A(n_911),
.B(n_922),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_877),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_984),
.B(n_817),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_843),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_872),
.A2(n_692),
.B(n_763),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_927),
.B(n_396),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_848),
.A2(n_735),
.B1(n_730),
.B2(n_329),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_911),
.B(n_790),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_903),
.B(n_290),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_857),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_930),
.A2(n_529),
.B(n_603),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_930),
.A2(n_529),
.B(n_603),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_933),
.A2(n_529),
.B(n_603),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_919),
.A2(n_712),
.B1(n_708),
.B2(n_529),
.Y(n_1037)
);

BUFx12f_ASAP7_75t_L g1038 ( 
.A(n_828),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_862),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_862),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_855),
.B(n_399),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_862),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_985),
.A2(n_608),
.B(n_604),
.C(n_597),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_883),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_848),
.A2(n_286),
.B1(n_291),
.B2(n_302),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_933),
.A2(n_603),
.B(n_611),
.Y(n_1046)
);

OR2x6_ASAP7_75t_L g1047 ( 
.A(n_841),
.B(n_604),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_907),
.Y(n_1048)
);

AOI221xp5_ASAP7_75t_SL g1049 ( 
.A1(n_875),
.A2(n_990),
.B1(n_937),
.B2(n_993),
.C(n_858),
.Y(n_1049)
);

BUFx12f_ASAP7_75t_L g1050 ( 
.A(n_824),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_L g1051 ( 
.A(n_837),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_926),
.B(n_303),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_931),
.B(n_932),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_867),
.A2(n_376),
.B(n_3),
.C(n_4),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_922),
.B(n_376),
.Y(n_1055)
);

AND2x2_ASAP7_75t_SL g1056 ( 
.A(n_823),
.B(n_0),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_929),
.B(n_5),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_938),
.A2(n_450),
.B(n_65),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_R g1059 ( 
.A(n_960),
.B(n_56),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_SL g1060 ( 
.A1(n_980),
.A2(n_8),
.B(n_9),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_829),
.Y(n_1061)
);

XNOR2xp5_ASAP7_75t_L g1062 ( 
.A(n_997),
.B(n_69),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_832),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_868),
.A2(n_450),
.B(n_67),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_962),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_851),
.A2(n_11),
.B1(n_14),
.B2(n_16),
.Y(n_1066)
);

AND2x4_ASAP7_75t_SL g1067 ( 
.A(n_922),
.B(n_76),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_846),
.A2(n_11),
.B(n_14),
.C(n_17),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_851),
.A2(n_831),
.B1(n_827),
.B2(n_858),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_837),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_868),
.A2(n_450),
.B(n_90),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_962),
.Y(n_1072)
);

OR2x2_ASAP7_75t_L g1073 ( 
.A(n_844),
.B(n_17),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_1001),
.B(n_952),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_883),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_883),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_921),
.B(n_850),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_998),
.A2(n_95),
.B1(n_153),
.B2(n_152),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_917),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_923),
.B(n_150),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_983),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_888),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_852),
.B(n_450),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_941),
.Y(n_1084)
);

CKINVDCx16_ASAP7_75t_R g1085 ( 
.A(n_874),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_954),
.A2(n_132),
.B1(n_127),
.B2(n_121),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_948),
.B(n_19),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_861),
.Y(n_1088)
);

AOI33xp33_ASAP7_75t_L g1089 ( 
.A1(n_856),
.A2(n_20),
.A3(n_22),
.B1(n_24),
.B2(n_28),
.B3(n_29),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_895),
.B(n_20),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_948),
.B(n_22),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_827),
.A2(n_30),
.B(n_34),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_823),
.B(n_450),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_918),
.B(n_35),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_894),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_842),
.A2(n_833),
.B(n_953),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_896),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_897),
.B(n_35),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_923),
.B(n_118),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_899),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_852),
.B(n_36),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_945),
.A2(n_38),
.B(n_42),
.C(n_45),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_878),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_859),
.B(n_904),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_923),
.B(n_98),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_866),
.Y(n_1106)
);

O2A1O1Ixp5_ASAP7_75t_SL g1107 ( 
.A1(n_994),
.A2(n_995),
.B(n_826),
.C(n_920),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_853),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_941),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_935),
.A2(n_45),
.B(n_52),
.C(n_110),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_SL g1111 ( 
.A1(n_916),
.A2(n_942),
.B(n_934),
.C(n_914),
.Y(n_1111)
);

BUFx8_ASAP7_75t_L g1112 ( 
.A(n_972),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_951),
.A2(n_910),
.B(n_906),
.C(n_976),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_924),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_872),
.A2(n_833),
.B(n_854),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_842),
.A2(n_953),
.B(n_956),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_941),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_881),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_999),
.A2(n_902),
.B(n_957),
.C(n_986),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_999),
.A2(n_902),
.B(n_880),
.C(n_864),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_950),
.Y(n_1121)
);

OAI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_876),
.A2(n_860),
.B(n_956),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_859),
.B(n_880),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_976),
.A2(n_908),
.B(n_992),
.C(n_961),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_849),
.Y(n_1125)
);

AOI221xp5_ASAP7_75t_L g1126 ( 
.A1(n_996),
.A2(n_970),
.B1(n_949),
.B2(n_870),
.C(n_847),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_958),
.A2(n_876),
.B(n_939),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_L g1128 ( 
.A1(n_854),
.A2(n_939),
.B(n_958),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_954),
.A2(n_969),
.B1(n_968),
.B2(n_909),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_SL g1130 ( 
.A1(n_914),
.A2(n_982),
.B(n_869),
.C(n_845),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_891),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_940),
.A2(n_979),
.B1(n_908),
.B2(n_969),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_964),
.B(n_974),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_964),
.A2(n_974),
.B(n_967),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_871),
.A2(n_890),
.B1(n_882),
.B2(n_1000),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_885),
.A2(n_912),
.B(n_892),
.C(n_887),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_881),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_SL g1138 ( 
.A1(n_967),
.A2(n_912),
.B(n_885),
.C(n_887),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_925),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_905),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_892),
.A2(n_955),
.B(n_943),
.C(n_946),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_835),
.A2(n_834),
.B1(n_901),
.B2(n_977),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_928),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_940),
.B(n_979),
.Y(n_1144)
);

A2O1A1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_959),
.A2(n_971),
.B(n_988),
.C(n_987),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_977),
.B(n_849),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1077),
.A2(n_865),
.B1(n_928),
.B2(n_977),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1033),
.B(n_849),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_1018),
.Y(n_1149)
);

NAND3x1_ASAP7_75t_L g1150 ( 
.A(n_1126),
.B(n_889),
.C(n_936),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1053),
.B(n_973),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_1048),
.Y(n_1152)
);

INVx6_ASAP7_75t_L g1153 ( 
.A(n_1050),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1106),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1033),
.B(n_940),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1134),
.A2(n_1096),
.B(n_1133),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1116),
.A2(n_836),
.B(n_928),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1021),
.B(n_979),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1028),
.A2(n_836),
.B(n_928),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1028),
.A2(n_879),
.B(n_989),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_1108),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1127),
.A2(n_947),
.B(n_884),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1027),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1011),
.B(n_979),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1017),
.A2(n_915),
.B(n_853),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1038),
.B(n_853),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1002),
.A2(n_853),
.B(n_838),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1041),
.B(n_1013),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1123),
.B(n_853),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1004),
.A2(n_839),
.B(n_1005),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1009),
.A2(n_1144),
.B(n_1135),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1108),
.A2(n_1122),
.B(n_1136),
.Y(n_1172)
);

AO21x2_ASAP7_75t_L g1173 ( 
.A1(n_1122),
.A2(n_1115),
.B(n_1043),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1118),
.B(n_1137),
.Y(n_1174)
);

NAND2xp33_ASAP7_75t_R g1175 ( 
.A(n_1014),
.B(n_1059),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1070),
.B(n_1079),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1049),
.A2(n_1128),
.B(n_1113),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1069),
.A2(n_1120),
.B(n_1107),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_1037),
.A2(n_1069),
.A3(n_1092),
.B(n_1124),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1143),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_SL g1181 ( 
.A1(n_1015),
.A2(n_1060),
.B(n_1062),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1108),
.A2(n_1115),
.B(n_1130),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1012),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1022),
.A2(n_1119),
.B(n_1003),
.C(n_1011),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1087),
.A2(n_1091),
.B(n_1054),
.C(n_1094),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1056),
.B(n_1051),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1088),
.A2(n_1125),
.B1(n_1132),
.B2(n_1032),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1052),
.B(n_1029),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1025),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1034),
.A2(n_1036),
.B(n_1035),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1046),
.A2(n_1142),
.B(n_1111),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1082),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_SL g1193 ( 
.A(n_1143),
.B(n_1121),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_SL g1194 ( 
.A1(n_1101),
.A2(n_1099),
.B(n_1057),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1088),
.B(n_1074),
.Y(n_1195)
);

AO21x2_ASAP7_75t_L g1196 ( 
.A1(n_1020),
.A2(n_1141),
.B(n_1064),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1031),
.A2(n_1055),
.B(n_1019),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1026),
.A2(n_1051),
.B(n_1129),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1006),
.A2(n_1049),
.B(n_1060),
.C(n_1068),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1102),
.B(n_1110),
.C(n_1045),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_1027),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1104),
.B(n_1063),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1010),
.B(n_1081),
.Y(n_1203)
);

NAND3xp33_ASAP7_75t_L g1204 ( 
.A(n_1045),
.B(n_1066),
.C(n_1089),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1095),
.A2(n_1097),
.B1(n_1100),
.B2(n_1061),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1138),
.A2(n_1058),
.B(n_1071),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1024),
.A2(n_1109),
.B1(n_1084),
.B2(n_1117),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1030),
.A2(n_1066),
.A3(n_1145),
.B(n_1078),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1030),
.A2(n_1105),
.B(n_1080),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1139),
.B(n_1114),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1027),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1083),
.A2(n_1086),
.B(n_1103),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1065),
.B(n_1072),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1016),
.A2(n_1098),
.B(n_1090),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1073),
.B(n_1140),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_1131),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1047),
.Y(n_1217)
);

INVx8_ASAP7_75t_L g1218 ( 
.A(n_1039),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1093),
.A2(n_1146),
.B(n_1067),
.Y(n_1219)
);

INVx6_ASAP7_75t_L g1220 ( 
.A(n_1112),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1146),
.B(n_1047),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1023),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1040),
.A2(n_1076),
.B(n_1042),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1040),
.A2(n_1076),
.B(n_1044),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1042),
.B(n_1044),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1044),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1075),
.A2(n_1096),
.A3(n_1043),
.B(n_1116),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1085),
.A2(n_679),
.B1(n_1011),
.B2(n_345),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1075),
.A2(n_1008),
.B(n_800),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1075),
.B(n_1053),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1027),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1069),
.A2(n_1077),
.B(n_1120),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1077),
.A2(n_1053),
.B1(n_975),
.B2(n_680),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1022),
.A2(n_679),
.B(n_668),
.C(n_903),
.Y(n_1236)
);

AOI221x1_ASAP7_75t_L g1237 ( 
.A1(n_1066),
.A2(n_679),
.B1(n_886),
.B2(n_1068),
.C(n_1096),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1096),
.A2(n_1043),
.A3(n_1116),
.B(n_1037),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_L g1239 ( 
.A1(n_1031),
.A2(n_679),
.B(n_671),
.C(n_696),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1118),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1033),
.B(n_830),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1027),
.Y(n_1244)
);

NAND3x1_ASAP7_75t_L g1245 ( 
.A(n_1126),
.B(n_667),
.C(n_801),
.Y(n_1245)
);

NOR2xp67_ASAP7_75t_SL g1246 ( 
.A(n_1050),
.B(n_775),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1022),
.A2(n_679),
.B(n_668),
.C(n_903),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_SL g1248 ( 
.A1(n_1092),
.A2(n_1132),
.B(n_1144),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1128),
.A2(n_1116),
.B(n_1035),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1011),
.A2(n_542),
.B1(n_975),
.B2(n_903),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1014),
.B(n_679),
.C(n_667),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1033),
.B(n_830),
.Y(n_1252)
);

OAI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1088),
.A2(n_667),
.B1(n_975),
.B2(n_903),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1011),
.A2(n_679),
.B1(n_345),
.B2(n_366),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1007),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1014),
.B(n_679),
.C(n_667),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1134),
.A2(n_670),
.B(n_1096),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_SL g1258 ( 
.A(n_1079),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1007),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_L g1261 ( 
.A(n_1077),
.B(n_716),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1134),
.A2(n_670),
.B(n_1096),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1134),
.A2(n_670),
.B(n_1096),
.Y(n_1263)
);

AO22x2_ASAP7_75t_L g1264 ( 
.A1(n_1060),
.A2(n_1066),
.B1(n_886),
.B2(n_1015),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1265)
);

OAI22x1_ASAP7_75t_L g1266 ( 
.A1(n_1088),
.A2(n_667),
.B1(n_975),
.B2(n_903),
.Y(n_1266)
);

INVxp67_ASAP7_75t_L g1267 ( 
.A(n_1018),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1128),
.A2(n_1116),
.B(n_1035),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1128),
.A2(n_1116),
.B(n_1035),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1049),
.A2(n_1096),
.B(n_1116),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1272)
);

BUFx3_ASAP7_75t_L g1273 ( 
.A(n_1079),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1007),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1053),
.B(n_1077),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1050),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1128),
.A2(n_1116),
.B(n_1035),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1128),
.A2(n_1116),
.B(n_1035),
.Y(n_1278)
);

A2O1A1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1022),
.A2(n_679),
.B(n_668),
.C(n_903),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1118),
.Y(n_1280)
);

AO32x2_ASAP7_75t_L g1281 ( 
.A1(n_1066),
.A2(n_1069),
.A3(n_1030),
.B1(n_1142),
.B2(n_1045),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1018),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1022),
.A2(n_679),
.B(n_668),
.C(n_903),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1118),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1033),
.B(n_822),
.Y(n_1285)
);

AOI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1011),
.A2(n_679),
.B1(n_345),
.B2(n_366),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1119),
.A2(n_679),
.B(n_544),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1232),
.B(n_1233),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1219),
.B(n_1229),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1285),
.B(n_1215),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1257),
.A2(n_1263),
.B(n_1262),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1254),
.A2(n_1286),
.B1(n_1251),
.B2(n_1256),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1168),
.B(n_1188),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1182),
.A2(n_1191),
.A3(n_1237),
.B(n_1172),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1179),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1264),
.A2(n_1287),
.B1(n_1204),
.B2(n_1200),
.Y(n_1296)
);

BUFx8_ASAP7_75t_L g1297 ( 
.A(n_1258),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1161),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1282),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1241),
.B(n_1242),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1247),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1156),
.A2(n_1157),
.B(n_1159),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1201),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1203),
.B(n_1149),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1259),
.B(n_1265),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1283),
.A2(n_1234),
.B(n_1184),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1154),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1165),
.A2(n_1249),
.B(n_1268),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1186),
.A2(n_1264),
.B1(n_1164),
.B2(n_1235),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1269),
.A2(n_1277),
.B(n_1278),
.Y(n_1310)
);

AND2x2_ASAP7_75t_SL g1311 ( 
.A(n_1166),
.B(n_1281),
.Y(n_1311)
);

OA21x2_ASAP7_75t_L g1312 ( 
.A1(n_1178),
.A2(n_1206),
.B(n_1160),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1190),
.A2(n_1162),
.B(n_1171),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1199),
.A2(n_1185),
.B(n_1275),
.C(n_1272),
.Y(n_1314)
);

INVx4_ASAP7_75t_SL g1315 ( 
.A(n_1220),
.Y(n_1315)
);

NAND2x1p5_ASAP7_75t_L g1316 ( 
.A(n_1201),
.B(n_1211),
.Y(n_1316)
);

INVxp33_ASAP7_75t_L g1317 ( 
.A(n_1195),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1228),
.A2(n_1253),
.B1(n_1266),
.B2(n_1220),
.Y(n_1318)
);

AO32x2_ASAP7_75t_L g1319 ( 
.A1(n_1281),
.A2(n_1205),
.A3(n_1147),
.B1(n_1179),
.B2(n_1248),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1194),
.A2(n_1197),
.B(n_1167),
.Y(n_1320)
);

OAI222xp33_ASAP7_75t_L g1321 ( 
.A1(n_1250),
.A2(n_1271),
.B1(n_1174),
.B2(n_1280),
.C1(n_1240),
.C2(n_1284),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1183),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1270),
.A2(n_1170),
.B(n_1196),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1189),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1179),
.Y(n_1325)
);

AO21x2_ASAP7_75t_L g1326 ( 
.A1(n_1173),
.A2(n_1155),
.B(n_1209),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1239),
.A2(n_1284),
.B(n_1280),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1151),
.B(n_1158),
.Y(n_1328)
);

OAI21xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1169),
.A2(n_1230),
.B(n_1202),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1176),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1217),
.A2(n_1214),
.B(n_1260),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1227),
.Y(n_1332)
);

OA21x2_ASAP7_75t_L g1333 ( 
.A1(n_1255),
.A2(n_1274),
.B(n_1210),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1175),
.A2(n_1245),
.B1(n_1181),
.B2(n_1187),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1267),
.A2(n_1148),
.B(n_1261),
.C(n_1152),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1276),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1209),
.A2(n_1212),
.B(n_1225),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1177),
.A2(n_1270),
.B(n_1221),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1213),
.B(n_1176),
.Y(n_1339)
);

AO31x2_ASAP7_75t_L g1340 ( 
.A1(n_1238),
.A2(n_1177),
.A3(n_1227),
.B(n_1208),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1238),
.A2(n_1227),
.B(n_1180),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1150),
.B(n_1208),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1223),
.A2(n_1207),
.B(n_1224),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1222),
.A2(n_1193),
.B(n_1246),
.C(n_1218),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1226),
.B(n_1211),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1163),
.B(n_1231),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1211),
.A2(n_1218),
.B(n_1163),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1153),
.A2(n_1216),
.B1(n_1244),
.B2(n_1258),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1153),
.A2(n_1287),
.B(n_1247),
.C(n_1279),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1244),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1244),
.A2(n_1287),
.B(n_1256),
.C(n_1251),
.Y(n_1351)
);

NAND3xp33_ASAP7_75t_L g1352 ( 
.A(n_1287),
.B(n_679),
.C(n_1251),
.Y(n_1352)
);

OAI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1257),
.A2(n_1263),
.B(n_1262),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1179),
.Y(n_1354)
);

OAI211xp5_ASAP7_75t_L g1355 ( 
.A1(n_1287),
.A2(n_667),
.B(n_1014),
.C(n_804),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1251),
.A2(n_1256),
.B1(n_667),
.B2(n_1264),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1251),
.A2(n_1256),
.B1(n_667),
.B2(n_1264),
.Y(n_1357)
);

AO31x2_ASAP7_75t_L g1358 ( 
.A1(n_1182),
.A2(n_1191),
.A3(n_1237),
.B(n_1172),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1192),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1257),
.A2(n_1263),
.B(n_1262),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1232),
.B(n_1233),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1219),
.B(n_1229),
.Y(n_1362)
);

NAND2x1p5_ASAP7_75t_L g1363 ( 
.A(n_1161),
.B(n_1108),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1243),
.B(n_1252),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1251),
.A2(n_1256),
.B1(n_667),
.B2(n_1264),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1257),
.A2(n_1263),
.B(n_1262),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1201),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1285),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1232),
.B(n_1233),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1287),
.B(n_679),
.C(n_1251),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1192),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1161),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1243),
.B(n_1252),
.Y(n_1373)
);

INVx5_ASAP7_75t_L g1374 ( 
.A(n_1161),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1236),
.A2(n_1279),
.B(n_1247),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1287),
.A2(n_1236),
.B(n_1279),
.C(n_1247),
.Y(n_1376)
);

AOI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1172),
.A2(n_1182),
.B(n_1159),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1216),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1251),
.A2(n_1256),
.B1(n_667),
.B2(n_1264),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1176),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1248),
.A2(n_1092),
.B(n_1198),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1273),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1254),
.A2(n_1011),
.B1(n_1286),
.B2(n_1256),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1273),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1243),
.B(n_1252),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1250),
.B(n_345),
.Y(n_1386)
);

INVx5_ASAP7_75t_L g1387 ( 
.A(n_1161),
.Y(n_1387)
);

OAI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1254),
.A2(n_1011),
.B1(n_1286),
.B2(n_1256),
.Y(n_1388)
);

CKINVDCx9p33_ASAP7_75t_R g1389 ( 
.A(n_1195),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1191),
.A2(n_1178),
.B(n_1172),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1232),
.A2(n_680),
.B1(n_1241),
.B2(n_1233),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1287),
.A2(n_1256),
.B(n_1251),
.C(n_679),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1219),
.B(n_1229),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1276),
.B(n_824),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1287),
.A2(n_1256),
.B(n_1251),
.C(n_679),
.Y(n_1395)
);

BUFx2_ASAP7_75t_L g1396 ( 
.A(n_1176),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1273),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1327),
.Y(n_1398)
);

AOI221x1_ASAP7_75t_SL g1399 ( 
.A1(n_1292),
.A2(n_1383),
.B1(n_1388),
.B2(n_1386),
.C(n_1370),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1288),
.B(n_1300),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1364),
.B(n_1373),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1368),
.B(n_1290),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1288),
.B(n_1300),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1328),
.B(n_1385),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1391),
.A2(n_1395),
.B(n_1392),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1305),
.B(n_1361),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1305),
.B(n_1361),
.Y(n_1407)
);

O2A1O1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1292),
.A2(n_1383),
.B(n_1388),
.C(n_1355),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1334),
.B(n_1328),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1339),
.B(n_1293),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1309),
.B(n_1330),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1309),
.B(n_1380),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1396),
.B(n_1315),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1369),
.B(n_1314),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1317),
.A2(n_1296),
.B1(n_1379),
.B2(n_1357),
.Y(n_1415)
);

BUFx3_ASAP7_75t_L g1416 ( 
.A(n_1382),
.Y(n_1416)
);

NOR2x1_ASAP7_75t_SL g1417 ( 
.A(n_1289),
.B(n_1362),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1296),
.A2(n_1357),
.B1(n_1365),
.B2(n_1356),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1391),
.A2(n_1349),
.B(n_1344),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1299),
.B(n_1307),
.Y(n_1420)
);

CKINVDCx6p67_ASAP7_75t_R g1421 ( 
.A(n_1336),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1350),
.B(n_1307),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1302),
.A2(n_1306),
.B(n_1291),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1315),
.B(n_1345),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1299),
.B(n_1304),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1359),
.Y(n_1426)
);

BUFx12f_ASAP7_75t_L g1427 ( 
.A(n_1297),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1318),
.A2(n_1352),
.B1(n_1306),
.B2(n_1351),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1301),
.A2(n_1375),
.B(n_1323),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1322),
.B(n_1324),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1311),
.A2(n_1342),
.B1(n_1393),
.B2(n_1362),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1303),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1301),
.A2(n_1375),
.B(n_1323),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_R g1434 ( 
.A(n_1394),
.B(n_1378),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1329),
.B(n_1349),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1335),
.B(n_1371),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1342),
.A2(n_1311),
.B(n_1343),
.C(n_1320),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1331),
.B(n_1333),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1313),
.A2(n_1341),
.B(n_1353),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1341),
.A2(n_1360),
.B(n_1366),
.Y(n_1440)
);

NOR2xp67_ASAP7_75t_L g1441 ( 
.A(n_1298),
.B(n_1372),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1397),
.Y(n_1442)
);

AOI21xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1289),
.A2(n_1393),
.B(n_1362),
.Y(n_1443)
);

AOI221xp5_ASAP7_75t_L g1444 ( 
.A1(n_1376),
.A2(n_1321),
.B1(n_1381),
.B2(n_1348),
.C(n_1325),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1345),
.B(n_1390),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1315),
.B(n_1346),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1338),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1294),
.B(n_1358),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1326),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1319),
.B(n_1298),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1316),
.A2(n_1367),
.B(n_1303),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1294),
.B(n_1358),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1389),
.A2(n_1384),
.B1(n_1316),
.B2(n_1367),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1303),
.A2(n_1367),
.B1(n_1363),
.B2(n_1387),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1294),
.B(n_1358),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1347),
.B(n_1387),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1374),
.B(n_1387),
.Y(n_1457)
);

NOR2xp33_ASAP7_75t_R g1458 ( 
.A(n_1297),
.B(n_1387),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1363),
.A2(n_1374),
.B1(n_1354),
.B2(n_1332),
.Y(n_1459)
);

AOI21x1_ASAP7_75t_SL g1460 ( 
.A1(n_1319),
.A2(n_1377),
.B(n_1326),
.Y(n_1460)
);

O2A1O1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1337),
.A2(n_1312),
.B(n_1319),
.C(n_1340),
.Y(n_1461)
);

O2A1O1Ixp33_ASAP7_75t_L g1462 ( 
.A1(n_1312),
.A2(n_1319),
.B(n_1340),
.C(n_1374),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1374),
.A2(n_667),
.B1(n_1292),
.B2(n_1306),
.C(n_1287),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1308),
.Y(n_1464)
);

O2A1O1Ixp5_ASAP7_75t_L g1465 ( 
.A1(n_1340),
.A2(n_1287),
.B(n_1306),
.C(n_1301),
.Y(n_1465)
);

AOI21x1_ASAP7_75t_SL g1466 ( 
.A1(n_1310),
.A2(n_1342),
.B(n_1144),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1382),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1386),
.A2(n_1287),
.B(n_679),
.C(n_1256),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1330),
.B(n_1221),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1288),
.B(n_1300),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1386),
.A2(n_1286),
.B1(n_1254),
.B2(n_1245),
.Y(n_1471)
);

O2A1O1Ixp5_ASAP7_75t_L g1472 ( 
.A1(n_1306),
.A2(n_1287),
.B(n_1375),
.C(n_1301),
.Y(n_1472)
);

AOI21x1_ASAP7_75t_SL g1473 ( 
.A1(n_1342),
.A2(n_1144),
.B(n_1295),
.Y(n_1473)
);

NOR2x1_ASAP7_75t_SL g1474 ( 
.A(n_1289),
.B(n_1362),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1292),
.A2(n_1287),
.B(n_1395),
.C(n_1392),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1288),
.B(n_1300),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1303),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1330),
.B(n_1221),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1327),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1382),
.Y(n_1480)
);

NOR2x1_ASAP7_75t_SL g1481 ( 
.A(n_1289),
.B(n_1362),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1429),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1443),
.B(n_1423),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1448),
.B(n_1452),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1455),
.B(n_1398),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1445),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1417),
.B(n_1474),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1435),
.B(n_1400),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1426),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1429),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1479),
.B(n_1447),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1481),
.B(n_1464),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

INVx1_ASAP7_75t_SL g1496 ( 
.A(n_1425),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1437),
.B(n_1462),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1461),
.B(n_1465),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1464),
.B(n_1456),
.Y(n_1499)
);

AO21x2_ASAP7_75t_L g1500 ( 
.A1(n_1405),
.A2(n_1419),
.B(n_1468),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1440),
.Y(n_1501)
);

AO21x2_ASAP7_75t_L g1502 ( 
.A1(n_1475),
.A2(n_1459),
.B(n_1431),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1439),
.B(n_1430),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1472),
.A2(n_1444),
.B(n_1463),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1466),
.A2(n_1460),
.B(n_1473),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1409),
.B(n_1422),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1463),
.A2(n_1475),
.B(n_1414),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1457),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1408),
.A2(n_1428),
.B(n_1418),
.Y(n_1509)
);

OAI211xp5_ASAP7_75t_L g1510 ( 
.A1(n_1408),
.A2(n_1471),
.B(n_1444),
.C(n_1415),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1402),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1436),
.Y(n_1512)
);

BUFx2_ASAP7_75t_R g1513 ( 
.A(n_1480),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1403),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1406),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1407),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1495),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1494),
.B(n_1412),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1512),
.B(n_1470),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1490),
.Y(n_1521)
);

INVx3_ASAP7_75t_SL g1522 ( 
.A(n_1483),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1494),
.B(n_1411),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1482),
.B(n_1491),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1512),
.B(n_1476),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1503),
.B(n_1401),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1482),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1487),
.B(n_1399),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1487),
.B(n_1410),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1509),
.A2(n_1404),
.B1(n_1478),
.B2(n_1469),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1487),
.B(n_1420),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1488),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1501),
.Y(n_1533)
);

INVx2_ASAP7_75t_SL g1534 ( 
.A(n_1492),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1510),
.A2(n_1453),
.B1(n_1413),
.B2(n_1424),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1484),
.B(n_1441),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1493),
.B(n_1446),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_L g1538 ( 
.A(n_1500),
.B(n_1451),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1528),
.A2(n_1510),
.B1(n_1507),
.B2(n_1513),
.Y(n_1539)
);

AOI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1528),
.A2(n_1504),
.B1(n_1507),
.B2(n_1497),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1521),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1533),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1538),
.B(n_1489),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1532),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1517),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1530),
.A2(n_1500),
.B1(n_1509),
.B2(n_1504),
.Y(n_1546)
);

INVx5_ASAP7_75t_SL g1547 ( 
.A(n_1527),
.Y(n_1547)
);

OAI211xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1520),
.A2(n_1489),
.B(n_1511),
.C(n_1496),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1533),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1533),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1538),
.B(n_1483),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1535),
.A2(n_1509),
.B1(n_1500),
.B2(n_1504),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1521),
.Y(n_1553)
);

AOI33xp33_ASAP7_75t_L g1554 ( 
.A1(n_1530),
.A2(n_1497),
.A3(n_1498),
.B1(n_1511),
.B2(n_1515),
.B3(n_1514),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.B(n_1484),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1538),
.A2(n_1497),
.B(n_1504),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1521),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1531),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1535),
.A2(n_1500),
.B1(n_1509),
.B2(n_1504),
.Y(n_1559)
);

OAI31xp33_ASAP7_75t_L g1560 ( 
.A1(n_1520),
.A2(n_1500),
.A3(n_1509),
.B(n_1498),
.Y(n_1560)
);

AO21x1_ASAP7_75t_SL g1561 ( 
.A1(n_1536),
.A2(n_1485),
.B(n_1486),
.Y(n_1561)
);

AOI222xp33_ASAP7_75t_L g1562 ( 
.A1(n_1525),
.A2(n_1427),
.B1(n_1498),
.B2(n_1516),
.C1(n_1514),
.C2(n_1515),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1531),
.B(n_1506),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1534),
.B(n_1484),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1525),
.A2(n_1513),
.B1(n_1504),
.B2(n_1483),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1537),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1537),
.Y(n_1567)
);

OAI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1522),
.A2(n_1483),
.B1(n_1508),
.B2(n_1516),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1527),
.Y(n_1569)
);

INVxp67_ASAP7_75t_SL g1570 ( 
.A(n_1543),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1561),
.B(n_1524),
.Y(n_1571)
);

INVx4_ASAP7_75t_SL g1572 ( 
.A(n_1551),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

INVx1_ASAP7_75t_SL g1574 ( 
.A(n_1545),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1542),
.Y(n_1575)
);

OAI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1539),
.A2(n_1483),
.B(n_1536),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_SL g1577 ( 
.A1(n_1539),
.A2(n_1552),
.B(n_1560),
.Y(n_1577)
);

AND2x2_ASAP7_75t_SL g1578 ( 
.A(n_1554),
.B(n_1488),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

AND2x6_ASAP7_75t_L g1580 ( 
.A(n_1547),
.B(n_1488),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1544),
.Y(n_1582)
);

INVxp67_ASAP7_75t_SL g1583 ( 
.A(n_1542),
.Y(n_1583)
);

INVx4_ASAP7_75t_L g1584 ( 
.A(n_1569),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1549),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1541),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1540),
.A2(n_1483),
.B(n_1505),
.Y(n_1587)
);

BUFx3_ASAP7_75t_L g1588 ( 
.A(n_1569),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1569),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1569),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1553),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1561),
.B(n_1524),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1553),
.Y(n_1593)
);

INVx4_ASAP7_75t_SL g1594 ( 
.A(n_1551),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1557),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1555),
.B(n_1564),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1540),
.B(n_1526),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1544),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1550),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1551),
.B(n_1483),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1566),
.B(n_1519),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1573),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1570),
.B(n_1562),
.Y(n_1605)
);

OR2x6_ASAP7_75t_L g1606 ( 
.A(n_1577),
.B(n_1551),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1597),
.B(n_1558),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1597),
.B(n_1574),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1570),
.B(n_1562),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1578),
.B(n_1560),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1573),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1571),
.B(n_1566),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1586),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1586),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1572),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1596),
.B(n_1563),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1574),
.B(n_1529),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1591),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1572),
.B(n_1566),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1578),
.B(n_1526),
.Y(n_1621)
);

NOR2x1p5_ASAP7_75t_L g1622 ( 
.A(n_1571),
.B(n_1421),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1582),
.B(n_1599),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1572),
.B(n_1567),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1579),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1571),
.B(n_1567),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1592),
.B(n_1581),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1579),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1592),
.B(n_1567),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1577),
.B(n_1552),
.C(n_1559),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1578),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1593),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1576),
.A2(n_1578),
.B1(n_1565),
.B2(n_1502),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1572),
.B(n_1532),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1547),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1582),
.B(n_1526),
.Y(n_1638)
);

CKINVDCx14_ASAP7_75t_R g1639 ( 
.A(n_1580),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1599),
.B(n_1523),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1588),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1585),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1595),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1623),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1643),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1622),
.B(n_1572),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1523),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1607),
.B(n_1595),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1623),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1627),
.B(n_1581),
.Y(n_1650)
);

NAND3xp33_ASAP7_75t_L g1651 ( 
.A(n_1631),
.B(n_1576),
.C(n_1587),
.Y(n_1651)
);

NOR2x1_ASAP7_75t_L g1652 ( 
.A(n_1610),
.B(n_1584),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1625),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1609),
.B(n_1416),
.Y(n_1654)
);

OAI21xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1610),
.A2(n_1587),
.B(n_1602),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1628),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1630),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1627),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1633),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1603),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1603),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1613),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_L g1664 ( 
.A(n_1608),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1632),
.B(n_1523),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1635),
.B(n_1518),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1594),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1614),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1641),
.B(n_1518),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1641),
.B(n_1518),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1617),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1634),
.B(n_1594),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1606),
.Y(n_1673)
);

NAND2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1637),
.B(n_1434),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1619),
.Y(n_1675)
);

INVx1_ASAP7_75t_SL g1676 ( 
.A(n_1618),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1642),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1642),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1620),
.B(n_1594),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1649),
.B(n_1607),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1667),
.B(n_1606),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1651),
.A2(n_1606),
.B1(n_1601),
.B2(n_1639),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1644),
.B(n_1606),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1653),
.Y(n_1684)
);

AND3x2_ASAP7_75t_L g1685 ( 
.A(n_1664),
.B(n_1637),
.C(n_1624),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1667),
.B(n_1612),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1672),
.B(n_1612),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1672),
.B(n_1650),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1659),
.Y(n_1689)
);

NOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1652),
.B(n_1649),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1652),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1655),
.A2(n_1502),
.B1(n_1556),
.B2(n_1546),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1674),
.A2(n_1601),
.B1(n_1639),
.B2(n_1502),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1657),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1653),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1650),
.B(n_1626),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1679),
.B(n_1620),
.Y(n_1697)
);

INVxp67_ASAP7_75t_L g1698 ( 
.A(n_1654),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1645),
.B(n_1620),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1676),
.B(n_1616),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1657),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1646),
.B(n_1626),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1621),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1657),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1646),
.B(n_1629),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1699),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1680),
.B(n_1647),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1688),
.B(n_1659),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1699),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1689),
.Y(n_1710)
);

INVxp67_ASAP7_75t_L g1711 ( 
.A(n_1688),
.Y(n_1711)
);

AOI21xp33_ASAP7_75t_L g1712 ( 
.A1(n_1683),
.A2(n_1657),
.B(n_1663),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1692),
.A2(n_1666),
.B1(n_1646),
.B2(n_1679),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1701),
.B(n_1645),
.Y(n_1714)
);

AOI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1692),
.A2(n_1679),
.B1(n_1624),
.B2(n_1636),
.Y(n_1715)
);

AOI211xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1698),
.A2(n_1679),
.B(n_1663),
.C(n_1675),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1689),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1686),
.A2(n_1624),
.B1(n_1636),
.B2(n_1601),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1691),
.A2(n_1670),
.B1(n_1669),
.B2(n_1636),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1689),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1681),
.B(n_1668),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1681),
.B(n_1668),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1694),
.B(n_1671),
.Y(n_1723)
);

OAI31xp33_ASAP7_75t_L g1724 ( 
.A1(n_1691),
.A2(n_1671),
.A3(n_1675),
.B(n_1548),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1690),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1711),
.B(n_1704),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1710),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1716),
.B(n_1696),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1717),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1713),
.A2(n_1686),
.B1(n_1687),
.B2(n_1705),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1707),
.B(n_1680),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1708),
.B(n_1696),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1720),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1721),
.B(n_1694),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1722),
.B(n_1687),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1719),
.A2(n_1705),
.B1(n_1702),
.B2(n_1682),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1706),
.B(n_1694),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1735),
.B(n_1709),
.Y(n_1738)
);

OAI211xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1728),
.A2(n_1712),
.B(n_1724),
.C(n_1690),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1726),
.Y(n_1740)
);

AOI211xp5_ASAP7_75t_L g1741 ( 
.A1(n_1734),
.A2(n_1725),
.B(n_1724),
.C(n_1714),
.Y(n_1741)
);

OAI222xp33_ASAP7_75t_L g1742 ( 
.A1(n_1736),
.A2(n_1715),
.B1(n_1718),
.B2(n_1730),
.C1(n_1694),
.C2(n_1693),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1731),
.B(n_1697),
.Y(n_1743)
);

OAI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1732),
.A2(n_1700),
.B1(n_1703),
.B2(n_1702),
.Y(n_1744)
);

AOI211xp5_ASAP7_75t_L g1745 ( 
.A1(n_1726),
.A2(n_1697),
.B(n_1723),
.C(n_1700),
.Y(n_1745)
);

AOI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1737),
.A2(n_1723),
.B(n_1695),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1727),
.B(n_1648),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1729),
.A2(n_1695),
.B1(n_1684),
.B2(n_1697),
.C(n_1656),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1747),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1739),
.A2(n_1733),
.B1(n_1684),
.B2(n_1656),
.C(n_1658),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1738),
.B(n_1697),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1740),
.A2(n_1685),
.B1(n_1434),
.B2(n_1458),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1745),
.B(n_1658),
.Y(n_1753)
);

XOR2xp5_ASAP7_75t_L g1754 ( 
.A(n_1743),
.B(n_1744),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1741),
.A2(n_1660),
.B1(n_1594),
.B2(n_1580),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1749),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1753),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1754),
.A2(n_1742),
.B(n_1748),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1751),
.B(n_1746),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1750),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1755),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1752),
.B(n_1648),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1754),
.A2(n_1660),
.B1(n_1677),
.B2(n_1662),
.C(n_1678),
.Y(n_1763)
);

AOI322xp5_ASAP7_75t_L g1764 ( 
.A1(n_1759),
.A2(n_1678),
.A3(n_1677),
.B1(n_1661),
.B2(n_1662),
.C1(n_1665),
.C2(n_1629),
.Y(n_1764)
);

INVx1_ASAP7_75t_SL g1765 ( 
.A(n_1756),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1758),
.A2(n_1661),
.B1(n_1584),
.B2(n_1588),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1760),
.Y(n_1767)
);

OA211x2_ASAP7_75t_L g1768 ( 
.A1(n_1763),
.A2(n_1640),
.B(n_1638),
.C(n_1556),
.Y(n_1768)
);

AND4x1_ASAP7_75t_L g1769 ( 
.A(n_1767),
.B(n_1757),
.C(n_1762),
.D(n_1761),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1765),
.Y(n_1770)
);

OA22x2_ASAP7_75t_L g1771 ( 
.A1(n_1766),
.A2(n_1584),
.B1(n_1604),
.B2(n_1611),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1770),
.B(n_1442),
.Y(n_1772)
);

AOI322xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1769),
.A3(n_1768),
.B1(n_1771),
.B2(n_1764),
.C1(n_1589),
.C2(n_1588),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1773),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1773),
.B(n_1467),
.Y(n_1775)
);

NAND2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1775),
.B(n_1413),
.Y(n_1776)
);

AO22x2_ASAP7_75t_L g1777 ( 
.A1(n_1774),
.A2(n_1604),
.B1(n_1611),
.B2(n_1584),
.Y(n_1777)
);

AOI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1584),
.B(n_1590),
.Y(n_1778)
);

AO22x2_ASAP7_75t_L g1779 ( 
.A1(n_1776),
.A2(n_1589),
.B1(n_1594),
.B2(n_1598),
.Y(n_1779)
);

OAI22xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1779),
.A2(n_1458),
.B1(n_1590),
.B2(n_1589),
.Y(n_1780)
);

INVxp33_ASAP7_75t_SL g1781 ( 
.A(n_1780),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1781),
.B(n_1778),
.Y(n_1782)
);

AOI322xp5_ASAP7_75t_L g1783 ( 
.A1(n_1782),
.A2(n_1590),
.A3(n_1575),
.B1(n_1583),
.B2(n_1602),
.C1(n_1568),
.C2(n_1600),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1590),
.B1(n_1575),
.B2(n_1583),
.Y(n_1784)
);

AOI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1454),
.B(n_1432),
.C(n_1477),
.Y(n_1785)
);


endmodule