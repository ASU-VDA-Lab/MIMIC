module fake_jpeg_31067_n_121 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_1),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_5),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_5),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_3),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_24),
.Y(n_49)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_15),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_32),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_57),
.B(n_59),
.C(n_62),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_26),
.B1(n_28),
.B2(n_19),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_40),
.B1(n_44),
.B2(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_23),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_36),
.B1(n_27),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_60),
.A2(n_64),
.B1(n_66),
.B2(n_68),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_13),
.B(n_17),
.C(n_16),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_16),
.B1(n_22),
.B2(n_31),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_16),
.B1(n_14),
.B2(n_24),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_22),
.B1(n_14),
.B2(n_1),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_4),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_57),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_40),
.B1(n_44),
.B2(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_79),
.A2(n_65),
.B1(n_62),
.B2(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_87),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_54),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_88),
.C(n_65),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_60),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_74),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.C(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_96),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_70),
.C(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_70),
.B(n_74),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_53),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_80),
.B1(n_64),
.B2(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_95),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_2),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_52),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_104),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_106),
.B(n_102),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_53),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_114),
.B(n_6),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.C(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_110),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_4),
.B(n_7),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_8),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g121 ( 
.A(n_120),
.Y(n_121)
);


endmodule