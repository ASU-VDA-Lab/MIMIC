module fake_netlist_6_3768_n_726 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_726);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_726;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_608;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_527;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g153 ( 
.A(n_34),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_68),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_86),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_20),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_41),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_15),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_48),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_44),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_35),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_7),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_13),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_0),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_66),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_4),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_7),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_9),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_83),
.Y(n_184)
);

BUFx8_ASAP7_75t_SL g185 ( 
.A(n_130),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_42),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_124),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_131),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_36),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_69),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_101),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_62),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_100),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_33),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_73),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_43),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_102),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_64),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g211 ( 
.A(n_156),
.B(n_0),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_159),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_1),
.B(n_2),
.Y(n_214)
);

OAI22x1_ASAP7_75t_L g215 ( 
.A1(n_172),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_3),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_204),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_175),
.B(n_8),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

OAI21x1_ASAP7_75t_L g233 ( 
.A1(n_179),
.A2(n_84),
.B(n_151),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_9),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g238 ( 
.A(n_168),
.B(n_10),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

BUFx8_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_186),
.B(n_10),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

CKINVDCx11_ASAP7_75t_R g245 ( 
.A(n_158),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_174),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_246)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_158),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_11),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_154),
.B(n_12),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_205),
.Y(n_253)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_208),
.Y(n_257)
);

AO21x2_ASAP7_75t_L g258 ( 
.A1(n_229),
.A2(n_200),
.B(n_203),
.Y(n_258)
);

NAND2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_155),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_164),
.Y(n_260)
);

BUFx10_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_213),
.B(n_166),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

NAND2xp33_ASAP7_75t_SL g266 ( 
.A(n_215),
.B(n_196),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_224),
.B(n_167),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_232),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_230),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_212),
.A2(n_206),
.B(n_201),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_232),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_211),
.A2(n_196),
.B1(n_199),
.B2(n_197),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_169),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_173),
.Y(n_276)
);

NAND3xp33_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_194),
.C(n_193),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_238),
.B(n_180),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_238),
.B(n_184),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_223),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_210),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_220),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_219),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_248),
.B(n_246),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_221),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

OR2x6_ASAP7_75t_L g296 ( 
.A(n_217),
.B(n_185),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

NAND2xp33_ASAP7_75t_L g298 ( 
.A(n_220),
.B(n_235),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g299 ( 
.A(n_228),
.B(n_188),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_226),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_237),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_218),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_262),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_249),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_220),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_192),
.B1(n_240),
.B2(n_209),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_240),
.C(n_209),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_214),
.B1(n_266),
.B2(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_294),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_235),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_235),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_236),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_269),
.B(n_247),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_236),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_261),
.B(n_236),
.Y(n_320)
);

AND3x2_ASAP7_75t_SL g321 ( 
.A(n_299),
.B(n_247),
.C(n_245),
.Y(n_321)
);

AND2x2_ASAP7_75t_SL g322 ( 
.A(n_259),
.B(n_214),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_236),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g327 ( 
.A1(n_253),
.A2(n_214),
.B1(n_244),
.B2(n_239),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_261),
.B(n_239),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_266),
.B(n_250),
.C(n_244),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_285),
.B(n_239),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_261),
.B(n_239),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_244),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_258),
.A2(n_250),
.B1(n_244),
.B2(n_233),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_288),
.B(n_250),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_254),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_250),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_297),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g340 ( 
.A1(n_299),
.A2(n_185),
.B1(n_245),
.B2(n_16),
.Y(n_340)
);

NOR3xp33_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_14),
.C(n_15),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_279),
.B(n_14),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_279),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_263),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_288),
.B(n_19),
.Y(n_349)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_277),
.B(n_17),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_286),
.B(n_18),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_270),
.B(n_21),
.Y(n_353)
);

NOR3xp33_ASAP7_75t_L g354 ( 
.A(n_259),
.B(n_22),
.C(n_23),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_286),
.B(n_24),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_287),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_296),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_286),
.B(n_28),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_263),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_296),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_302),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_280),
.B(n_273),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_265),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_298),
.C(n_296),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_305),
.B(n_287),
.Y(n_368)
);

NOR2x1_ASAP7_75t_L g369 ( 
.A(n_329),
.B(n_296),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_271),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_304),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_268),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_313),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_319),
.B(n_268),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_310),
.B(n_273),
.Y(n_379)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_342),
.A2(n_298),
.B(n_291),
.C(n_283),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_307),
.B(n_325),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_320),
.B(n_287),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_325),
.B(n_280),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_327),
.A2(n_291),
.B(n_283),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_301),
.A2(n_29),
.B(n_30),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_311),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_343),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_311),
.A2(n_38),
.B1(n_40),
.B2(n_45),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_334),
.A2(n_46),
.B(n_50),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_152),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_322),
.B(n_51),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_322),
.B(n_52),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_320),
.B(n_328),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_360),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_353),
.A2(n_54),
.B(n_55),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_56),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_353),
.A2(n_57),
.B(n_58),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_351),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_331),
.B(n_65),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_347),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_348),
.Y(n_406)
);

AO22x1_ASAP7_75t_L g407 ( 
.A1(n_341),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_334),
.A2(n_74),
.B(n_75),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_315),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_351),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_331),
.B(n_79),
.Y(n_412)
);

OAI21xp33_ASAP7_75t_L g413 ( 
.A1(n_344),
.A2(n_82),
.B(n_85),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_318),
.B(n_87),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_354),
.B(n_88),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_344),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_352),
.A2(n_92),
.B(n_93),
.C(n_94),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_349),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_356),
.A2(n_316),
.B(n_317),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_324),
.A2(n_103),
.B(n_104),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_300),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

AND2x4_ASAP7_75t_SL g425 ( 
.A(n_340),
.B(n_108),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_336),
.A2(n_109),
.B(n_111),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_362),
.B(n_349),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_381),
.B(n_335),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_323),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_376),
.B(n_340),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_424),
.B(n_333),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_378),
.Y(n_432)
);

AOI221x1_ASAP7_75t_L g433 ( 
.A1(n_395),
.A2(n_396),
.B1(n_389),
.B2(n_387),
.C(n_413),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_358),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_333),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_377),
.A2(n_355),
.B(n_357),
.Y(n_436)
);

OAI21x1_ASAP7_75t_L g437 ( 
.A1(n_365),
.A2(n_114),
.B(n_116),
.Y(n_437)
);

O2A1O1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_416),
.A2(n_357),
.B(n_321),
.C(n_120),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_384),
.A2(n_117),
.B(n_119),
.Y(n_439)
);

NAND2x1_ASAP7_75t_L g440 ( 
.A(n_378),
.B(n_122),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_372),
.B(n_123),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_383),
.A2(n_125),
.B(n_126),
.Y(n_442)
);

INVx4_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_369),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_373),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_321),
.B1(n_128),
.B2(n_129),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_127),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_132),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_L g449 ( 
.A1(n_414),
.A2(n_133),
.B(n_134),
.Y(n_449)
);

AO21x2_ASAP7_75t_L g450 ( 
.A1(n_400),
.A2(n_150),
.B(n_137),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_136),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_380),
.A2(n_138),
.B(n_139),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_404),
.B(n_141),
.C(n_142),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_425),
.B(n_143),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_371),
.B(n_146),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_419),
.A2(n_402),
.B(n_366),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_363),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_392),
.A2(n_148),
.B(n_149),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_382),
.A2(n_394),
.B1(n_367),
.B2(n_388),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_401),
.Y(n_461)
);

AO31x2_ASAP7_75t_L g462 ( 
.A1(n_417),
.A2(n_411),
.A3(n_403),
.B(n_418),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_399),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_386),
.A2(n_375),
.B1(n_406),
.B2(n_397),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_408),
.A2(n_405),
.B(n_393),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_379),
.B(n_368),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_391),
.A2(n_415),
.B(n_422),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_390),
.A2(n_409),
.B(n_385),
.C(n_408),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

O2A1O1Ixp5_ASAP7_75t_L g470 ( 
.A1(n_385),
.A2(n_390),
.B(n_409),
.C(n_420),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_420),
.B(n_426),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_376),
.B(n_326),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_376),
.B(n_326),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_376),
.A2(n_340),
.B1(n_228),
.B2(n_204),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_373),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_376),
.B(n_326),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g477 ( 
.A1(n_383),
.A2(n_381),
.B(n_365),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_472),
.B(n_476),
.Y(n_479)
);

OAI33xp33_ASAP7_75t_L g480 ( 
.A1(n_474),
.A2(n_430),
.A3(n_446),
.B1(n_445),
.B2(n_453),
.B3(n_475),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_465),
.A2(n_477),
.B(n_470),
.Y(n_481)
);

AO21x2_ASAP7_75t_L g482 ( 
.A1(n_457),
.A2(n_436),
.B(n_452),
.Y(n_482)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_433),
.A2(n_435),
.B(n_439),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_444),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_473),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_427),
.A2(n_478),
.B1(n_431),
.B2(n_469),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_458),
.Y(n_487)
);

AND2x6_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_461),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_456),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_437),
.A2(n_468),
.B(n_471),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_460),
.B(n_441),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_429),
.B(n_464),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_447),
.A2(n_448),
.B(n_451),
.Y(n_493)
);

NAND2x1p5_ASAP7_75t_L g494 ( 
.A(n_443),
.B(n_440),
.Y(n_494)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_443),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_428),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_469),
.A2(n_432),
.B1(n_461),
.B2(n_434),
.Y(n_498)
);

OA21x2_ASAP7_75t_L g499 ( 
.A1(n_449),
.A2(n_454),
.B(n_442),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_466),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g501 ( 
.A(n_461),
.Y(n_501)
);

BUFx8_ASAP7_75t_SL g502 ( 
.A(n_438),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_449),
.B(n_462),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g504 ( 
.A(n_450),
.B(n_462),
.Y(n_504)
);

NAND2x1p5_ASAP7_75t_L g505 ( 
.A(n_459),
.B(n_454),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_443),
.B(n_438),
.Y(n_507)
);

A2O1A1Ixp33_ASAP7_75t_L g508 ( 
.A1(n_438),
.A2(n_342),
.B(n_413),
.C(n_425),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

A2O1A1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_438),
.A2(n_342),
.B(n_413),
.C(n_425),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_435),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_430),
.B(n_376),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_443),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_472),
.B(n_376),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_427),
.B(n_362),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_458),
.B(n_364),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_472),
.B(n_376),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_478),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_472),
.B(n_305),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_445),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_516),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_511),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_506),
.A2(n_482),
.B(n_481),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_511),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_515),
.B(n_518),
.Y(n_526)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_484),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_513),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_521),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_485),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

OAI21x1_ASAP7_75t_SL g533 ( 
.A1(n_493),
.A2(n_486),
.B(n_498),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_488),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_492),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_485),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_496),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_509),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_505),
.A2(n_490),
.B(n_494),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_496),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_501),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_488),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_488),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_488),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_479),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

CKINVDCx6p67_ASAP7_75t_R g548 ( 
.A(n_519),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_508),
.A2(n_510),
.B(n_504),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_500),
.B(n_512),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_483),
.A2(n_499),
.B(n_514),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_482),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_507),
.B(n_517),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_517),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_522),
.B(n_510),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_536),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_525),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_508),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_525),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_529),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_531),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_529),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_546),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_523),
.B(n_507),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_532),
.B(n_507),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_499),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_535),
.B(n_499),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_520),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_535),
.B(n_491),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_550),
.B(n_491),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_530),
.B(n_480),
.Y(n_575)
);

INVx1_ASAP7_75t_SL g576 ( 
.A(n_526),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_480),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_552),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_552),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_541),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_526),
.B(n_502),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_495),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_553),
.B(n_495),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_537),
.B(n_495),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_578),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_565),
.B(n_542),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_555),
.B(n_556),
.Y(n_587)
);

CKINVDCx6p67_ASAP7_75t_R g588 ( 
.A(n_558),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_576),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_580),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_580),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_581),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_563),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_L g594 ( 
.A1(n_575),
.A2(n_554),
.B(n_540),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_574),
.B(n_524),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_578),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_574),
.B(n_524),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_565),
.B(n_542),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_568),
.B(n_549),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_549),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_554),
.Y(n_601)
);

AND2x4_ASAP7_75t_SL g602 ( 
.A(n_570),
.B(n_583),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_559),
.Y(n_603)
);

AND2x4_ASAP7_75t_SL g604 ( 
.A(n_570),
.B(n_548),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_559),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_561),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_577),
.B(n_566),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_566),
.B(n_549),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_579),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_555),
.B(n_540),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_571),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_567),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_579),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_551),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_570),
.B(n_537),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_582),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_567),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_561),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_562),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_572),
.B(n_551),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_562),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_595),
.B(n_569),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_595),
.B(n_569),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_597),
.B(n_557),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_585),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_597),
.B(n_557),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_560),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_607),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_619),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_605),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_606),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_607),
.B(n_560),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_585),
.Y(n_634)
);

NAND2x1p5_ASAP7_75t_L g635 ( 
.A(n_614),
.B(n_539),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_593),
.B(n_573),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_618),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_596),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_596),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_609),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_613),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_586),
.B(n_556),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_613),
.Y(n_643)
);

NOR2x1p5_ASAP7_75t_L g644 ( 
.A(n_588),
.B(n_581),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_598),
.B(n_589),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_599),
.B(n_600),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_591),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_634),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_634),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_646),
.B(n_600),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_641),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_646),
.B(n_629),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_629),
.B(n_612),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_625),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_624),
.B(n_617),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_624),
.B(n_626),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_625),
.B(n_612),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_626),
.B(n_617),
.Y(n_659)
);

OR2x2_ASAP7_75t_L g660 ( 
.A(n_622),
.B(n_620),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_645),
.B(n_621),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_627),
.B(n_587),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_640),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_622),
.B(n_620),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_641),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_627),
.B(n_587),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_628),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_661),
.B(n_644),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_662),
.B(n_592),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_649),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_650),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_623),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_623),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_652),
.Y(n_674)
);

OAI222xp33_ASAP7_75t_L g675 ( 
.A1(n_656),
.A2(n_633),
.B1(n_636),
.B2(n_615),
.C1(n_642),
.C2(n_601),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_667),
.A2(n_648),
.B(n_647),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_665),
.Y(n_677)
);

XNOR2x1_ASAP7_75t_L g678 ( 
.A(n_672),
.B(n_611),
.Y(n_678)
);

AOI322xp5_ASAP7_75t_L g679 ( 
.A1(n_668),
.A2(n_657),
.A3(n_633),
.B1(n_664),
.B2(n_654),
.C1(n_651),
.C2(n_659),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_670),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_668),
.A2(n_502),
.B1(n_616),
.B2(n_611),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_671),
.Y(n_682)
);

OAI21xp33_ASAP7_75t_SL g683 ( 
.A1(n_672),
.A2(n_657),
.B(n_654),
.Y(n_683)
);

OAI22xp5_ASAP7_75t_L g684 ( 
.A1(n_669),
.A2(n_660),
.B1(n_666),
.B2(n_588),
.Y(n_684)
);

NOR2x1_ASAP7_75t_L g685 ( 
.A(n_678),
.B(n_675),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_679),
.B(n_673),
.Y(n_686)
);

NOR2x1_ASAP7_75t_L g687 ( 
.A(n_680),
.B(n_674),
.Y(n_687)
);

OAI21xp33_ASAP7_75t_L g688 ( 
.A1(n_681),
.A2(n_676),
.B(n_677),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_684),
.A2(n_604),
.B(n_630),
.Y(n_689)
);

AOI221xp5_ASAP7_75t_L g690 ( 
.A1(n_683),
.A2(n_664),
.B1(n_673),
.B2(n_658),
.C(n_631),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_687),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_685),
.B(n_689),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_688),
.B(n_682),
.C(n_583),
.Y(n_693)
);

NAND4xp75_ASAP7_75t_L g694 ( 
.A(n_686),
.B(n_637),
.C(n_632),
.D(n_582),
.Y(n_694)
);

OAI21xp33_ASAP7_75t_L g695 ( 
.A1(n_692),
.A2(n_690),
.B(n_616),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_691),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_693),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_SL g698 ( 
.A(n_695),
.B(n_697),
.C(n_696),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_696),
.Y(n_699)
);

AND3x2_ASAP7_75t_L g700 ( 
.A(n_696),
.B(n_527),
.C(n_694),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_699),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_698),
.B(n_651),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_700),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_699),
.B(n_604),
.Y(n_704)
);

XNOR2x1_ASAP7_75t_L g705 ( 
.A(n_700),
.B(n_527),
.Y(n_705)
);

OAI221xp5_ASAP7_75t_L g706 ( 
.A1(n_703),
.A2(n_705),
.B1(n_702),
.B2(n_701),
.C(n_704),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_703),
.B(n_584),
.C(n_564),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_701),
.B(n_548),
.Y(n_709)
);

HB1xp67_ASAP7_75t_L g710 ( 
.A(n_702),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_704),
.B(n_658),
.Y(n_711)
);

OA22x2_ASAP7_75t_L g712 ( 
.A1(n_710),
.A2(n_602),
.B1(n_658),
.B2(n_533),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_707),
.Y(n_713)
);

XNOR2x1_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_527),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_711),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_SL g716 ( 
.A1(n_714),
.A2(n_706),
.B(n_709),
.Y(n_716)
);

NAND4xp25_ASAP7_75t_L g717 ( 
.A(n_715),
.B(n_584),
.C(n_594),
.D(n_534),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_713),
.A2(n_663),
.B1(n_655),
.B2(n_635),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_712),
.A2(n_602),
.B1(n_610),
.B2(n_635),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_663),
.B1(n_655),
.B2(n_635),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_718),
.A2(n_643),
.B1(n_639),
.B2(n_638),
.Y(n_721)
);

AOI221xp5_ASAP7_75t_L g722 ( 
.A1(n_716),
.A2(n_533),
.B1(n_544),
.B2(n_547),
.C(n_543),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_722),
.B(n_717),
.Y(n_723)
);

AOI21xp5_ASAP7_75t_L g724 ( 
.A1(n_723),
.A2(n_720),
.B(n_721),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_724),
.B(n_534),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_725),
.A2(n_547),
.B1(n_543),
.B2(n_545),
.Y(n_726)
);


endmodule