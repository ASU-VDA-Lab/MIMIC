module fake_jpeg_10519_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_41),
.B1(n_28),
.B2(n_24),
.Y(n_45)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_50),
.B1(n_33),
.B2(n_1),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_26),
.B1(n_22),
.B2(n_23),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_48),
.B(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_34),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_36),
.A2(n_24),
.B1(n_32),
.B2(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_16),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_56),
.B(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_27),
.B1(n_17),
.B2(n_32),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_78),
.B(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_62),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_65),
.B1(n_70),
.B2(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_20),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_64),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_50),
.A2(n_37),
.B1(n_36),
.B2(n_41),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_75),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_37),
.B(n_18),
.C(n_31),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_2),
.B(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_52),
.B(n_38),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_41),
.B1(n_40),
.B2(n_30),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_41),
.B1(n_40),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_74),
.B1(n_44),
.B2(n_53),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_40),
.B1(n_25),
.B2(n_23),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_22),
.B1(n_19),
.B2(n_18),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_19),
.B1(n_21),
.B2(n_2),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_14),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_81),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_4),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_55),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_87),
.C(n_89),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_54),
.C(n_55),
.Y(n_87)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_95),
.B(n_7),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_100),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_54),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_68),
.B1(n_63),
.B2(n_78),
.Y(n_120)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_102),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_60),
.B(n_5),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_98),
.B(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_109),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_61),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_103),
.Y(n_111)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_112),
.B(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_130),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_121),
.Y(n_139)
);

AO21x2_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_65),
.B(n_83),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_68),
.B1(n_58),
.B2(n_64),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_97),
.B1(n_96),
.B2(n_98),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_128),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_71),
.B1(n_57),
.B2(n_67),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_110),
.A2(n_122),
.B(n_117),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_88),
.B(n_86),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_85),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_137),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_93),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_138),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_147),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_88),
.B1(n_99),
.B2(n_67),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_110),
.B1(n_116),
.B2(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_113),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_152),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_116),
.A2(n_92),
.B1(n_97),
.B2(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_155),
.A2(n_71),
.B1(n_88),
.B2(n_86),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_89),
.B(n_105),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_124),
.B1(n_118),
.B2(n_92),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_159),
.A2(n_161),
.B1(n_140),
.B2(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_152),
.B(n_87),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_139),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_89),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_81),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_165),
.B1(n_135),
.B2(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_135),
.B1(n_155),
.B2(n_150),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_132),
.B(n_75),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_153),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_177),
.B(n_182),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_158),
.B(n_171),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_136),
.C(n_144),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_156),
.C(n_162),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_184),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_134),
.B1(n_143),
.B2(n_137),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_188),
.B(n_166),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_143),
.B1(n_154),
.B2(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_189),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_153),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_173),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_133),
.B1(n_71),
.B2(n_102),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_72),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_197),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_156),
.C(n_166),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_176),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_182),
.B(n_188),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_170),
.C(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_179),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_159),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_201),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_174),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_208),
.C(n_210),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_209),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_179),
.B(n_184),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_185),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_177),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_192),
.C(n_190),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_72),
.C(n_14),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_201),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_214),
.B(n_217),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_199),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_206),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_198),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_222),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_213),
.A2(n_218),
.B1(n_216),
.B2(n_215),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_209),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_223),
.Y(n_224)
);

AOI21x1_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_8),
.B(n_9),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_13),
.C2(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_223),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

OAI321xp33_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_224),
.A3(n_11),
.B1(n_10),
.B2(n_72),
.C(n_225),
.Y(n_230)
);

BUFx24_ASAP7_75t_SL g232 ( 
.A(n_230),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_231),
.Y(n_233)
);

XNOR2x2_ASAP7_75t_SL g234 ( 
.A(n_233),
.B(n_72),
.Y(n_234)
);


endmodule