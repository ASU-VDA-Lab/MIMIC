module fake_jpeg_28076_n_322 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_36),
.B(n_20),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_31),
.Y(n_60)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_32),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_36),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_61),
.B(n_35),
.C(n_34),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_36),
.B(n_40),
.C(n_41),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_40),
.B(n_41),
.C(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_63),
.B(n_78),
.Y(n_132)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_65),
.B(n_40),
.Y(n_116)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_74),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_70),
.B(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_39),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_80),
.Y(n_122)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_48),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_99),
.B1(n_103),
.B2(n_28),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx2_ASAP7_75t_SL g126 ( 
.A(n_79),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_46),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_29),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

OR2x4_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_15),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_92),
.C(n_18),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_38),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_22),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_25),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_25),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_45),
.A2(n_42),
.B1(n_40),
.B2(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_15),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_37),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_18),
.B1(n_24),
.B2(n_42),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_40),
.B1(n_18),
.B2(n_23),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_49),
.B(n_27),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_104),
.A2(n_116),
.B(n_134),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_110),
.A2(n_30),
.B(n_112),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_99),
.B1(n_79),
.B2(n_94),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_129),
.B1(n_73),
.B2(n_98),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_133),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_91),
.A2(n_100),
.B1(n_66),
.B2(n_82),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_64),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_62),
.C(n_65),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_61),
.B(n_65),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_20),
.B(n_26),
.C(n_37),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_135),
.A2(n_154),
.B1(n_35),
.B2(n_34),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_62),
.C(n_68),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_143),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_144),
.A2(n_119),
.B1(n_105),
.B2(n_35),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_92),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_62),
.C(n_73),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_35),
.C(n_33),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_85),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_76),
.B1(n_83),
.B2(n_101),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_162),
.B1(n_93),
.B2(n_34),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_63),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_131),
.A2(n_110),
.B1(n_118),
.B2(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_85),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_30),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_113),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_0),
.B(n_20),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_161),
.B(n_163),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_26),
.B(n_37),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_101),
.B1(n_67),
.B2(n_88),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_93),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_35),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_164),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_176),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_138),
.A2(n_127),
.B(n_117),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_167),
.B(n_172),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_115),
.B(n_125),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_105),
.B1(n_125),
.B2(n_67),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_195),
.B1(n_33),
.B2(n_41),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_115),
.B(n_87),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_140),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_183),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_119),
.B(n_111),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_190),
.B(n_194),
.Y(n_219)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_196),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_185),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_182),
.B1(n_184),
.B2(n_186),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_37),
.C(n_15),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_144),
.A2(n_136),
.B1(n_152),
.B2(n_148),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_145),
.B1(n_143),
.B2(n_155),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_188),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_21),
.B1(n_14),
.B2(n_17),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_21),
.B1(n_14),
.B2(n_17),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_141),
.B(n_34),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_161),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_175),
.B(n_167),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_201),
.B(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_194),
.A2(n_141),
.B1(n_135),
.B2(n_139),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_203),
.A2(n_190),
.B1(n_182),
.B2(n_177),
.Y(n_230)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_206),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_160),
.C(n_34),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_225),
.C(n_183),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_41),
.CI(n_33),
.CON(n_211),
.SN(n_211)
);

NAND2xp33_ASAP7_75t_R g233 ( 
.A(n_211),
.B(n_222),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_21),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_212),
.A2(n_213),
.B1(n_218),
.B2(n_221),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_171),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_178),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_220),
.B(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_169),
.B(n_21),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_172),
.A2(n_41),
.B(n_14),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_41),
.C(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_168),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_189),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_226),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_187),
.C(n_191),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_230),
.A2(n_247),
.B1(n_216),
.B2(n_221),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_191),
.C(n_209),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_219),
.C(n_203),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_241),
.C(n_218),
.Y(n_264)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_204),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_201),
.A2(n_197),
.B1(n_189),
.B2(n_174),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_207),
.B1(n_215),
.B2(n_212),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_174),
.C(n_2),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_1),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_243),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_1),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_216),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_250),
.B(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_262),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_223),
.B1(n_199),
.B2(n_222),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_267),
.B1(n_232),
.B2(n_228),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_207),
.B(n_208),
.Y(n_262)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_264),
.B(n_266),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_211),
.B1(n_4),
.B2(n_5),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_211),
.C(n_4),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_277),
.Y(n_292)
);

BUFx12_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

INVx11_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_242),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_261),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g280 ( 
.A(n_261),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_284),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_257),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_264),
.C(n_266),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_288),
.C(n_296),
.Y(n_304)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_248),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_293),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_256),
.B(n_227),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_294),
.B(n_295),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_268),
.B(n_252),
.Y(n_293)
);

A2O1A1Ixp33_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_260),
.B(n_254),
.C(n_259),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_267),
.B(n_245),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_235),
.C(n_263),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_275),
.B1(n_279),
.B2(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_300),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_244),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_277),
.C(n_278),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_302),
.C(n_305),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_270),
.C(n_274),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_291),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_5),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_289),
.B(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_294),
.B(n_293),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_294),
.C(n_8),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_8),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_301),
.C(n_302),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_314),
.C(n_307),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_315),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_8),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_9),
.Y(n_322)
);


endmodule