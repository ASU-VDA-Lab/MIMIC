module fake_jpeg_449_n_51 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_51);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_51;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_SL g7 ( 
.A(n_6),
.Y(n_7)
);

BUFx4f_ASAP7_75t_SL g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_20),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_11),
.A2(n_4),
.B1(n_0),
.B2(n_1),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_22),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_21),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_9),
.Y(n_23)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_16),
.B1(n_10),
.B2(n_8),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_26),
.Y(n_28)
);

CKINVDCx9p33_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_25),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_22),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_18),
.B1(n_13),
.B2(n_21),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_20),
.C(n_23),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_26),
.C(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_10),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_41),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_30),
.Y(n_43)
);

AOI322xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_14),
.A3(n_28),
.B1(n_8),
.B2(n_27),
.C1(n_15),
.C2(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_15),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_44),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_43),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_49),
.A2(n_48),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_17),
.Y(n_51)
);


endmodule