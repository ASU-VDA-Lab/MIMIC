module fake_ariane_199_n_751 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_751);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_751;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_670;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_151;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

BUFx3_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_52),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_21),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_2),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_133),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_44),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_30),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_6),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_31),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_77),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_15),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_2),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_131),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_20),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_86),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_78),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_67),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_139),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_53),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_73),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_108),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_23),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_14),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_13),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_8),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_97),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_45),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_35),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_122),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_153),
.B(n_191),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_0),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_148),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_174),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_165),
.B(n_0),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_1),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_151),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_19),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_200),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_1),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_178),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_172),
.B(n_3),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_182),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_22),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_186),
.B(n_197),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_195),
.B(n_3),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_154),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_198),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

BUFx6f_ASAP7_75t_SL g249 ( 
.A(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_220),
.B(n_157),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_224),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_202),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_205),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

NAND2xp33_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_158),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_220),
.B(n_164),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_210),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_228),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_201),
.B(n_199),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_207),
.B(n_212),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_218),
.B(n_166),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_169),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_209),
.B(n_177),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_204),
.B(n_183),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g275 ( 
.A(n_221),
.B(n_152),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

AND3x2_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_196),
.C(n_189),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_203),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_203),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_223),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_237),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_207),
.B(n_187),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_217),
.B(n_152),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_237),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_207),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_207),
.B(n_190),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_4),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_206),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

AND2x4_ASAP7_75t_L g297 ( 
.A(n_254),
.B(n_218),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_222),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_253),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_247),
.A2(n_243),
.B1(n_219),
.B2(n_241),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_247),
.B(n_207),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_218),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_219),
.C(n_236),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_222),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_247),
.B(n_212),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_231),
.C(n_245),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_254),
.B(n_212),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_280),
.Y(n_309)
);

OR2x4_ASAP7_75t_L g310 ( 
.A(n_293),
.B(n_208),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_247),
.A2(n_243),
.B1(n_241),
.B2(n_240),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_285),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_247),
.B(n_212),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_212),
.Y(n_316)
);

AOI22x1_ASAP7_75t_L g317 ( 
.A1(n_252),
.A2(n_243),
.B1(n_269),
.B2(n_274),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_251),
.A2(n_217),
.B1(n_189),
.B2(n_196),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_251),
.B(n_222),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_262),
.B(n_217),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_211),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g324 ( 
.A1(n_261),
.A2(n_272),
.B(n_273),
.C(n_278),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_261),
.B(n_235),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_272),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_260),
.B(n_246),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_275),
.A2(n_156),
.B1(n_176),
.B2(n_185),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_277),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_290),
.B(n_246),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_265),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_270),
.B(n_246),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_246),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_275),
.A2(n_156),
.B1(n_240),
.B2(n_235),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_258),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_249),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_259),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_216),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_249),
.A2(n_241),
.B1(n_239),
.B2(n_238),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_233),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_282),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_279),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_270),
.B(n_230),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_294),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_252),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_279),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_271),
.A2(n_295),
.B1(n_281),
.B2(n_233),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_233),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_292),
.A2(n_216),
.B(n_229),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_324),
.A2(n_292),
.B(n_264),
.Y(n_357)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_298),
.B(n_267),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_305),
.B(n_270),
.Y(n_360)
);

A2O1A1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_303),
.A2(n_232),
.B(n_213),
.C(n_208),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_302),
.A2(n_276),
.B(n_270),
.Y(n_362)
);

NAND2x1p5_ASAP7_75t_L g363 ( 
.A(n_299),
.B(n_285),
.Y(n_363)
);

AOI21x1_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_274),
.B(n_232),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_353),
.B(n_285),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_300),
.B(n_270),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_276),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_356),
.A2(n_276),
.B(n_225),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_307),
.A2(n_213),
.B1(n_225),
.B2(n_276),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_340),
.B(n_276),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_318),
.B(n_4),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_319),
.A2(n_326),
.B(n_349),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_309),
.B(n_5),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_225),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_329),
.Y(n_375)
);

OR2x6_ASAP7_75t_SL g376 ( 
.A(n_330),
.B(n_337),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_225),
.B(n_69),
.Y(n_378)
);

OAI21xp33_ASAP7_75t_L g379 ( 
.A1(n_296),
.A2(n_5),
.B(n_6),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_297),
.B(n_7),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_312),
.A2(n_72),
.B(n_145),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_7),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_304),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_297),
.B(n_10),
.Y(n_384)
);

O2A1O1Ixp5_ASAP7_75t_L g385 ( 
.A1(n_311),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_325),
.B(n_11),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_325),
.B(n_12),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_316),
.B(n_14),
.Y(n_388)
);

O2A1O1Ixp5_ASAP7_75t_L g389 ( 
.A1(n_313),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_310),
.B(n_16),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_18),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_328),
.B(n_18),
.Y(n_394)
);

O2A1O1Ixp33_ASAP7_75t_L g395 ( 
.A1(n_348),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_395)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_336),
.A2(n_27),
.B(n_28),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_334),
.A2(n_32),
.B(n_33),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_310),
.Y(n_399)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_314),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_338),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_331),
.B(n_38),
.Y(n_402)
);

BUFx8_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_320),
.B(n_146),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_352),
.A2(n_39),
.B(n_40),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_344),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_322),
.A2(n_46),
.B(n_47),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_333),
.A2(n_48),
.B(n_49),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_343),
.B(n_50),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_327),
.Y(n_412)
);

NOR3xp33_ASAP7_75t_L g413 ( 
.A(n_332),
.B(n_347),
.C(n_346),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_345),
.A2(n_54),
.B(n_56),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_354),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_415)
);

OAI21x1_ASAP7_75t_L g416 ( 
.A1(n_317),
.A2(n_61),
.B(n_62),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_301),
.A2(n_63),
.B(n_64),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_301),
.B(n_143),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_306),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_418),
.A2(n_416),
.B(n_368),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_399),
.B(n_314),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_359),
.A2(n_315),
.B(n_308),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_412),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_375),
.Y(n_424)
);

A2O1A1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_371),
.A2(n_355),
.B(n_79),
.C(n_81),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_361),
.A2(n_75),
.B(n_82),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_381),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_90),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_403),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_372),
.A2(n_91),
.B(n_93),
.Y(n_430)
);

BUFx4f_ASAP7_75t_SL g431 ( 
.A(n_403),
.Y(n_431)
);

A2O1A1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_379),
.A2(n_95),
.B(n_96),
.C(n_99),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_367),
.A2(n_100),
.B(n_101),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_366),
.A2(n_105),
.B(n_109),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_110),
.Y(n_435)
);

AO31x2_ASAP7_75t_L g436 ( 
.A1(n_396),
.A2(n_111),
.A3(n_112),
.B(n_113),
.Y(n_436)
);

AOI21x1_ASAP7_75t_L g437 ( 
.A1(n_360),
.A2(n_115),
.B(n_117),
.Y(n_437)
);

AO21x2_ASAP7_75t_L g438 ( 
.A1(n_357),
.A2(n_118),
.B(n_119),
.Y(n_438)
);

OAI21x1_ASAP7_75t_L g439 ( 
.A1(n_364),
.A2(n_120),
.B(n_121),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_386),
.A2(n_123),
.B(n_124),
.C(n_125),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_374),
.A2(n_127),
.B(n_128),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_377),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_365),
.A2(n_129),
.B(n_130),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_378),
.A2(n_132),
.B(n_134),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_388),
.B(n_135),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_402),
.B(n_136),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_385),
.A2(n_137),
.B(n_138),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_400),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_387),
.B(n_142),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_413),
.B(n_394),
.C(n_383),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_388),
.B(n_398),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_376),
.B(n_384),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_362),
.A2(n_417),
.B(n_405),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_414),
.A2(n_407),
.B(n_408),
.Y(n_457)
);

O2A1O1Ixp5_ASAP7_75t_L g458 ( 
.A1(n_393),
.A2(n_410),
.B(n_404),
.C(n_380),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_377),
.B(n_406),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_409),
.A2(n_406),
.B(n_397),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_400),
.A2(n_395),
.B(n_358),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_370),
.B(n_369),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_419),
.A2(n_415),
.B(n_389),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_358),
.B(n_392),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_401),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_323),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_388),
.B(n_337),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_359),
.A2(n_367),
.B(n_372),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_359),
.A2(n_367),
.B(n_372),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_416),
.B(n_368),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_391),
.B(n_298),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_359),
.A2(n_367),
.B(n_372),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_361),
.A2(n_372),
.B(n_378),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_423),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_471),
.B(n_467),
.Y(n_477)
);

CKINVDCx11_ASAP7_75t_R g478 ( 
.A(n_424),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_429),
.Y(n_479)
);

INVx3_ASAP7_75t_SL g480 ( 
.A(n_466),
.Y(n_480)
);

OAI21x1_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_456),
.B(n_420),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

OA21x2_ASAP7_75t_L g483 ( 
.A1(n_470),
.A2(n_473),
.B(n_469),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_454),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_464),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_455),
.B(n_475),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_441),
.C(n_426),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_444),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_457),
.A2(n_472),
.B(n_468),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_464),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_465),
.B(n_458),
.Y(n_492)
);

OR3x4_ASAP7_75t_SL g493 ( 
.A(n_431),
.B(n_435),
.C(n_448),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_448),
.A2(n_427),
.B1(n_453),
.B2(n_426),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_449),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_421),
.B(n_447),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_421),
.B(n_451),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_451),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_473),
.A2(n_422),
.B(n_463),
.Y(n_499)
);

AO31x2_ASAP7_75t_L g500 ( 
.A1(n_427),
.A2(n_432),
.A3(n_425),
.B(n_452),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_428),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_459),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_461),
.A2(n_430),
.B(n_450),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_450),
.B(n_430),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_438),
.A2(n_434),
.B1(n_440),
.B2(n_445),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_438),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_439),
.A2(n_446),
.B(n_442),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_433),
.B(n_437),
.Y(n_509)
);

AO31x2_ASAP7_75t_L g510 ( 
.A1(n_436),
.A2(n_427),
.A3(n_469),
.B(n_468),
.Y(n_510)
);

OA21x2_ASAP7_75t_L g511 ( 
.A1(n_436),
.A2(n_470),
.B(n_420),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_436),
.A2(n_359),
.B(n_468),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_467),
.A2(n_371),
.B1(n_455),
.B2(n_275),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_424),
.B(n_329),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_376),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_454),
.Y(n_516)
);

NAND2x1p5_ASAP7_75t_L g517 ( 
.A(n_464),
.B(n_451),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_423),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_454),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_420),
.A2(n_470),
.B(n_357),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_424),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_513),
.A2(n_515),
.B1(n_507),
.B2(n_494),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_485),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_488),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

AO21x2_ASAP7_75t_L g527 ( 
.A1(n_504),
.A2(n_505),
.B(n_512),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_476),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_482),
.Y(n_529)
);

AO21x2_ASAP7_75t_L g530 ( 
.A1(n_505),
.A2(n_499),
.B(n_506),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_519),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_501),
.B(n_520),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_513),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_501),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_519),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_495),
.Y(n_537)
);

BUFx4f_ASAP7_75t_SL g538 ( 
.A(n_522),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_481),
.A2(n_490),
.B(n_508),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_477),
.B(n_480),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_494),
.A2(n_487),
.B(n_492),
.Y(n_541)
);

NOR2x1_ASAP7_75t_SL g542 ( 
.A(n_492),
.B(n_521),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_491),
.B(n_480),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_491),
.B(n_520),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_514),
.Y(n_545)
);

BUFx4f_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

BUFx5_ASAP7_75t_L g547 ( 
.A(n_496),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_483),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_483),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_485),
.B(n_520),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_478),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_521),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_511),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_520),
.B(n_517),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_484),
.Y(n_558)
);

INVxp33_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_555),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_530),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_538),
.B(n_502),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_511),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_555),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_556),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_533),
.B(n_500),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_529),
.B(n_500),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_556),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_534),
.B(n_497),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_540),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_526),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_526),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_529),
.B(n_500),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_530),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_536),
.B(n_500),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_540),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_532),
.B(n_498),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_554),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_525),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_554),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_536),
.B(n_503),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_479),
.Y(n_585)
);

BUFx2_ASAP7_75t_SL g586 ( 
.A(n_547),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_541),
.B(n_493),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_547),
.B(n_508),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_547),
.B(n_508),
.Y(n_589)
);

NOR2x1_ASAP7_75t_L g590 ( 
.A(n_534),
.B(n_509),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_532),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_546),
.A2(n_523),
.B1(n_545),
.B2(n_547),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_547),
.B(n_546),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_547),
.B(n_546),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_547),
.B(n_528),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_548),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_548),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_552),
.B(n_544),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_551),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_524),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_549),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_562),
.B(n_559),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_571),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_563),
.B(n_527),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_581),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_581),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_572),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_573),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_583),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_574),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_588),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_531),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_601),
.B(n_553),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_580),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_578),
.B(n_553),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_587),
.B(n_535),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_563),
.B(n_567),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_567),
.B(n_527),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_568),
.B(n_527),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_568),
.B(n_542),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_574),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_575),
.B(n_542),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_564),
.B(n_576),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_552),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_575),
.B(n_551),
.Y(n_627)
);

AOI221xp5_ASAP7_75t_L g628 ( 
.A1(n_576),
.A2(n_550),
.B1(n_543),
.B2(n_544),
.C(n_537),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_579),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_577),
.B(n_543),
.Y(n_630)
);

NAND2x1p5_ASAP7_75t_L g631 ( 
.A(n_580),
.B(n_593),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_598),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_584),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_600),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_560),
.B(n_539),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_598),
.B(n_539),
.Y(n_636)
);

NOR2x1_ASAP7_75t_L g637 ( 
.A(n_616),
.B(n_590),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_605),
.Y(n_638)
);

NAND2x1p5_ASAP7_75t_L g639 ( 
.A(n_634),
.B(n_600),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_618),
.B(n_588),
.Y(n_640)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_603),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_605),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_632),
.B(n_569),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_606),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_633),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_618),
.B(n_612),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_606),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_612),
.B(n_589),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_579),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_608),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_580),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_624),
.B(n_586),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_636),
.B(n_589),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_608),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_636),
.B(n_561),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_SL g656 ( 
.A(n_604),
.B(n_590),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_629),
.B(n_580),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_604),
.B(n_561),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_610),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_630),
.B(n_561),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_630),
.B(n_619),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_617),
.B(n_619),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_627),
.B(n_570),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_627),
.Y(n_665)
);

AND2x2_ASAP7_75t_SL g666 ( 
.A(n_624),
.B(n_591),
.Y(n_666)
);

AND2x4_ASAP7_75t_SL g667 ( 
.A(n_652),
.B(n_625),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_641),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_646),
.B(n_625),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_665),
.B(n_662),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_662),
.B(n_620),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_645),
.B(n_620),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_646),
.B(n_625),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_637),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_638),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_640),
.B(n_623),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_640),
.B(n_623),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_649),
.B(n_614),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_643),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_642),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_647),
.Y(n_682)
);

INVxp33_ASAP7_75t_L g683 ( 
.A(n_649),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_652),
.B(n_621),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_650),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_654),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_659),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_653),
.B(n_648),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_664),
.B(n_621),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_686),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_683),
.A2(n_592),
.B1(n_652),
.B2(n_666),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_668),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_686),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_675),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_669),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_678),
.A2(n_584),
.B1(n_594),
.B2(n_593),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_683),
.A2(n_652),
.B1(n_666),
.B2(n_657),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_668),
.B(n_661),
.C(n_655),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_674),
.B(n_663),
.Y(n_699)
);

INVx1_ASAP7_75t_SL g700 ( 
.A(n_672),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_692),
.B(n_679),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_L g702 ( 
.A1(n_698),
.A2(n_678),
.B(n_689),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_L g703 ( 
.A(n_690),
.B(n_670),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_699),
.A2(n_667),
.B(n_602),
.C(n_671),
.Y(n_704)
);

OAI21xp33_ASAP7_75t_L g705 ( 
.A1(n_693),
.A2(n_681),
.B(n_687),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_694),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_695),
.B(n_667),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_SL g708 ( 
.A1(n_702),
.A2(n_691),
.B(n_696),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_704),
.A2(n_696),
.B1(n_697),
.B2(n_684),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_706),
.A2(n_700),
.B1(n_658),
.B2(n_628),
.Y(n_710)
);

OAI322xp33_ASAP7_75t_L g711 ( 
.A1(n_701),
.A2(n_685),
.A3(n_682),
.B1(n_680),
.B2(n_677),
.C1(n_676),
.C2(n_673),
.Y(n_711)
);

AOI211xp5_ASAP7_75t_L g712 ( 
.A1(n_703),
.A2(n_684),
.B(n_648),
.C(n_655),
.Y(n_712)
);

AOI211xp5_ASAP7_75t_SL g713 ( 
.A1(n_705),
.A2(n_657),
.B(n_651),
.C(n_615),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_707),
.A2(n_585),
.B(n_688),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_711),
.Y(n_715)
);

NOR4xp75_ASAP7_75t_L g716 ( 
.A(n_709),
.B(n_653),
.C(n_615),
.D(n_660),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_708),
.B(n_660),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_714),
.A2(n_594),
.B(n_657),
.Y(n_718)
);

NOR3xp33_ASAP7_75t_L g719 ( 
.A(n_715),
.B(n_712),
.C(n_713),
.Y(n_719)
);

AOI211xp5_ASAP7_75t_L g720 ( 
.A1(n_717),
.A2(n_651),
.B(n_710),
.C(n_579),
.Y(n_720)
);

NOR4xp25_ASAP7_75t_L g721 ( 
.A(n_716),
.B(n_570),
.C(n_635),
.D(n_569),
.Y(n_721)
);

NAND2x1p5_ASAP7_75t_L g722 ( 
.A(n_721),
.B(n_718),
.Y(n_722)
);

NOR3xp33_ASAP7_75t_L g723 ( 
.A(n_719),
.B(n_600),
.C(n_579),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_720),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_721),
.B(n_658),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_725),
.B(n_656),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_724),
.Y(n_727)
);

INVxp33_ASAP7_75t_L g728 ( 
.A(n_723),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_722),
.Y(n_729)
);

AND2x2_ASAP7_75t_SL g730 ( 
.A(n_723),
.B(n_600),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_722),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_729),
.B(n_639),
.Y(n_732)
);

XNOR2x1_ASAP7_75t_L g733 ( 
.A(n_731),
.B(n_727),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_727),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_728),
.B(n_656),
.Y(n_735)
);

OAI222xp33_ASAP7_75t_L g736 ( 
.A1(n_726),
.A2(n_609),
.B1(n_607),
.B2(n_611),
.C1(n_622),
.C2(n_626),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_733),
.A2(n_730),
.B1(n_586),
.B2(n_651),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_734),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_735),
.Y(n_739)
);

OAI322xp33_ASAP7_75t_L g740 ( 
.A1(n_732),
.A2(n_635),
.A3(n_566),
.B1(n_565),
.B2(n_560),
.C1(n_597),
.C2(n_599),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_738),
.A2(n_736),
.B1(n_639),
.B2(n_634),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_739),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_740),
.A2(n_582),
.B1(n_537),
.B2(n_595),
.Y(n_743)
);

OAI321xp33_ASAP7_75t_L g744 ( 
.A1(n_741),
.A2(n_737),
.A3(n_524),
.B1(n_557),
.B2(n_631),
.C(n_565),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_742),
.A2(n_634),
.B1(n_566),
.B2(n_631),
.Y(n_745)
);

NAND3x2_ASAP7_75t_L g746 ( 
.A(n_743),
.B(n_597),
.C(n_599),
.Y(n_746)
);

NOR2x1_ASAP7_75t_SL g747 ( 
.A(n_745),
.B(n_634),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_744),
.B(n_634),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_747),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_749),
.B(n_748),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_750),
.A2(n_746),
.B(n_596),
.Y(n_751)
);


endmodule