module fake_netlist_5_196_n_41 (n_8, n_4, n_5, n_7, n_0, n_2, n_3, n_6, n_1, n_41);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_2;
input n_3;
input n_6;
input n_1;

output n_41;

wire n_29;
wire n_16;
wire n_12;
wire n_9;
wire n_36;
wire n_25;
wire n_18;
wire n_27;
wire n_22;
wire n_10;
wire n_24;
wire n_28;
wire n_21;
wire n_40;
wire n_34;
wire n_38;
wire n_35;
wire n_32;
wire n_11;
wire n_17;
wire n_19;
wire n_37;
wire n_15;
wire n_26;
wire n_30;
wire n_20;
wire n_33;
wire n_14;
wire n_31;
wire n_23;
wire n_13;
wire n_39;

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_0),
.Y(n_12)
);

OAI21x1_ASAP7_75t_L g13 ( 
.A1(n_8),
.A2(n_2),
.B(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

XNOR2x2_ASAP7_75t_SL g16 ( 
.A(n_15),
.B(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_R g23 ( 
.A(n_10),
.B(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_9),
.B1(n_15),
.B2(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

OAI31xp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_18),
.A3(n_20),
.B(n_22),
.Y(n_27)
);

OAI33xp33_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_22),
.A3(n_20),
.B1(n_23),
.B2(n_16),
.B3(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_13),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_21),
.B1(n_7),
.B2(n_8),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_24),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR3xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.C(n_31),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_32),
.Y(n_37)
);

NOR3xp33_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_27),
.C(n_34),
.Y(n_38)
);

INVxp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_7),
.A3(n_32),
.B1(n_38),
.B2(n_39),
.C1(n_19),
.C2(n_21),
.Y(n_41)
);


endmodule