module fake_ariane_1927_n_1724 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1724);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1724;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_66),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_108),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_83),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_21),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_19),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_40),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_91),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_5),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_76),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_111),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_37),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_89),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_95),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_45),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_42),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_105),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_52),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_137),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_147),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_100),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_32),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_64),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_51),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_37),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_90),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_23),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_77),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_73),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_63),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_54),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_16),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_96),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_92),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_68),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_46),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_22),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_88),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_45),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_38),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_9),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_27),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_41),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_18),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_30),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_11),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_124),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_62),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_43),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_72),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_51),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_1),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_87),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_41),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_2),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_122),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_31),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_145),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_30),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_47),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_38),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_110),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_4),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_33),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_4),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_14),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_17),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_118),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_78),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_58),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_27),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_146),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_67),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_48),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_46),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_40),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_39),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_69),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_94),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_52),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_113),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_149),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_107),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_48),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_57),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_16),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_132),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_19),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_133),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_85),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_47),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_18),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_82),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_115),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_103),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_6),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_29),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_130),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_127),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_140),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_93),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_138),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_135),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_125),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_7),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_75),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_53),
.Y(n_278)
);

BUFx10_ASAP7_75t_L g279 ( 
.A(n_20),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_99),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_7),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_49),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_71),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_104),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_109),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_20),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_25),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_8),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_58),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_65),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_81),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_1),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_35),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_79),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_86),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_28),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_150),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

BUFx2_ASAP7_75t_SL g302 ( 
.A(n_173),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_243),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_175),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_226),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_185),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_207),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_190),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_253),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_227),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_156),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_155),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_254),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_159),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_162),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_230),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_231),
.B(n_0),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_165),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_166),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_254),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_232),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_163),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_170),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_163),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_178),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_172),
.B(n_180),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_172),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_156),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_180),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_191),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_193),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_198),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_241),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_169),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_278),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_226),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_199),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_184),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_202),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_205),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_187),
.B(n_2),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_187),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_206),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_192),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_209),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_192),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_197),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_161),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_197),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_182),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_204),
.B(n_3),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_161),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_218),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_204),
.Y(n_363)
);

INVxp33_ASAP7_75t_L g364 ( 
.A(n_169),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_284),
.B(n_3),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_188),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_219),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_183),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_213),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_221),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_222),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_203),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_331),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_327),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_333),
.B(n_213),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_216),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_301),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_183),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_303),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_216),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_304),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_215),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_211),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_234),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_316),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_318),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_338),
.B(n_234),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_338),
.B(n_215),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_307),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_307),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_325),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_211),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_223),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_358),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_182),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_352),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_354),
.A2(n_252),
.B(n_225),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_354),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_355),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_355),
.B(n_176),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_306),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_357),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_369),
.B(n_182),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_203),
.Y(n_426)
);

INVx5_ASAP7_75t_L g427 ( 
.A(n_302),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_315),
.B(n_182),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_302),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_344),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_315),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_317),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_385),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_382),
.B(n_223),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_319),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_436),
.A2(n_309),
.B1(n_323),
.B2(n_335),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_385),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_420),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_400),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_321),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_436),
.A2(n_323),
.B1(n_342),
.B2(n_366),
.Y(n_455)
);

NOR2x1p5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_311),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_385),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_420),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_420),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_420),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_429),
.A2(n_312),
.B1(n_276),
.B2(n_262),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_422),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_382),
.B(n_324),
.Y(n_463)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_422),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_382),
.A2(n_356),
.B1(n_361),
.B2(n_368),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_422),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_427),
.B(n_326),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_402),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_436),
.A2(n_245),
.B1(n_249),
.B2(n_255),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_435),
.B(n_330),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_332),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_390),
.B(n_342),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_401),
.B(n_403),
.Y(n_473)
);

NAND3xp33_ASAP7_75t_L g474 ( 
.A(n_436),
.B(n_200),
.C(n_182),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_337),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_402),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_401),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_339),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_385),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_422),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_422),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_436),
.A2(n_366),
.B1(n_269),
.B2(n_266),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_422),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_402),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_373),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_403),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_427),
.B(n_340),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_422),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_435),
.B(n_266),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_436),
.A2(n_269),
.B1(n_282),
.B2(n_188),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_402),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_419),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_422),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

OAI21xp33_ASAP7_75t_SL g498 ( 
.A1(n_432),
.A2(n_228),
.B(n_210),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_387),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_402),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_387),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_435),
.B(n_345),
.Y(n_502)
);

AND2x6_ASAP7_75t_L g503 ( 
.A(n_390),
.B(n_225),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_347),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_427),
.B(n_348),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_427),
.B(n_351),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_390),
.B(n_353),
.Y(n_507)
);

INVxp33_ASAP7_75t_SL g508 ( 
.A(n_419),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_383),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_437),
.B(n_359),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_390),
.A2(n_157),
.B1(n_261),
.B2(n_287),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_406),
.B(n_210),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_427),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_437),
.B(n_362),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_389),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_375),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_375),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_413),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_413),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_402),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_389),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_437),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_389),
.Y(n_527)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_389),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_406),
.A2(n_267),
.B1(n_256),
.B2(n_244),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_375),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_373),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_437),
.B(n_367),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_394),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_437),
.B(n_370),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_427),
.B(n_371),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_426),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_388),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_434),
.B(n_220),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_415),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_406),
.B(n_260),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_437),
.B(n_240),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_388),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_434),
.B(n_265),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_427),
.B(n_181),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_394),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_427),
.B(n_181),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_406),
.B(n_224),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_394),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_376),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_374),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_415),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_426),
.B(n_425),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_376),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_437),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_437),
.B(n_275),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_437),
.B(n_277),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_426),
.B(n_181),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_437),
.B(n_260),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_375),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_425),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_376),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_376),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_377),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_377),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_374),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_377),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_426),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_433),
.A2(n_282),
.B1(n_281),
.B2(n_299),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_388),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_388),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_374),
.B(n_181),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_425),
.B(n_228),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_425),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_377),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_374),
.B(n_208),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_418),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_433),
.B(n_176),
.Y(n_581)
);

NAND2xp33_ASAP7_75t_L g582 ( 
.A(n_433),
.B(n_152),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_433),
.B(n_432),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_432),
.A2(n_258),
.B1(n_233),
.B2(n_299),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_428),
.A2(n_258),
.B1(n_233),
.B2(n_281),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_447),
.A2(n_374),
.B1(n_378),
.B2(n_428),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_470),
.B(n_478),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_553),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_502),
.B(n_428),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_510),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_510),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_447),
.A2(n_374),
.B1(n_378),
.B2(n_428),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_374),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_448),
.B(n_428),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_540),
.B(n_428),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_522),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_545),
.B(n_428),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_558),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_447),
.B(n_416),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_447),
.B(n_416),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_447),
.B(n_416),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_517),
.B(n_553),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_522),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_523),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_447),
.B(n_416),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_553),
.B(n_379),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_447),
.B(n_430),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_557),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_581),
.A2(n_418),
.B1(n_386),
.B2(n_407),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_430),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_553),
.B(n_379),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_508),
.B(n_495),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_503),
.B(n_430),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_503),
.B(n_430),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_472),
.B(n_379),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_468),
.B(n_412),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_523),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_517),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_473),
.B(n_379),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_517),
.B(n_379),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_538),
.B(n_308),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_517),
.B(n_379),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_565),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_571),
.B(n_310),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_569),
.Y(n_627)
);

O2A1O1Ixp5_ASAP7_75t_L g628 ( 
.A1(n_438),
.A2(n_392),
.B(n_380),
.C(n_399),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_503),
.B(n_542),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_463),
.B(n_507),
.C(n_495),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_503),
.A2(n_379),
.B1(n_384),
.B2(n_391),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_473),
.B(n_384),
.Y(n_632)
);

NOR2x1p5_ASAP7_75t_L g633 ( 
.A(n_507),
.B(n_386),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_569),
.B(n_384),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_520),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_534),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_446),
.B(n_314),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_503),
.B(n_388),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_558),
.A2(n_407),
.B1(n_397),
.B2(n_412),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_503),
.B(n_388),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_542),
.B(n_384),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_534),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_542),
.B(n_384),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_520),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_569),
.B(n_384),
.Y(n_645)
);

NOR2xp67_ASAP7_75t_L g646 ( 
.A(n_468),
.B(n_412),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_542),
.B(n_384),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_565),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_R g649 ( 
.A(n_550),
.B(n_322),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_542),
.B(n_583),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_542),
.B(n_391),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_542),
.B(n_391),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_453),
.B(n_328),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_564),
.B(n_391),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_566),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_541),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_497),
.B(n_341),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_567),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_498),
.A2(n_424),
.B1(n_421),
.B2(n_412),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_564),
.B(n_391),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_526),
.B(n_380),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_456),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_477),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_530),
.B(n_513),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_577),
.B(n_391),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_577),
.B(n_391),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_567),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_515),
.A2(n_396),
.B1(n_417),
.B2(n_423),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_508),
.B(n_343),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_568),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_455),
.B(n_396),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_477),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_456),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_561),
.B(n_396),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_560),
.B(n_396),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_561),
.B(n_396),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_556),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_575),
.B(n_396),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_489),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_575),
.B(n_396),
.Y(n_683)
);

O2A1O1Ixp5_ASAP7_75t_L g684 ( 
.A1(n_454),
.A2(n_395),
.B(n_380),
.C(n_381),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_471),
.A2(n_392),
.B(n_381),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_489),
.B(n_288),
.C(n_286),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_450),
.B(n_381),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_475),
.B(n_392),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_556),
.B(n_305),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_554),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_570),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_512),
.B(n_393),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_530),
.B(n_397),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_518),
.B(n_533),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_514),
.B(n_393),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_536),
.B(n_393),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_543),
.B(n_395),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_513),
.B(n_421),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_514),
.Y(n_700)
);

AOI22xp5_ASAP7_75t_L g701 ( 
.A1(n_498),
.A2(n_424),
.B1(n_421),
.B2(n_423),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_476),
.B(n_421),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_465),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_461),
.B(n_395),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_559),
.B(n_399),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_515),
.A2(n_424),
.B1(n_423),
.B2(n_411),
.Y(n_706)
);

NAND2x1_ASAP7_75t_L g707 ( 
.A(n_539),
.B(n_544),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_439),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_570),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_578),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_526),
.B(n_399),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_439),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_487),
.B(n_405),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_SL g714 ( 
.A(n_476),
.B(n_173),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_579),
.B(n_405),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_555),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_485),
.B(n_173),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_515),
.B(n_405),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_485),
.B(n_424),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_492),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_487),
.B(n_417),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_494),
.B(n_417),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_578),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_444),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_444),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_494),
.B(n_411),
.Y(n_726)
);

O2A1O1Ixp5_ASAP7_75t_L g727 ( 
.A1(n_546),
.A2(n_423),
.B(n_411),
.C(n_264),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_539),
.A2(n_414),
.B(n_423),
.C(n_411),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_515),
.B(n_398),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_492),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_451),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_515),
.A2(n_423),
.B1(n_411),
.B2(n_173),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_451),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_L g734 ( 
.A(n_520),
.B(n_383),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_492),
.B(n_411),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_457),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_576),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_457),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_492),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_532),
.B(n_411),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_532),
.B(n_423),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_539),
.B(n_375),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_544),
.B(n_375),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_544),
.B(n_398),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_479),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_573),
.B(n_375),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_573),
.B(n_375),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_492),
.B(n_414),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_479),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_500),
.B(n_208),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_480),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_480),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_573),
.B(n_398),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_500),
.B(n_208),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_574),
.B(n_398),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_520),
.Y(n_756)
);

O2A1O1Ixp33_ASAP7_75t_L g757 ( 
.A1(n_587),
.A2(n_582),
.B(n_469),
.C(n_555),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_483),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_593),
.B(n_585),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_666),
.A2(n_580),
.B1(n_549),
.B2(n_572),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_586),
.A2(n_574),
.B1(n_580),
.B2(n_528),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_633),
.A2(n_584),
.B1(n_524),
.B2(n_504),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_588),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_680),
.B(n_574),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_696),
.B(n_576),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_588),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_590),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_680),
.B(n_493),
.Y(n_768)
);

AO21x1_ASAP7_75t_L g769 ( 
.A1(n_695),
.A2(n_562),
.B(n_490),
.Y(n_769)
);

A2O1A1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_704),
.A2(n_414),
.B(n_551),
.C(n_548),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_588),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_737),
.B(n_524),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_617),
.B(n_486),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_665),
.B(n_288),
.C(n_286),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_208),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_700),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_637),
.B(n_474),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_688),
.A2(n_697),
.B(n_693),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_742),
.A2(n_516),
.B(n_505),
.Y(n_779)
);

AO21x1_ASAP7_75t_L g780 ( 
.A1(n_677),
.A2(n_506),
.B(n_467),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_664),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_743),
.A2(n_516),
.B(n_537),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_617),
.B(n_486),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_674),
.Y(n_784)
);

INVx3_ASAP7_75t_L g785 ( 
.A(n_712),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_746),
.A2(n_516),
.B(n_501),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_676),
.B(n_499),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_628),
.A2(n_501),
.B(n_499),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_682),
.B(n_474),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_747),
.A2(n_516),
.B(n_519),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_676),
.B(n_519),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_671),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_678),
.B(n_525),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_586),
.A2(n_528),
.B1(n_551),
.B2(n_548),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_663),
.A2(n_527),
.B(n_525),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_633),
.A2(n_529),
.B1(n_547),
.B2(n_535),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_663),
.A2(n_529),
.B(n_527),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_678),
.B(n_595),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_597),
.B(n_535),
.Y(n_799)
);

O2A1O1Ixp5_ASAP7_75t_L g800 ( 
.A1(n_694),
.A2(n_684),
.B(n_594),
.C(n_611),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_698),
.A2(n_547),
.B(n_521),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_705),
.A2(n_563),
.B(n_521),
.Y(n_802)
);

BUFx2_ASAP7_75t_SL g803 ( 
.A(n_664),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_620),
.B(n_563),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_626),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_590),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_598),
.B(n_452),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_728),
.A2(n_441),
.B(n_440),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_685),
.A2(n_563),
.B(n_521),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_712),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_681),
.A2(n_296),
.B(n_293),
.C(n_291),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_598),
.B(n_452),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_591),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_621),
.B(n_452),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_589),
.B(n_520),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_671),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_711),
.A2(n_563),
.B(n_531),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_621),
.B(n_521),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_718),
.B(n_563),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_592),
.A2(n_729),
.B1(n_630),
.B2(n_624),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_592),
.B(n_521),
.Y(n_821)
);

AND2x2_ASAP7_75t_SL g822 ( 
.A(n_714),
.B(n_264),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_708),
.B(n_531),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_607),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_734),
.A2(n_531),
.B(n_441),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_649),
.Y(n_826)
);

AND2x2_ASAP7_75t_SL g827 ( 
.A(n_717),
.B(n_270),
.Y(n_827)
);

OAI21xp33_ASAP7_75t_L g828 ( 
.A1(n_715),
.A2(n_238),
.B(n_237),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_650),
.A2(n_442),
.B(n_440),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_609),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_734),
.A2(n_531),
.B(n_443),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_744),
.A2(n_531),
.B(n_443),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_635),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_632),
.B(n_442),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_708),
.B(n_683),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_708),
.B(n_620),
.Y(n_836)
);

A2O1A1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_591),
.A2(n_414),
.B(n_291),
.C(n_296),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_622),
.A2(n_528),
.B1(n_509),
.B2(n_496),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_753),
.A2(n_449),
.B(n_445),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_755),
.A2(n_449),
.B(n_445),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_627),
.B(n_458),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_638),
.A2(n_640),
.B(n_713),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_707),
.A2(n_466),
.B(n_458),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_690),
.B(n_279),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_627),
.A2(n_528),
.B1(n_466),
.B2(n_509),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_596),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_596),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_632),
.B(n_459),
.Y(n_848)
);

AND2x2_ASAP7_75t_SL g849 ( 
.A(n_629),
.B(n_270),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_603),
.A2(n_619),
.B(n_604),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_707),
.A2(n_482),
.B(n_496),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_654),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_602),
.A2(n_482),
.B(n_491),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_603),
.A2(n_619),
.B(n_604),
.Y(n_854)
);

O2A1O1Ixp5_ASAP7_75t_L g855 ( 
.A1(n_639),
.A2(n_459),
.B(n_491),
.C(n_488),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_606),
.B(n_460),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_636),
.A2(n_462),
.B(n_488),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_636),
.A2(n_484),
.B(n_481),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_606),
.B(n_613),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_659),
.Y(n_860)
);

OAI21xp33_ASAP7_75t_L g861 ( 
.A1(n_686),
.A2(n_295),
.B(n_242),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_703),
.B(n_279),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_642),
.A2(n_460),
.B1(n_484),
.B2(n_481),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_SL g864 ( 
.A1(n_642),
.A2(n_462),
.B(n_297),
.C(n_274),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_606),
.B(n_398),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_613),
.B(n_511),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_613),
.B(n_398),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_703),
.B(n_279),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_653),
.A2(n_511),
.B(n_464),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_653),
.A2(n_511),
.B(n_464),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_658),
.A2(n_290),
.B(n_293),
.C(n_289),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_740),
.A2(n_741),
.B(n_716),
.C(n_691),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_689),
.B(n_511),
.Y(n_873)
);

NOR2xp67_ASAP7_75t_L g874 ( 
.A(n_675),
.B(n_274),
.Y(n_874)
);

AOI21x1_ASAP7_75t_L g875 ( 
.A1(n_689),
.A2(n_409),
.B(n_408),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_691),
.B(n_511),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_675),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_716),
.A2(n_511),
.B(n_464),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_724),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_655),
.A2(n_464),
.B(n_283),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_662),
.A2(n_289),
.B(n_290),
.C(n_285),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_667),
.A2(n_283),
.B(n_297),
.C(n_280),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_668),
.A2(n_464),
.B(n_404),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_610),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_721),
.A2(n_464),
.B(n_404),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_599),
.A2(n_383),
.B(n_404),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_600),
.A2(n_383),
.B(n_404),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_706),
.B(n_375),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_701),
.A2(n_285),
.B(n_280),
.C(n_263),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_735),
.B(n_398),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_699),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_720),
.A2(n_263),
.B1(n_398),
.B2(n_236),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_634),
.B(n_383),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_601),
.A2(n_383),
.B(n_404),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_605),
.A2(n_644),
.B(n_635),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_748),
.A2(n_252),
.B(n_408),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_720),
.A2(n_229),
.B1(n_154),
.B2(n_158),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_735),
.B(n_383),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_635),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_724),
.Y(n_900)
);

NOR2xp67_ASAP7_75t_L g901 ( 
.A(n_701),
.B(n_409),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_730),
.A2(n_235),
.B1(n_160),
.B2(n_164),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_670),
.B(n_383),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_712),
.B(n_383),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_635),
.A2(n_404),
.B(n_153),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_739),
.B(n_404),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_625),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_725),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_739),
.B(n_404),
.Y(n_909)
);

OAI21xp33_ASAP7_75t_L g910 ( 
.A1(n_661),
.A2(n_179),
.B(n_167),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_661),
.A2(n_409),
.B(n_179),
.C(n_408),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_635),
.B(n_404),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_641),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_643),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_644),
.A2(n_756),
.B(n_731),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_644),
.B(n_404),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_644),
.B(n_410),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_625),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_645),
.B(n_408),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_648),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_750),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_754),
.B(n_168),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_608),
.B(n_279),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_612),
.A2(n_616),
.B(n_615),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_631),
.B(n_673),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_644),
.A2(n_239),
.B(n_300),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_756),
.A2(n_217),
.B(n_298),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_647),
.A2(n_652),
.B(n_651),
.C(n_726),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_687),
.B(n_171),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_725),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_731),
.A2(n_246),
.B(n_294),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_756),
.A2(n_752),
.B(n_751),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_732),
.B(n_174),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_722),
.A2(n_6),
.B(n_8),
.C(n_10),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_756),
.A2(n_247),
.B1(n_292),
.B2(n_273),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_805),
.B(n_733),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_778),
.A2(n_756),
.B(n_748),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_815),
.A2(n_719),
.B(n_702),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_852),
.B(n_736),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_822),
.B(n_618),
.Y(n_940)
);

INVx4_ASAP7_75t_SL g941 ( 
.A(n_899),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_784),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_776),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_860),
.B(n_736),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_765),
.B(n_738),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_822),
.B(n_618),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_781),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_800),
.A2(n_889),
.B(n_872),
.C(n_928),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_770),
.A2(n_752),
.B(n_751),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_816),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_798),
.A2(n_889),
.B(n_871),
.C(n_811),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_899),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_862),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_757),
.A2(n_727),
.B(n_749),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_816),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_772),
.B(n_738),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_810),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_827),
.B(n_646),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_850),
.A2(n_646),
.B(n_749),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_781),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_L g961 ( 
.A(n_844),
.B(n_745),
.C(n_723),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_767),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_827),
.A2(n_745),
.B1(n_723),
.B2(n_710),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_820),
.B(n_648),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_770),
.A2(n_710),
.B(n_709),
.Y(n_965)
);

NAND2x1p5_ASAP7_75t_L g966 ( 
.A(n_810),
.B(n_709),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_914),
.B(n_913),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_834),
.A2(n_848),
.B1(n_821),
.B2(n_818),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_868),
.A2(n_775),
.B1(n_792),
.B2(n_759),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_865),
.A2(n_692),
.B1(n_679),
.B2(n_672),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_806),
.Y(n_971)
);

BUFx10_ASAP7_75t_L g972 ( 
.A(n_826),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_809),
.A2(n_692),
.B(n_679),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_834),
.A2(n_672),
.B1(n_669),
.B2(n_660),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_848),
.B(n_669),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_877),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_859),
.B(n_656),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_854),
.A2(n_660),
.B(n_657),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_764),
.B(n_657),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_764),
.B(n_656),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_803),
.Y(n_981)
);

BUFx8_ASAP7_75t_SL g982 ( 
.A(n_833),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_813),
.B(n_12),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_874),
.B(n_410),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_865),
.A2(n_212),
.B1(n_272),
.B2(n_271),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_846),
.B(n_13),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_L g987 ( 
.A(n_828),
.B(n_410),
.C(n_268),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_810),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_763),
.B(n_410),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_774),
.B(n_410),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_763),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_869),
.A2(n_410),
.B(n_259),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_847),
.B(n_14),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_802),
.A2(n_808),
.B(n_858),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_760),
.A2(n_410),
.B(n_257),
.C(n_251),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_921),
.B(n_177),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_879),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_900),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_891),
.Y(n_999)
);

OA22x2_ASAP7_75t_L g1000 ( 
.A1(n_861),
.A2(n_186),
.B1(n_189),
.B2(n_194),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_833),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_766),
.B(n_771),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_897),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_910),
.A2(n_410),
.B(n_250),
.C(n_248),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_817),
.A2(n_410),
.B(n_201),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_777),
.A2(n_410),
.B(n_196),
.C(n_195),
.Y(n_1006)
);

INVx6_ASAP7_75t_L g1007 ( 
.A(n_919),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_823),
.A2(n_15),
.B(n_17),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_898),
.B(n_21),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_766),
.B(n_22),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_890),
.B(n_24),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_812),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_789),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_762),
.A2(n_25),
.B(n_26),
.C(n_29),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_824),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_801),
.A2(n_26),
.B(n_32),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_L g1017 ( 
.A(n_934),
.B(n_33),
.C(n_34),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_SL g1018 ( 
.A(n_849),
.B(n_901),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_819),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_SL g1020 ( 
.A1(n_933),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_867),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_779),
.A2(n_43),
.B(n_44),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_849),
.B(n_50),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_842),
.A2(n_50),
.B(n_53),
.C(n_54),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_824),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_833),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_902),
.B(n_55),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_908),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_SL g1029 ( 
.A1(n_893),
.A2(n_788),
.B(n_814),
.C(n_807),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_925),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_1030)
);

NAND2xp33_ASAP7_75t_SL g1031 ( 
.A(n_771),
.B(n_56),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_807),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_814),
.A2(n_59),
.B(n_60),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_871),
.B(n_151),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_782),
.A2(n_61),
.B(n_70),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_867),
.A2(n_74),
.B1(n_80),
.B2(n_97),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_923),
.B(n_112),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_785),
.B(n_114),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_773),
.B(n_117),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_783),
.B(n_121),
.Y(n_1040)
);

A2O1A1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_893),
.A2(n_129),
.B(n_131),
.C(n_134),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_761),
.A2(n_139),
.B1(n_142),
.B2(n_143),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_830),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_929),
.B(n_148),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_866),
.B(n_856),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_832),
.A2(n_790),
.B(n_786),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_785),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_768),
.B(n_758),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_880),
.A2(n_882),
.B(n_924),
.C(n_829),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_769),
.A2(n_780),
.B(n_855),
.C(n_804),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_796),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_835),
.B(n_931),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_787),
.B(n_791),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_839),
.A2(n_840),
.B(n_885),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_935),
.B(n_930),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_793),
.B(n_918),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_896),
.A2(n_932),
.B(n_915),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_888),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_881),
.A2(n_911),
.B(n_795),
.C(n_797),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_884),
.B(n_907),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_912),
.A2(n_916),
.B(n_851),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_922),
.B(n_804),
.C(n_904),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_841),
.A2(n_836),
.B1(n_863),
.B2(n_903),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_949),
.A2(n_896),
.B(n_875),
.Y(n_1064)
);

AOI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_951),
.A2(n_911),
.B(n_799),
.Y(n_1065)
);

NOR2xp67_ASAP7_75t_L g1066 ( 
.A(n_1047),
.B(n_906),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1027),
.A2(n_892),
.B(n_895),
.C(n_909),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_939),
.B(n_920),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_SL g1069 ( 
.A(n_1045),
.B(n_904),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_994),
.A2(n_825),
.B(n_831),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_994),
.A2(n_912),
.B(n_916),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_952),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_962),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1014),
.A2(n_864),
.B(n_837),
.C(n_794),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_965),
.A2(n_857),
.B(n_843),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_942),
.Y(n_1076)
);

AO31x2_ASAP7_75t_L g1077 ( 
.A1(n_965),
.A2(n_918),
.A3(n_873),
.B(n_876),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_937),
.A2(n_917),
.B(n_845),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1003),
.B(n_927),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_944),
.B(n_926),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_1023),
.A2(n_838),
.B(n_883),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_937),
.A2(n_917),
.B(n_886),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_936),
.B(n_864),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_968),
.A2(n_887),
.B(n_894),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_971),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_953),
.B(n_905),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_L g1087 ( 
.A(n_1020),
.B(n_853),
.C(n_870),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_SL g1088 ( 
.A1(n_1018),
.A2(n_878),
.B1(n_1000),
.B2(n_1051),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_969),
.A2(n_1000),
.B1(n_950),
.B2(n_1034),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1054),
.A2(n_975),
.B(n_1049),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_952),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1054),
.A2(n_1046),
.B(n_948),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_1050),
.A2(n_1059),
.B(n_1063),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1044),
.A2(n_951),
.B(n_1033),
.C(n_1009),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1050),
.A2(n_938),
.B(n_1061),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_973),
.A2(n_1057),
.B(n_1046),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_1024),
.B(n_1030),
.C(n_1022),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_SL g1098 ( 
.A(n_947),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_955),
.B(n_943),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_952),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1053),
.A2(n_1029),
.B(n_1040),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1039),
.A2(n_1052),
.B(n_945),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_973),
.A2(n_959),
.B(n_1061),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_964),
.A2(n_978),
.B(n_992),
.Y(n_1104)
);

OR2x6_ASAP7_75t_L g1105 ( 
.A(n_960),
.B(n_999),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_978),
.A2(n_992),
.B(n_980),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1013),
.B(n_1032),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_997),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_998),
.Y(n_1109)
);

CKINVDCx11_ASAP7_75t_R g1110 ( 
.A(n_972),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_1037),
.A2(n_1011),
.B(n_1055),
.C(n_961),
.Y(n_1111)
);

BUFx5_ASAP7_75t_L g1112 ( 
.A(n_1038),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1021),
.B(n_1010),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_979),
.A2(n_974),
.B(n_1005),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1005),
.A2(n_1002),
.B(n_1035),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1035),
.A2(n_954),
.B(n_1031),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1028),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_967),
.B(n_996),
.Y(n_1118)
);

AO32x2_ASAP7_75t_L g1119 ( 
.A1(n_1019),
.A2(n_1042),
.A3(n_1012),
.B1(n_1036),
.B2(n_991),
.Y(n_1119)
);

AO31x2_ASAP7_75t_L g1120 ( 
.A1(n_995),
.A2(n_1004),
.A3(n_1048),
.B(n_1058),
.Y(n_1120)
);

AO21x2_ASAP7_75t_L g1121 ( 
.A1(n_938),
.A2(n_1006),
.B(n_1062),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_976),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1022),
.A2(n_1016),
.B(n_966),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_991),
.A2(n_1056),
.B(n_1038),
.Y(n_1124)
);

AO22x2_ASAP7_75t_L g1125 ( 
.A1(n_940),
.A2(n_958),
.B1(n_946),
.B2(n_1025),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_957),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_956),
.B(n_1045),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_981),
.B(n_1010),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_972),
.Y(n_1129)
);

AND2x6_ASAP7_75t_L g1130 ( 
.A(n_957),
.B(n_988),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_988),
.A2(n_977),
.B(n_970),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_983),
.B(n_993),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_986),
.A2(n_1008),
.B(n_1017),
.C(n_1041),
.Y(n_1133)
);

OAI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1045),
.A2(n_960),
.B1(n_985),
.B2(n_1007),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_989),
.A2(n_1047),
.B(n_987),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_989),
.A2(n_1047),
.B(n_1026),
.Y(n_1136)
);

BUFx8_ASAP7_75t_L g1137 ( 
.A(n_1001),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_963),
.A2(n_990),
.B(n_1060),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1007),
.B(n_941),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1007),
.B(n_1015),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1001),
.A2(n_984),
.B(n_1043),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_941),
.A2(n_965),
.B(n_949),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_984),
.A2(n_587),
.B(n_778),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_941),
.A2(n_587),
.B(n_1027),
.C(n_1023),
.Y(n_1144)
);

BUFx2_ASAP7_75t_SL g1145 ( 
.A(n_947),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_942),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_941),
.B(n_859),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_950),
.B(n_665),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_949),
.A2(n_965),
.B(n_973),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_942),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_953),
.B(n_665),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_939),
.B(n_805),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_972),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_968),
.A2(n_587),
.B1(n_765),
.B2(n_592),
.Y(n_1154)
);

NOR2x1_ASAP7_75t_R g1155 ( 
.A(n_960),
.B(n_495),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1023),
.A2(n_666),
.B1(n_1027),
.B2(n_587),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1018),
.B(n_822),
.Y(n_1158)
);

NOR2xp67_ASAP7_75t_L g1159 ( 
.A(n_1047),
.B(n_957),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_962),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_968),
.B(n_1053),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_949),
.A2(n_965),
.B(n_973),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1018),
.B(n_822),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_939),
.B(n_805),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_SL g1166 ( 
.A1(n_1029),
.A2(n_587),
.B(n_948),
.C(n_968),
.Y(n_1166)
);

OA21x2_ASAP7_75t_L g1167 ( 
.A1(n_1046),
.A2(n_1050),
.B(n_965),
.Y(n_1167)
);

NAND2x1p5_ASAP7_75t_L g1168 ( 
.A(n_952),
.B(n_810),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_SL g1169 ( 
.A(n_1003),
.B(n_495),
.C(n_614),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1027),
.A2(n_587),
.B(n_1023),
.C(n_1044),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_949),
.A2(n_965),
.B(n_973),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_972),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1027),
.A2(n_587),
.B(n_1023),
.C(n_1044),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_952),
.Y(n_1174)
);

OA21x2_ASAP7_75t_L g1175 ( 
.A1(n_1046),
.A2(n_1050),
.B(n_965),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_962),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1046),
.A2(n_1050),
.B(n_965),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_982),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_952),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1183)
);

OAI21x1_ASAP7_75t_L g1184 ( 
.A1(n_949),
.A2(n_965),
.B(n_973),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_972),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_942),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_949),
.A2(n_965),
.A3(n_770),
.B(n_769),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_994),
.A2(n_587),
.B(n_778),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_968),
.B(n_1053),
.Y(n_1191)
);

NOR2xp67_ASAP7_75t_L g1192 ( 
.A(n_1047),
.B(n_957),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_972),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_962),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_948),
.A2(n_587),
.B(n_1049),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_949),
.A2(n_965),
.B(n_973),
.Y(n_1196)
);

INVx6_ASAP7_75t_L g1197 ( 
.A(n_1137),
.Y(n_1197)
);

INVx6_ASAP7_75t_L g1198 ( 
.A(n_1137),
.Y(n_1198)
);

INVx6_ASAP7_75t_L g1199 ( 
.A(n_1072),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1073),
.Y(n_1200)
);

CKINVDCx6p67_ASAP7_75t_R g1201 ( 
.A(n_1178),
.Y(n_1201)
);

OAI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1156),
.A2(n_1158),
.B1(n_1164),
.B2(n_1154),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1151),
.B(n_1152),
.Y(n_1203)
);

BUFx8_ASAP7_75t_L g1204 ( 
.A(n_1098),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1165),
.B(n_1146),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1158),
.A2(n_1164),
.B1(n_1156),
.B2(n_1089),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1088),
.A2(n_1154),
.B1(n_1097),
.B2(n_1079),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1097),
.A2(n_1086),
.B1(n_1132),
.B2(n_1169),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1161),
.A2(n_1191),
.B1(n_1195),
.B2(n_1093),
.Y(n_1209)
);

INVx8_ASAP7_75t_L g1210 ( 
.A(n_1105),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1085),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1161),
.A2(n_1191),
.B1(n_1195),
.B2(n_1093),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1083),
.A2(n_1125),
.B1(n_1065),
.B2(n_1117),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1118),
.A2(n_1081),
.B1(n_1146),
.B2(n_1148),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1125),
.A2(n_1065),
.B1(n_1109),
.B2(n_1108),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1150),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1185),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1170),
.A2(n_1173),
.B1(n_1144),
.B2(n_1113),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1112),
.A2(n_1138),
.B1(n_1116),
.B2(n_1094),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1160),
.A2(n_1194),
.B1(n_1176),
.B2(n_1134),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1111),
.A2(n_1076),
.B1(n_1186),
.B2(n_1107),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1081),
.A2(n_1127),
.B1(n_1080),
.B2(n_1105),
.Y(n_1222)
);

BUFx8_ASAP7_75t_SL g1223 ( 
.A(n_1098),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1112),
.A2(n_1138),
.B1(n_1069),
.B2(n_1127),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1092),
.A2(n_1187),
.B(n_1181),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1129),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1099),
.A2(n_1128),
.B1(n_1124),
.B2(n_1122),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1140),
.A2(n_1087),
.B1(n_1112),
.B2(n_1068),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1110),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1091),
.B(n_1139),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1091),
.B(n_1112),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1100),
.B(n_1174),
.Y(n_1232)
);

CKINVDCx6p67_ASAP7_75t_R g1233 ( 
.A(n_1178),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_1178),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1145),
.B(n_1100),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1153),
.Y(n_1236)
);

INVx6_ASAP7_75t_L g1237 ( 
.A(n_1100),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_1172),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1147),
.A2(n_1101),
.B1(n_1141),
.B2(n_1121),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1133),
.A2(n_1074),
.B(n_1090),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1157),
.A2(n_1188),
.B1(n_1190),
.B2(n_1180),
.Y(n_1241)
);

BUFx12f_ASAP7_75t_L g1242 ( 
.A(n_1182),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1182),
.B(n_1193),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_SL g1244 ( 
.A1(n_1121),
.A2(n_1095),
.B1(n_1102),
.B2(n_1114),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1067),
.A2(n_1163),
.B1(n_1179),
.B2(n_1183),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1143),
.A2(n_1095),
.B1(n_1104),
.B2(n_1066),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1066),
.A2(n_1106),
.B1(n_1078),
.B2(n_1177),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1126),
.A2(n_1192),
.B1(n_1159),
.B2(n_1136),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1126),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1131),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1166),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1130),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1135),
.A2(n_1130),
.B1(n_1115),
.B2(n_1192),
.Y(n_1253)
);

OAI21xp33_ASAP7_75t_L g1254 ( 
.A1(n_1084),
.A2(n_1070),
.B(n_1071),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1168),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1123),
.A2(n_1119),
.B1(n_1175),
.B2(n_1167),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1167),
.A2(n_1177),
.B1(n_1175),
.B2(n_1130),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1142),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1120),
.Y(n_1259)
);

BUFx12f_ASAP7_75t_L g1260 ( 
.A(n_1155),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1082),
.A2(n_1119),
.B1(n_1064),
.B2(n_1075),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1096),
.A2(n_1103),
.B(n_1162),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1119),
.A2(n_1149),
.B1(n_1171),
.B2(n_1184),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1196),
.A2(n_1120),
.B1(n_1077),
.B2(n_1189),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1189),
.A2(n_1156),
.B1(n_1164),
.B2(n_1158),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1152),
.B(n_1165),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1156),
.A2(n_1164),
.B1(n_1158),
.B2(n_1154),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1073),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1073),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1073),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1110),
.Y(n_1271)
);

INVx5_ASAP7_75t_L g1272 ( 
.A(n_1130),
.Y(n_1272)
);

INVx3_ASAP7_75t_SL g1273 ( 
.A(n_1105),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1156),
.A2(n_1158),
.B1(n_1164),
.B2(n_1170),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_1110),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1110),
.Y(n_1276)
);

CKINVDCx6p67_ASAP7_75t_R g1277 ( 
.A(n_1178),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1170),
.A2(n_1173),
.B1(n_1156),
.B2(n_1154),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1156),
.A2(n_666),
.B1(n_1164),
.B2(n_1158),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1152),
.B(n_1165),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1156),
.A2(n_1164),
.B1(n_1158),
.B2(n_1154),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1156),
.A2(n_1164),
.B1(n_1158),
.B2(n_1154),
.Y(n_1282)
);

BUFx3_ASAP7_75t_L g1283 ( 
.A(n_1185),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1073),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_1098),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1073),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1158),
.A2(n_1164),
.B1(n_1018),
.B2(n_827),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1158),
.A2(n_1164),
.B1(n_1018),
.B2(n_827),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1156),
.A2(n_1158),
.B1(n_1164),
.B2(n_1170),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1156),
.A2(n_1164),
.B1(n_1158),
.B2(n_1154),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1158),
.A2(n_1164),
.B1(n_822),
.B2(n_827),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1156),
.A2(n_666),
.B1(n_1164),
.B2(n_1158),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1156),
.A2(n_666),
.B1(n_1164),
.B2(n_1158),
.Y(n_1293)
);

BUFx12f_ASAP7_75t_L g1294 ( 
.A(n_1110),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1110),
.Y(n_1295)
);

CKINVDCx11_ASAP7_75t_R g1296 ( 
.A(n_1110),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1073),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1073),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1152),
.B(n_1165),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1073),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1156),
.A2(n_816),
.B1(n_671),
.B2(n_1020),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1073),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1158),
.A2(n_1164),
.B1(n_1018),
.B2(n_827),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1158),
.A2(n_1164),
.B1(n_1018),
.B2(n_827),
.Y(n_1304)
);

INVxp67_ASAP7_75t_SL g1305 ( 
.A(n_1092),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1156),
.A2(n_1173),
.B(n_1170),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1073),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1200),
.B(n_1211),
.Y(n_1308)
);

AO21x1_ASAP7_75t_L g1309 ( 
.A1(n_1202),
.A2(n_1281),
.B(n_1267),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1305),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1250),
.Y(n_1311)
);

INVx2_ASAP7_75t_SL g1312 ( 
.A(n_1210),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1268),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1301),
.A2(n_1287),
.B1(n_1304),
.B2(n_1303),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1307),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1269),
.Y(n_1316)
);

OR2x6_ASAP7_75t_L g1317 ( 
.A(n_1252),
.B(n_1259),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1245),
.A2(n_1278),
.A3(n_1225),
.B(n_1262),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1270),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1284),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1286),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_1272),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1247),
.A2(n_1261),
.B(n_1263),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1258),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1297),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1298),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1300),
.Y(n_1327)
);

BUFx12f_ASAP7_75t_L g1328 ( 
.A(n_1271),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1251),
.A2(n_1248),
.B(n_1227),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1302),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1272),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1209),
.B(n_1212),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1305),
.Y(n_1333)
);

INVx2_ASAP7_75t_SL g1334 ( 
.A(n_1210),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1247),
.A2(n_1246),
.B(n_1257),
.Y(n_1335)
);

AO21x2_ASAP7_75t_L g1336 ( 
.A1(n_1265),
.A2(n_1214),
.B(n_1241),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1265),
.A2(n_1214),
.B(n_1241),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1246),
.A2(n_1257),
.B(n_1264),
.Y(n_1338)
);

INVx1_ASAP7_75t_SL g1339 ( 
.A(n_1238),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1209),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1212),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1252),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1231),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1287),
.A2(n_1304),
.B1(n_1303),
.B2(n_1288),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1254),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1249),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1266),
.B(n_1280),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1240),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1299),
.B(n_1205),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1216),
.Y(n_1350)
);

INVx4_ASAP7_75t_SL g1351 ( 
.A(n_1273),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1222),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1222),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1244),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1273),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1221),
.A2(n_1255),
.B(n_1232),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1244),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1219),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1213),
.A2(n_1306),
.B(n_1215),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1219),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1203),
.B(n_1213),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1256),
.B(n_1207),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1256),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1215),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1242),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1208),
.B(n_1289),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1199),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1199),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1218),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1239),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1199),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1224),
.Y(n_1372)
);

INVx1_ASAP7_75t_SL g1373 ( 
.A(n_1230),
.Y(n_1373)
);

INVx1_ASAP7_75t_SL g1374 ( 
.A(n_1226),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1243),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1274),
.B(n_1282),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1253),
.A2(n_1228),
.B(n_1293),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1224),
.Y(n_1378)
);

OR2x6_ASAP7_75t_L g1379 ( 
.A(n_1197),
.B(n_1198),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1220),
.Y(n_1380)
);

AOI21xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1202),
.A2(n_1281),
.B(n_1290),
.Y(n_1381)
);

AOI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1235),
.A2(n_1267),
.B(n_1290),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1279),
.B(n_1293),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1282),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1279),
.B(n_1292),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1375),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1348),
.A2(n_1292),
.B(n_1288),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1350),
.B(n_1236),
.Y(n_1388)
);

BUFx4f_ASAP7_75t_SL g1389 ( 
.A(n_1328),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1350),
.B(n_1234),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1348),
.B(n_1206),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1349),
.B(n_1277),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1322),
.B(n_1197),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1332),
.B(n_1201),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1308),
.B(n_1233),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1333),
.Y(n_1396)
);

BUFx12f_ASAP7_75t_L g1397 ( 
.A(n_1328),
.Y(n_1397)
);

NOR2x1_ASAP7_75t_SL g1398 ( 
.A(n_1322),
.B(n_1294),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1313),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1381),
.A2(n_1291),
.B(n_1295),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1351),
.B(n_1217),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1351),
.B(n_1217),
.Y(n_1402)
);

CKINVDCx14_ASAP7_75t_R g1403 ( 
.A(n_1328),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1381),
.A2(n_1283),
.B(n_1204),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1355),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1314),
.A2(n_1237),
.B1(n_1260),
.B2(n_1275),
.Y(n_1406)
);

NAND4xp25_ASAP7_75t_L g1407 ( 
.A(n_1332),
.B(n_1276),
.C(n_1296),
.D(n_1229),
.Y(n_1407)
);

NAND2xp33_ASAP7_75t_L g1408 ( 
.A(n_1342),
.B(n_1223),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1343),
.B(n_1285),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1333),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1373),
.B(n_1285),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1345),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1376),
.A2(n_1360),
.B(n_1358),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1329),
.A2(n_1356),
.B(n_1345),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1309),
.A2(n_1344),
.B1(n_1359),
.B2(n_1385),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1351),
.B(n_1317),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1347),
.B(n_1343),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_SL g1418 ( 
.A(n_1379),
.B(n_1342),
.Y(n_1418)
);

AO21x1_ASAP7_75t_L g1419 ( 
.A1(n_1366),
.A2(n_1362),
.B(n_1358),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1367),
.B(n_1371),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1367),
.B(n_1371),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1335),
.A2(n_1323),
.B(n_1338),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1363),
.B(n_1354),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1370),
.A2(n_1354),
.B(n_1357),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1369),
.A2(n_1383),
.B1(n_1385),
.B2(n_1360),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1315),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1383),
.A2(n_1369),
.B1(n_1359),
.B2(n_1384),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1340),
.A2(n_1341),
.B(n_1362),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1357),
.A2(n_1363),
.B1(n_1340),
.B2(n_1341),
.C(n_1369),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1377),
.A2(n_1353),
.B(n_1352),
.C(n_1384),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1316),
.B(n_1319),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1377),
.A2(n_1352),
.B(n_1353),
.C(n_1378),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1323),
.A2(n_1338),
.B(n_1309),
.Y(n_1434)
);

BUFx12f_ASAP7_75t_L g1435 ( 
.A(n_1365),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1319),
.B(n_1320),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1320),
.B(n_1321),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1368),
.A2(n_1312),
.A3(n_1334),
.B1(n_1331),
.B2(n_1361),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1359),
.A2(n_1337),
.B1(n_1336),
.B2(n_1380),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_SL g1440 ( 
.A1(n_1374),
.A2(n_1310),
.B(n_1339),
.C(n_1334),
.Y(n_1440)
);

NAND4xp25_ASAP7_75t_L g1441 ( 
.A(n_1346),
.B(n_1327),
.C(n_1326),
.D(n_1325),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1396),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1430),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1422),
.B(n_1318),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1396),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1417),
.B(n_1412),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_L g1447 ( 
.A(n_1441),
.B(n_1336),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1412),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1410),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1387),
.A2(n_1359),
.B(n_1382),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1422),
.B(n_1318),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1410),
.B(n_1337),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1399),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1438),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1386),
.B(n_1337),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_L g1456 ( 
.A(n_1393),
.B(n_1337),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1422),
.B(n_1318),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1432),
.B(n_1318),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1438),
.B(n_1318),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1436),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1439),
.B(n_1437),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1431),
.B(n_1325),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1438),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1414),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1438),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1430),
.B(n_1318),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1420),
.B(n_1311),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1431),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1434),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1433),
.B(n_1330),
.Y(n_1471)
);

INVxp67_ASAP7_75t_SL g1472 ( 
.A(n_1434),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1433),
.B(n_1330),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1421),
.B(n_1311),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1423),
.B(n_1326),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1427),
.B(n_1346),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1434),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1446),
.B(n_1423),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1442),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1454),
.B(n_1390),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1442),
.Y(n_1481)
);

INVx5_ASAP7_75t_SL g1482 ( 
.A(n_1470),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1445),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1445),
.Y(n_1484)
);

AOI322xp5_ASAP7_75t_L g1485 ( 
.A1(n_1447),
.A2(n_1415),
.A3(n_1427),
.B1(n_1429),
.B2(n_1391),
.C1(n_1394),
.C2(n_1403),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_SL g1486 ( 
.A(n_1455),
.B(n_1419),
.C(n_1415),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1454),
.B(n_1460),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1446),
.B(n_1424),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1460),
.B(n_1388),
.Y(n_1489)
);

AOI33xp33_ASAP7_75t_L g1490 ( 
.A1(n_1460),
.A2(n_1458),
.A3(n_1444),
.B1(n_1451),
.B2(n_1469),
.B3(n_1466),
.Y(n_1490)
);

BUFx2_ASAP7_75t_L g1491 ( 
.A(n_1448),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1446),
.B(n_1468),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1447),
.B(n_1418),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1409),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1462),
.A2(n_1455),
.B1(n_1472),
.B2(n_1469),
.C(n_1476),
.Y(n_1495)
);

OAI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1462),
.A2(n_1450),
.B1(n_1476),
.B2(n_1400),
.C(n_1471),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1449),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1449),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1416),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1453),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1474),
.B(n_1464),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1456),
.B(n_1416),
.Y(n_1502)
);

AND2x4_ASAP7_75t_L g1503 ( 
.A(n_1443),
.B(n_1416),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1464),
.B(n_1395),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1466),
.B(n_1405),
.Y(n_1505)
);

AOI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1463),
.A2(n_1440),
.B(n_1408),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1448),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1475),
.B(n_1407),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1450),
.A2(n_1364),
.B1(n_1428),
.B2(n_1372),
.Y(n_1509)
);

AND2x4_ASAP7_75t_SL g1510 ( 
.A(n_1467),
.B(n_1393),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1470),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1475),
.B(n_1424),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1471),
.A2(n_1364),
.B1(n_1378),
.B2(n_1372),
.Y(n_1513)
);

OAI211xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1465),
.A2(n_1403),
.B(n_1392),
.C(n_1411),
.Y(n_1514)
);

OAI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1473),
.A2(n_1413),
.B1(n_1406),
.B2(n_1425),
.C(n_1394),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1453),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_L g1517 ( 
.A(n_1452),
.B(n_1393),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1493),
.B(n_1472),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1493),
.B(n_1467),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1478),
.B(n_1452),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1493),
.B(n_1467),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1487),
.B(n_1444),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1500),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1487),
.B(n_1444),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1507),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1490),
.B(n_1461),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1511),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1492),
.B(n_1451),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1500),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1511),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.B(n_1451),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1516),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1511),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1491),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1482),
.Y(n_1535)
);

NOR3xp33_ASAP7_75t_SL g1536 ( 
.A(n_1514),
.B(n_1404),
.C(n_1389),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1479),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1479),
.B(n_1461),
.Y(n_1538)
);

INVx3_ASAP7_75t_L g1539 ( 
.A(n_1482),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1481),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1481),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1501),
.B(n_1458),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1483),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1483),
.B(n_1459),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1484),
.B(n_1459),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1489),
.B(n_1458),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1489),
.B(n_1459),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1512),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1501),
.B(n_1465),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1484),
.B(n_1457),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1491),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1482),
.B(n_1443),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1497),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1535),
.Y(n_1554)
);

OAI31xp33_ASAP7_75t_L g1555 ( 
.A1(n_1526),
.A2(n_1496),
.A3(n_1515),
.B(n_1506),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1522),
.B(n_1480),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1527),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1526),
.A2(n_1486),
.B1(n_1515),
.B2(n_1495),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1535),
.B(n_1493),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1535),
.B(n_1480),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1523),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1535),
.B(n_1510),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1523),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1535),
.B(n_1503),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1523),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1529),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1535),
.B(n_1508),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1539),
.B(n_1510),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1539),
.B(n_1504),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1544),
.B(n_1478),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1529),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1532),
.Y(n_1575)
);

NAND2x2_ASAP7_75t_L g1576 ( 
.A(n_1536),
.B(n_1389),
.Y(n_1576)
);

AOI211xp5_ASAP7_75t_L g1577 ( 
.A1(n_1518),
.A2(n_1440),
.B(n_1473),
.C(n_1463),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1527),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1534),
.A2(n_1485),
.B(n_1509),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1544),
.B(n_1497),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1527),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1545),
.B(n_1498),
.Y(n_1582)
);

NAND2xp33_ASAP7_75t_SL g1583 ( 
.A(n_1536),
.B(n_1494),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1539),
.B(n_1522),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1545),
.B(n_1498),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1522),
.B(n_1505),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1527),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1532),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1534),
.A2(n_1477),
.B(n_1517),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1537),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1538),
.B(n_1457),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1520),
.B(n_1488),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1539),
.B(n_1510),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1524),
.B(n_1504),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1532),
.Y(n_1595)
);

NOR2x1p5_ASAP7_75t_SL g1596 ( 
.A(n_1557),
.B(n_1548),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1573),
.B(n_1520),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1562),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1590),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1590),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1567),
.B(n_1397),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1562),
.B(n_1549),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1561),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1562),
.B(n_1570),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1549),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1561),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1579),
.A2(n_1513),
.B1(n_1518),
.B2(n_1502),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1555),
.B(n_1534),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1567),
.B(n_1397),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1555),
.B(n_1551),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1570),
.B(n_1549),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1558),
.A2(n_1519),
.B1(n_1521),
.B2(n_1524),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1558),
.B(n_1551),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1563),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1579),
.A2(n_1518),
.B1(n_1499),
.B2(n_1502),
.Y(n_1615)
);

INVxp33_ASAP7_75t_L g1616 ( 
.A(n_1570),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1563),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_SL g1618 ( 
.A(n_1570),
.B(n_1435),
.Y(n_1618)
);

OAI33xp33_ASAP7_75t_L g1619 ( 
.A1(n_1565),
.A2(n_1553),
.A3(n_1537),
.B1(n_1540),
.B2(n_1541),
.B3(n_1543),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1593),
.B(n_1519),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1557),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1593),
.B(n_1572),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1593),
.B(n_1524),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1593),
.B(n_1542),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1551),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1565),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1572),
.B(n_1542),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1584),
.B(n_1519),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1583),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1577),
.B(n_1547),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1599),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1604),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1599),
.Y(n_1633)
);

XNOR2x2_ASAP7_75t_L g1634 ( 
.A(n_1608),
.B(n_1589),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1604),
.B(n_1560),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1607),
.A2(n_1518),
.B1(n_1584),
.B2(n_1560),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1610),
.B(n_1554),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1625),
.A2(n_1589),
.B(n_1485),
.Y(n_1640)
);

AOI322xp5_ASAP7_75t_L g1641 ( 
.A1(n_1613),
.A2(n_1615),
.A3(n_1630),
.B1(n_1629),
.B2(n_1542),
.C1(n_1556),
.C2(n_1546),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1598),
.B(n_1594),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1598),
.B(n_1594),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1596),
.A2(n_1518),
.B(n_1592),
.C(n_1488),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1622),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1596),
.A2(n_1518),
.B(n_1592),
.C(n_1542),
.Y(n_1646)
);

OAI211xp5_ASAP7_75t_SL g1647 ( 
.A1(n_1600),
.A2(n_1612),
.B(n_1554),
.C(n_1626),
.Y(n_1647)
);

AOI222xp33_ASAP7_75t_L g1648 ( 
.A1(n_1619),
.A2(n_1548),
.B1(n_1556),
.B2(n_1477),
.C1(n_1587),
.C2(n_1578),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1616),
.A2(n_1576),
.B1(n_1559),
.B2(n_1556),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1603),
.A2(n_1569),
.B(n_1566),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_SL g1651 ( 
.A(n_1609),
.B(n_1576),
.C(n_1569),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1622),
.B(n_1547),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1621),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1603),
.Y(n_1654)
);

NAND2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1602),
.B(n_1564),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1640),
.A2(n_1637),
.B1(n_1645),
.B2(n_1646),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1653),
.Y(n_1657)
);

OAI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1634),
.A2(n_1618),
.B1(n_1576),
.B2(n_1597),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1653),
.Y(n_1659)
);

AOI32xp33_ASAP7_75t_L g1660 ( 
.A1(n_1647),
.A2(n_1602),
.A3(n_1605),
.B1(n_1611),
.B2(n_1627),
.Y(n_1660)
);

AOI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1639),
.A2(n_1621),
.B1(n_1623),
.B2(n_1605),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1642),
.B(n_1597),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1632),
.B(n_1627),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1643),
.B(n_1611),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1641),
.A2(n_1554),
.B(n_1606),
.C(n_1626),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1631),
.Y(n_1666)
);

NAND2x1_ASAP7_75t_L g1667 ( 
.A(n_1651),
.B(n_1620),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1635),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1654),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1639),
.A2(n_1614),
.B(n_1606),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1633),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1638),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1652),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1636),
.B(n_1620),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1668),
.B(n_1651),
.Y(n_1675)
);

XNOR2x1_ASAP7_75t_L g1676 ( 
.A(n_1658),
.B(n_1649),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1656),
.A2(n_1648),
.B1(n_1650),
.B2(n_1628),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1673),
.B(n_1624),
.Y(n_1678)
);

AND3x4_ASAP7_75t_L g1679 ( 
.A(n_1667),
.B(n_1620),
.C(n_1628),
.Y(n_1679)
);

AND3x1_ASAP7_75t_L g1680 ( 
.A(n_1674),
.B(n_1554),
.C(n_1623),
.Y(n_1680)
);

AOI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1658),
.A2(n_1665),
.B(n_1670),
.C(n_1659),
.Y(n_1681)
);

OAI21xp33_ASAP7_75t_L g1682 ( 
.A1(n_1661),
.A2(n_1644),
.B(n_1617),
.Y(n_1682)
);

INVxp67_ASAP7_75t_L g1683 ( 
.A(n_1657),
.Y(n_1683)
);

OAI211xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1660),
.A2(n_1614),
.B(n_1617),
.C(n_1655),
.Y(n_1684)
);

AOI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1671),
.A2(n_1672),
.B(n_1669),
.Y(n_1685)
);

AO22x2_ASAP7_75t_SL g1686 ( 
.A1(n_1662),
.A2(n_1624),
.B1(n_1564),
.B2(n_1568),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1678),
.Y(n_1687)
);

AND2x4_ASAP7_75t_SL g1688 ( 
.A(n_1675),
.B(n_1666),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1686),
.B(n_1663),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1679),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1680),
.B(n_1664),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_L g1692 ( 
.A(n_1682),
.B(n_1666),
.Y(n_1692)
);

OAI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1677),
.A2(n_1578),
.B1(n_1581),
.B2(n_1587),
.C(n_1557),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1683),
.Y(n_1694)
);

NAND4xp25_ASAP7_75t_L g1695 ( 
.A(n_1681),
.B(n_1685),
.C(n_1684),
.D(n_1682),
.Y(n_1695)
);

NAND3xp33_ASAP7_75t_SL g1696 ( 
.A(n_1690),
.B(n_1676),
.C(n_1365),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1693),
.A2(n_1628),
.B1(n_1581),
.B2(n_1578),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1695),
.A2(n_1587),
.B1(n_1581),
.B2(n_1566),
.C(n_1574),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1695),
.A2(n_1595),
.B1(n_1574),
.B2(n_1575),
.C(n_1588),
.Y(n_1699)
);

NOR3x1_ASAP7_75t_L g1700 ( 
.A(n_1689),
.B(n_1687),
.C(n_1694),
.Y(n_1700)
);

AOI221xp5_ASAP7_75t_L g1701 ( 
.A1(n_1698),
.A2(n_1692),
.B1(n_1691),
.B2(n_1688),
.C(n_1575),
.Y(n_1701)
);

AOI221xp5_ASAP7_75t_L g1702 ( 
.A1(n_1696),
.A2(n_1595),
.B1(n_1588),
.B2(n_1548),
.C(n_1530),
.Y(n_1702)
);

A2O1A1Ixp33_ASAP7_75t_SL g1703 ( 
.A1(n_1700),
.A2(n_1568),
.B(n_1571),
.C(n_1540),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1699),
.A2(n_1548),
.B1(n_1533),
.B2(n_1530),
.C(n_1525),
.Y(n_1704)
);

AOI222xp33_ASAP7_75t_L g1705 ( 
.A1(n_1697),
.A2(n_1533),
.B1(n_1530),
.B2(n_1525),
.C1(n_1546),
.C2(n_1547),
.Y(n_1705)
);

OA211x2_ASAP7_75t_L g1706 ( 
.A1(n_1696),
.A2(n_1591),
.B(n_1538),
.C(n_1550),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1706),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1701),
.Y(n_1708)
);

NAND4xp75_ASAP7_75t_L g1709 ( 
.A(n_1702),
.B(n_1571),
.C(n_1517),
.D(n_1586),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1705),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1703),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1704),
.B1(n_1585),
.B2(n_1582),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1708),
.A2(n_1711),
.B(n_1707),
.C(n_1710),
.Y(n_1713)
);

AOI322xp5_ASAP7_75t_L g1714 ( 
.A1(n_1709),
.A2(n_1546),
.A3(n_1586),
.B1(n_1530),
.B2(n_1533),
.C1(n_1528),
.C2(n_1531),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1712),
.Y(n_1715)
);

AO22x2_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1713),
.B1(n_1714),
.B2(n_1580),
.Y(n_1716)
);

XNOR2x1_ASAP7_75t_L g1717 ( 
.A(n_1716),
.B(n_1379),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1717),
.A2(n_1435),
.B1(n_1573),
.B2(n_1582),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1718),
.A2(n_1591),
.B(n_1585),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1719),
.A2(n_1580),
.B(n_1398),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1553),
.B1(n_1537),
.B2(n_1540),
.Y(n_1721)
);

AO21x2_ASAP7_75t_L g1722 ( 
.A1(n_1721),
.A2(n_1553),
.B(n_1543),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_R g1723 ( 
.A1(n_1722),
.A2(n_1528),
.B1(n_1531),
.B2(n_1541),
.C(n_1552),
.Y(n_1723)
);

AOI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1723),
.A2(n_1408),
.B(n_1402),
.C(n_1401),
.Y(n_1724)
);


endmodule