module real_aes_4212_n_296 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_1109, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_296);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_1109;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_296;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_503;
wire n_357;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_1034;
wire n_923;
wire n_952;
wire n_429;
wire n_976;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_370;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1053;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_973;
wire n_1081;
wire n_1084;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_404;
wire n_756;
wire n_598;
wire n_1073;
wire n_728;
wire n_334;
wire n_735;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_1105;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1028;
wire n_1003;
wire n_1014;
wire n_366;
wire n_346;
wire n_1083;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_712;
wire n_312;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_307;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_396;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g839 ( .A1(n_0), .A2(n_57), .B1(n_832), .B2(n_836), .Y(n_839) );
AOI21xp33_ASAP7_75t_L g1071 ( .A1(n_1), .A2(n_640), .B(n_1072), .Y(n_1071) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_2), .Y(n_307) );
AND2x4_ASAP7_75t_L g826 ( .A(n_2), .B(n_827), .Y(n_826) );
AND2x4_ASAP7_75t_L g835 ( .A(n_2), .B(n_287), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_3), .A2(n_294), .B1(n_430), .B2(n_433), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g794 ( .A1(n_4), .A2(n_35), .B1(n_795), .B2(n_796), .Y(n_794) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_5), .A2(n_204), .B1(n_380), .B2(n_387), .Y(n_1090) );
AOI22x1_ASAP7_75t_L g401 ( .A1(n_6), .A2(n_154), .B1(n_402), .B2(n_407), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_7), .A2(n_560), .B(n_712), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_8), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_9), .A2(n_201), .B1(n_479), .B2(n_485), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_10), .A2(n_261), .B1(n_804), .B2(n_805), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_11), .A2(n_174), .B1(n_487), .B2(n_488), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_12), .A2(n_89), .B1(n_825), .B2(n_829), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_13), .A2(n_147), .B1(n_352), .B2(n_639), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_14), .A2(n_151), .B1(n_799), .B2(n_801), .Y(n_798) );
CKINVDCx5p33_ASAP7_75t_R g600 ( .A(n_15), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g319 ( .A1(n_16), .A2(n_320), .B(n_345), .C(n_379), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_17), .A2(n_65), .B1(n_479), .B2(n_482), .Y(n_1063) );
XNOR2x1_ASAP7_75t_L g566 ( .A(n_18), .B(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_19), .A2(n_31), .B1(n_347), .B2(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g862 ( .A(n_20), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_21), .A2(n_146), .B1(n_403), .B2(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_22), .A2(n_191), .B1(n_478), .B2(n_484), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_23), .A2(n_286), .B1(n_511), .B2(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_24), .A2(n_87), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_25), .A2(n_72), .B1(n_565), .B2(n_633), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_26), .A2(n_83), .B1(n_867), .B2(n_879), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_27), .A2(n_188), .B1(n_572), .B2(n_1101), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_28), .A2(n_78), .B1(n_412), .B2(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_29), .A2(n_102), .B1(n_467), .B2(n_471), .Y(n_569) );
INVx1_ASAP7_75t_SL g672 ( .A(n_30), .Y(n_672) );
INVx1_ASAP7_75t_SL g932 ( .A(n_32), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_33), .A2(n_71), .B1(n_487), .B2(n_488), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_34), .A2(n_125), .B1(n_403), .B2(n_454), .Y(n_1102) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_36), .B(n_227), .Y(n_305) );
INVx1_ASAP7_75t_L g342 ( .A(n_36), .Y(n_342) );
INVxp67_ASAP7_75t_L g371 ( .A(n_36), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_37), .A2(n_139), .B1(n_416), .B2(n_444), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_38), .A2(n_73), .B1(n_411), .B2(n_415), .C(n_418), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_39), .A2(n_229), .B1(n_467), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_40), .A2(n_164), .B1(n_419), .B2(n_512), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_41), .A2(n_59), .B1(n_407), .B2(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g658 ( .A(n_42), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_43), .A2(n_111), .B1(n_402), .B2(n_609), .Y(n_608) );
OA22x2_ASAP7_75t_L g747 ( .A1(n_44), .A2(n_748), .B1(n_759), .B2(n_760), .Y(n_747) );
INVx1_ASAP7_75t_L g760 ( .A(n_44), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_44), .A2(n_94), .B1(n_858), .B2(n_872), .Y(n_880) );
AOI21xp33_ASAP7_75t_SL g1097 ( .A1(n_45), .A2(n_592), .B(n_1098), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_46), .A2(n_62), .B1(n_487), .B2(n_488), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_47), .B(n_347), .Y(n_797) );
INVx1_ASAP7_75t_L g475 ( .A(n_48), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_49), .A2(n_560), .B(n_574), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_50), .A2(n_117), .B1(n_380), .B2(n_387), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_51), .B(n_327), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_52), .A2(n_119), .B1(n_411), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_53), .A2(n_259), .B1(n_498), .B2(n_633), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_54), .A2(n_242), .B1(n_467), .B2(n_1075), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_55), .A2(n_108), .B1(n_592), .B2(n_605), .Y(n_767) );
INVx1_ASAP7_75t_SL g661 ( .A(n_56), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_58), .A2(n_254), .B1(n_403), .B2(n_501), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_60), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_61), .A2(n_177), .B1(n_864), .B2(n_870), .Y(n_869) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_63), .A2(n_233), .B1(n_470), .B2(n_471), .Y(n_469) );
INVxp67_ASAP7_75t_R g865 ( .A(n_64), .Y(n_865) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_66), .A2(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_SL g669 ( .A(n_67), .Y(n_669) );
INVx2_ASAP7_75t_L g302 ( .A(n_68), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_69), .A2(n_186), .B1(n_467), .B2(n_468), .Y(n_466) );
INVx1_ASAP7_75t_SL g828 ( .A(n_70), .Y(n_828) );
AND2x4_ASAP7_75t_L g830 ( .A(n_70), .B(n_302), .Y(n_830) );
INVx1_ASAP7_75t_L g834 ( .A(n_70), .Y(n_834) );
INVx1_ASAP7_75t_L g1099 ( .A(n_74), .Y(n_1099) );
INVx1_ASAP7_75t_SL g666 ( .A(n_75), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_76), .A2(n_84), .B1(n_683), .B2(n_685), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_77), .A2(n_187), .B1(n_505), .B2(n_507), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_79), .A2(n_203), .B1(n_362), .B2(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_80), .A2(n_268), .B1(n_432), .B2(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g791 ( .A(n_81), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_81), .A2(n_217), .B1(n_825), .B2(n_829), .Y(n_824) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_82), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_85), .A2(n_93), .B1(n_403), .B2(n_501), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_86), .A2(n_232), .B1(n_487), .B2(n_488), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_88), .A2(n_210), .B1(n_565), .B2(n_811), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_90), .A2(n_281), .B1(n_468), .B2(n_470), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_91), .A2(n_295), .B1(n_481), .B2(n_485), .Y(n_579) );
INVx1_ASAP7_75t_L g766 ( .A(n_92), .Y(n_766) );
CKINVDCx16_ASAP7_75t_R g860 ( .A(n_95), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_96), .A2(n_182), .B1(n_858), .B2(n_918), .Y(n_917) );
AO22x1_ASAP7_75t_L g379 ( .A1(n_97), .A2(n_274), .B1(n_380), .B2(n_387), .Y(n_379) );
INVx1_ASAP7_75t_L g575 ( .A(n_98), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_99), .A2(n_183), .B1(n_631), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_100), .A2(n_257), .B1(n_478), .B2(n_484), .Y(n_752) );
INVx1_ASAP7_75t_L g328 ( .A(n_101), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_101), .B(n_226), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_103), .A2(n_194), .B1(n_529), .B2(n_531), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_104), .A2(n_285), .B1(n_444), .B2(n_525), .Y(n_598) );
INVx1_ASAP7_75t_L g597 ( .A(n_105), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_106), .A2(n_272), .B1(n_479), .B2(n_482), .Y(n_577) );
XNOR2x1_ASAP7_75t_L g705 ( .A(n_107), .B(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g555 ( .A1(n_109), .A2(n_166), .B1(n_556), .B2(n_558), .C(n_561), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_110), .A2(n_158), .B1(n_468), .B2(n_470), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_112), .A2(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_SL g689 ( .A(n_113), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_114), .A2(n_219), .B1(n_380), .B2(n_503), .Y(n_629) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_115), .A2(n_256), .B1(n_407), .B2(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_116), .A2(n_288), .B1(n_481), .B2(n_482), .Y(n_750) );
AOI221xp5_ASAP7_75t_SL g754 ( .A1(n_118), .A2(n_263), .B1(n_470), .B2(n_640), .C(n_755), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_120), .A2(n_167), .B1(n_456), .B2(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g846 ( .A(n_121), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_122), .A2(n_185), .B1(n_870), .B2(n_879), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_123), .A2(n_255), .B1(n_407), .B2(n_511), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_124), .B(n_1069), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_126), .A2(n_235), .B1(n_362), .B2(n_372), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g756 ( .A(n_127), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_128), .A2(n_196), .B1(n_467), .B2(n_471), .C(n_758), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_129), .A2(n_260), .B1(n_482), .B2(n_484), .Y(n_717) );
CKINVDCx14_ASAP7_75t_R g317 ( .A(n_130), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_131), .A2(n_163), .B1(n_444), .B2(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_132), .B(n_446), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_133), .B(n_640), .Y(n_710) );
INVx1_ASAP7_75t_L g603 ( .A(n_134), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_135), .A2(n_197), .B1(n_446), .B2(n_448), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_136), .A2(n_155), .B1(n_432), .B2(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g722 ( .A(n_137), .Y(n_722) );
NAND2xp33_ASAP7_75t_L g429 ( .A(n_138), .B(n_430), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_140), .A2(n_206), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g713 ( .A(n_141), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_142), .A2(n_175), .B1(n_479), .B2(n_485), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_143), .A2(n_179), .B1(n_511), .B2(n_631), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_144), .A2(n_190), .B1(n_864), .B2(n_867), .Y(n_933) );
INVx1_ASAP7_75t_L g651 ( .A(n_145), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_148), .A2(n_279), .B1(n_470), .B2(n_481), .Y(n_715) );
AO22x1_ASAP7_75t_L g418 ( .A1(n_149), .A2(n_211), .B1(n_419), .B2(n_421), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_150), .A2(n_152), .B1(n_481), .B2(n_485), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_153), .A2(n_237), .B1(n_467), .B2(n_468), .Y(n_709) );
INVx1_ASAP7_75t_L g1073 ( .A(n_156), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_157), .A2(n_225), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_159), .A2(n_161), .B1(n_503), .B2(n_631), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_160), .A2(n_208), .B1(n_478), .B2(n_484), .Y(n_578) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_162), .A2(n_202), .B1(n_533), .B2(n_535), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_165), .A2(n_270), .B1(n_403), .B2(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g660 ( .A(n_168), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_169), .A2(n_262), .B1(n_832), .B2(n_836), .Y(n_831) );
INVx1_ASAP7_75t_L g850 ( .A(n_170), .Y(n_850) );
AO22x1_ASAP7_75t_L g758 ( .A1(n_171), .A2(n_253), .B1(n_468), .B2(n_560), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_172), .A2(n_258), .B1(n_478), .B2(n_479), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_173), .A2(n_234), .B1(n_617), .B2(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g848 ( .A(n_176), .Y(n_848) );
INVx1_ASAP7_75t_L g1076 ( .A(n_177), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_177), .A2(n_1083), .B1(n_1103), .B2(n_1105), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_178), .A2(n_1084), .B1(n_1085), .B2(n_1086), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g1084 ( .A(n_178), .Y(n_1084) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_180), .A2(n_218), .B1(n_500), .B2(n_502), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_181), .A2(n_184), .B1(n_498), .B2(n_633), .Y(n_1089) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_182), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_189), .B(n_448), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_192), .A2(n_278), .B1(n_419), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_193), .A2(n_239), .B1(n_471), .B2(n_478), .Y(n_708) );
INVx1_ASAP7_75t_L g733 ( .A(n_195), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_198), .A2(n_267), .B1(n_395), .B2(n_614), .Y(n_613) );
OA22x2_ASAP7_75t_L g332 ( .A1(n_199), .A2(n_227), .B1(n_327), .B2(n_331), .Y(n_332) );
INVx1_ASAP7_75t_L g358 ( .A(n_199), .Y(n_358) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_200), .A2(n_222), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_205), .A2(n_243), .B1(n_347), .B2(n_731), .C(n_732), .Y(n_730) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_207), .A2(n_516), .B(n_520), .Y(n_515) );
AOI221x1_ASAP7_75t_L g764 ( .A1(n_209), .A2(n_250), .B1(n_518), .B2(n_668), .C(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_212), .A2(n_220), .B1(n_407), .B2(n_635), .Y(n_775) );
INVx1_ASAP7_75t_L g527 ( .A(n_213), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_214), .A2(n_230), .B1(n_391), .B2(n_395), .C(n_400), .Y(n_390) );
AOI221x1_ASAP7_75t_L g431 ( .A1(n_215), .A2(n_266), .B1(n_432), .B2(n_433), .C(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g523 ( .A(n_216), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_221), .A2(n_265), .B1(n_391), .B2(n_633), .Y(n_632) );
CKINVDCx6p67_ASAP7_75t_R g859 ( .A(n_223), .Y(n_859) );
AO22x2_ASAP7_75t_L g493 ( .A1(n_224), .A2(n_494), .B1(n_538), .B2(n_539), .Y(n_493) );
INVx1_ASAP7_75t_L g539 ( .A(n_224), .Y(n_539) );
INVx1_ASAP7_75t_L g344 ( .A(n_226), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_226), .B(n_356), .Y(n_378) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_227), .A2(n_240), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g434 ( .A(n_228), .B(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g871 ( .A1(n_231), .A2(n_245), .B1(n_858), .B2(n_872), .Y(n_871) );
INVx1_ASAP7_75t_SL g695 ( .A(n_236), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_238), .A2(n_252), .B1(n_736), .B2(n_737), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_240), .B(n_282), .Y(n_306) );
INVx1_ASAP7_75t_L g330 ( .A(n_240), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g692 ( .A(n_241), .Y(n_692) );
INVx1_ASAP7_75t_L g562 ( .A(n_244), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_246), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g462 ( .A(n_247), .Y(n_462) );
OAI21x1_ASAP7_75t_L g761 ( .A1(n_248), .A2(n_762), .B(n_780), .Y(n_761) );
INVx1_ASAP7_75t_L g783 ( .A(n_248), .Y(n_783) );
XNOR2x1_ASAP7_75t_L g543 ( .A(n_249), .B(n_544), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_251), .A2(n_292), .B1(n_736), .B2(n_805), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_264), .A2(n_269), .B1(n_510), .B2(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_271), .B(n_731), .Y(n_1096) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_273), .B(n_428), .C(n_436), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_273), .A2(n_436), .B1(n_442), .B2(n_1109), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g459 ( .A1(n_273), .A2(n_428), .B(n_451), .Y(n_459) );
INVx1_ASAP7_75t_SL g688 ( .A(n_275), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_276), .A2(n_290), .B1(n_352), .B2(n_592), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_277), .A2(n_284), .B1(n_511), .B2(n_813), .Y(n_812) );
AOI22xp5_ASAP7_75t_SL g1070 ( .A1(n_280), .A2(n_291), .B1(n_468), .B2(n_470), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_282), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_283), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g827 ( .A(n_287), .Y(n_827) );
INVx1_ASAP7_75t_L g622 ( .A(n_289), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_293), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_308), .B(n_817), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx4_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .C(n_307), .Y(n_299) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_300), .B(n_1080), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1104 ( .A(n_300), .B(n_1081), .Y(n_1104) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OA21x2_ASAP7_75t_L g1106 ( .A1(n_301), .A2(n_828), .B(n_1107), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND3x4_ASAP7_75t_L g825 ( .A(n_302), .B(n_826), .C(n_828), .Y(n_825) );
AND2x2_ASAP7_75t_L g833 ( .A(n_302), .B(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g1080 ( .A(n_303), .B(n_1081), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_304), .A2(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g1081 ( .A(n_307), .Y(n_1081) );
OAI22xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B1(n_700), .B2(n_701), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
XNOR2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_490), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
XNOR2x1_ASAP7_75t_L g314 ( .A(n_315), .B(n_424), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
XNOR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NAND3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_390), .C(n_410), .Y(n_318) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx3_ASAP7_75t_SL g731 ( .A(n_322), .Y(n_731) );
INVx2_ASAP7_75t_L g795 ( .A(n_322), .Y(n_795) );
INVx2_ASAP7_75t_L g1069 ( .A(n_322), .Y(n_1069) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g447 ( .A(n_323), .Y(n_447) );
BUFx3_ASAP7_75t_L g647 ( .A(n_323), .Y(n_647) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_333), .Y(n_323) );
AND2x2_ASAP7_75t_L g414 ( .A(n_324), .B(n_399), .Y(n_414) );
AND2x2_ASAP7_75t_L g420 ( .A(n_324), .B(n_405), .Y(n_420) );
AND2x4_ASAP7_75t_L g422 ( .A(n_324), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g435 ( .A(n_324), .B(n_405), .Y(n_435) );
AND2x4_ASAP7_75t_L g467 ( .A(n_324), .B(n_399), .Y(n_467) );
AND2x4_ASAP7_75t_L g481 ( .A(n_324), .B(n_405), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_324), .B(n_384), .Y(n_482) );
AND2x2_ASAP7_75t_L g560 ( .A(n_324), .B(n_333), .Y(n_560) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_332), .Y(n_324) );
INVx1_ASAP7_75t_L g351 ( .A(n_325), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_329), .Y(n_325) );
NAND2xp33_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g331 ( .A(n_327), .Y(n_331) );
INVx3_ASAP7_75t_L g337 ( .A(n_327), .Y(n_337) );
NAND2xp33_ASAP7_75t_L g343 ( .A(n_327), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_328), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_330), .A2(n_360), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g350 ( .A(n_332), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g383 ( .A(n_332), .Y(n_383) );
AND2x4_ASAP7_75t_L g349 ( .A(n_333), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g353 ( .A(n_333), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g394 ( .A(n_333), .B(n_382), .Y(n_394) );
AND2x4_ASAP7_75t_L g468 ( .A(n_333), .B(n_354), .Y(n_468) );
AND2x2_ASAP7_75t_L g473 ( .A(n_333), .B(n_350), .Y(n_473) );
AND2x4_ASAP7_75t_L g488 ( .A(n_333), .B(n_382), .Y(n_488) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_339), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g365 ( .A(n_335), .B(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g385 ( .A(n_335), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g399 ( .A(n_335), .B(n_339), .Y(n_399) );
AND2x4_ASAP7_75t_L g405 ( .A(n_335), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_337), .B(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g356 ( .A(n_337), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_338), .B(n_355), .C(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g386 ( .A(n_340), .Y(n_386) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_361), .Y(n_345) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g440 ( .A(n_349), .Y(n_440) );
BUFx8_ASAP7_75t_SL g530 ( .A(n_349), .Y(n_530) );
INVx2_ASAP7_75t_L g557 ( .A(n_349), .Y(n_557) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_349), .Y(n_572) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_349), .Y(n_640) );
AND2x4_ASAP7_75t_L g417 ( .A(n_350), .B(n_399), .Y(n_417) );
AND2x4_ASAP7_75t_L g470 ( .A(n_350), .B(n_399), .Y(n_470) );
AND2x4_ASAP7_75t_L g382 ( .A(n_351), .B(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g531 ( .A(n_352), .Y(n_531) );
INVx4_ASAP7_75t_L g670 ( .A(n_352), .Y(n_670) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_353), .Y(n_438) );
INVx3_ASAP7_75t_L g802 ( .A(n_353), .Y(n_802) );
AND2x4_ASAP7_75t_L g389 ( .A(n_354), .B(n_384), .Y(n_389) );
AND2x4_ASAP7_75t_L g409 ( .A(n_354), .B(n_405), .Y(n_409) );
AND2x4_ASAP7_75t_L g479 ( .A(n_354), .B(n_384), .Y(n_479) );
AND2x4_ASAP7_75t_L g485 ( .A(n_354), .B(n_405), .Y(n_485) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_359), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx4_ASAP7_75t_L g444 ( .A(n_363), .Y(n_444) );
INVx2_ASAP7_75t_L g522 ( .A(n_363), .Y(n_522) );
INVx2_ASAP7_75t_L g551 ( .A(n_363), .Y(n_551) );
INVx2_ASAP7_75t_L g737 ( .A(n_363), .Y(n_737) );
INVx5_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g650 ( .A(n_364), .Y(n_650) );
BUFx2_ASAP7_75t_L g805 ( .A(n_364), .Y(n_805) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_369), .Y(n_364) );
AND2x2_ASAP7_75t_L g471 ( .A(n_365), .B(n_369), .Y(n_471) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_365), .B(n_369), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVx1_ASAP7_75t_L g376 ( .A(n_367), .Y(n_376) );
INVx2_ASAP7_75t_L g734 ( .A(n_372), .Y(n_734) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_373), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_373), .B(n_713), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_373), .B(n_766), .Y(n_765) );
INVx4_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g526 ( .A(n_374), .Y(n_526) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_375), .Y(n_450) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_381), .Y(n_501) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_381), .Y(n_618) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
AND2x4_ASAP7_75t_L g398 ( .A(n_382), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g404 ( .A(n_382), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g478 ( .A(n_382), .B(n_423), .Y(n_478) );
AND2x4_ASAP7_75t_L g484 ( .A(n_382), .B(n_405), .Y(n_484) );
AND2x4_ASAP7_75t_L g487 ( .A(n_382), .B(n_399), .Y(n_487) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g423 ( .A(n_385), .Y(n_423) );
INVx1_ASAP7_75t_L g406 ( .A(n_386), .Y(n_406) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx5_ASAP7_75t_L g430 ( .A(n_388), .Y(n_430) );
INVx2_ASAP7_75t_L g621 ( .A(n_388), .Y(n_621) );
INVx3_ASAP7_75t_L g808 ( .A(n_388), .Y(n_808) );
INVx6_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx12f_ASAP7_75t_L g503 ( .A(n_389), .Y(n_503) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g615 ( .A(n_392), .Y(n_615) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx3_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
BUFx5_ASAP7_75t_L g498 ( .A(n_394), .Y(n_498) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_394), .Y(n_565) );
BUFx4f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g811 ( .A(n_397), .Y(n_811) );
INVx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx12f_ASAP7_75t_L g432 ( .A(n_398), .Y(n_432) );
BUFx6f_ASAP7_75t_L g633 ( .A(n_398), .Y(n_633) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx12f_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g681 ( .A(n_403), .Y(n_681) );
BUFx12f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_404), .Y(n_506) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_404), .Y(n_635) );
INVx4_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g454 ( .A(n_408), .Y(n_454) );
INVx2_ASAP7_75t_L g508 ( .A(n_408), .Y(n_508) );
INVx2_ASAP7_75t_SL g549 ( .A(n_408), .Y(n_549) );
INVx4_ASAP7_75t_L g610 ( .A(n_408), .Y(n_610) );
INVx2_ASAP7_75t_L g813 ( .A(n_408), .Y(n_813) );
INVx8_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g770 ( .A(n_412), .Y(n_770) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_413), .Y(n_664) );
INVx1_ASAP7_75t_L g736 ( .A(n_413), .Y(n_736) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g537 ( .A(n_414), .Y(n_537) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_414), .Y(n_804) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g643 ( .A(n_416), .Y(n_643) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx3_ASAP7_75t_L g534 ( .A(n_417), .Y(n_534) );
BUFx6f_ASAP7_75t_L g592 ( .A(n_417), .Y(n_592) );
INVx1_ASAP7_75t_L g800 ( .A(n_417), .Y(n_800) );
BUFx8_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_420), .Y(n_511) );
INVx1_ASAP7_75t_L g690 ( .A(n_421), .Y(n_690) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_422), .Y(n_456) );
BUFx12f_ASAP7_75t_L g513 ( .A(n_422), .Y(n_513) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_422), .Y(n_631) );
BUFx6f_ASAP7_75t_L g1094 ( .A(n_422), .Y(n_1094) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_460), .B2(n_461), .Y(n_424) );
INVx2_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
AO21x2_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_441), .B(n_457), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_432), .Y(n_694) );
BUFx4f_ASAP7_75t_L g547 ( .A(n_435), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_437), .B(n_439), .Y(n_436) );
BUFx3_ASAP7_75t_L g605 ( .A(n_438), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_451), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_445), .Y(n_442) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_447), .Y(n_519) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_450), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_450), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_SL g676 ( .A(n_450), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_450), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g796 ( .A(n_450), .Y(n_796) );
NAND2x1_ASAP7_75t_SL g451 ( .A(n_452), .B(n_455), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AO21x2_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B(n_489), .Y(n_461) );
NOR3xp33_ASAP7_75t_SL g489 ( .A(n_462), .B(n_464), .C(n_476), .Y(n_489) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_476), .Y(n_463) );
NAND4xp75_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .C(n_469), .D(n_472), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .C(n_483), .D(n_486), .Y(n_476) );
XNOR2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_585), .Y(n_490) );
XOR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_540), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
NOR2x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_514), .Y(n_494) );
NAND4xp25_ASAP7_75t_L g495 ( .A(n_496), .B(n_499), .C(n_504), .D(n_509), .Y(n_495) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_SL g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g687 ( .A(n_510), .Y(n_687) );
BUFx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_528), .C(n_532), .Y(n_514) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
OAI21xp33_ASAP7_75t_L g596 ( .A1(n_517), .A2(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g674 ( .A(n_519), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_523), .B1(n_524), .B2(n_527), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g1072 ( .A(n_526), .B(n_1073), .Y(n_1072) );
NOR2xp33_ASAP7_75t_L g1098 ( .A(n_526), .B(n_1099), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g595 ( .A(n_537), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_566), .B1(n_581), .B2(n_583), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g582 ( .A(n_543), .Y(n_582) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_546), .B(n_548), .C(n_550), .D(n_552), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .C(n_564), .Y(n_553) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g668 ( .A(n_557), .Y(n_668) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g696 ( .A(n_565), .Y(n_696) );
INVx2_ASAP7_75t_L g584 ( .A(n_566), .Y(n_584) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_576), .Y(n_567) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .C(n_571), .D(n_573), .Y(n_568) );
BUFx3_ASAP7_75t_L g602 ( .A(n_572), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .C(n_579), .D(n_580), .Y(n_576) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
XNOR2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_623), .Y(n_585) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_622), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_606), .Y(n_587) );
NOR3xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_596), .C(n_599), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_593), .B2(n_594), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_591), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
INVx4_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_601), .B1(n_603), .B2(n_604), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp67_ASAP7_75t_L g606 ( .A(n_607), .B(n_612), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .Y(n_607) );
BUFx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g684 ( .A(n_618), .Y(n_684) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g685 ( .A(n_620), .Y(n_685) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_654), .B1(n_655), .B2(n_699), .Y(n_623) );
INVx2_ASAP7_75t_L g699 ( .A(n_624), .Y(n_699) );
AO21x2_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B(n_653), .Y(n_624) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_625), .B(n_628), .C(n_637), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_636), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND4xp25_ASAP7_75t_SL g628 ( .A(n_629), .B(n_630), .C(n_632), .D(n_634), .Y(n_628) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .C(n_644), .Y(n_637) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI21xp5_ASAP7_75t_SL g648 ( .A1(n_649), .A2(n_651), .B(n_652), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx4_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AO22x2_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_657), .B1(n_677), .B2(n_697), .Y(n_655) );
NOR4xp25_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .C(n_665), .D(n_671), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g657 ( .A(n_658), .Y(n_657) );
NOR3xp33_ASAP7_75t_SL g698 ( .A(n_659), .B(n_665), .C(n_671), .Y(n_698) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_669), .B2(n_670), .Y(n_665) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_677), .B(n_698), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_686), .C(n_691), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_686) );
OAI22x1_ASAP7_75t_SL g691 ( .A1(n_692), .A2(n_693), .B1(n_695), .B2(n_696), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
XNOR2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_741), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_719), .B1(n_739), .B2(n_740), .Y(n_702) );
INVx2_ASAP7_75t_L g739 ( .A(n_703), .Y(n_739) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_714), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .C(n_710), .D(n_711), .Y(n_707) );
NAND4xp25_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .C(n_717), .D(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g740 ( .A(n_719), .Y(n_740) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
XNOR2x1_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_729), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .C(n_727), .D(n_728), .Y(n_724) );
NAND3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_735), .C(n_738), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_742), .A2(n_743), .B1(n_814), .B2(n_815), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_787), .B2(n_788), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
XNOR2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_761), .Y(n_746) );
INVx2_ASAP7_75t_L g816 ( .A(n_747), .Y(n_816) );
INVx1_ASAP7_75t_L g759 ( .A(n_748), .Y(n_759) );
NAND3xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_754), .C(n_757), .Y(n_748) );
AND4x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .C(n_752), .D(n_753), .Y(n_749) );
NOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_771), .Y(n_762) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_767), .C(n_768), .Y(n_763) );
INVx1_ASAP7_75t_L g785 ( .A(n_764), .Y(n_785) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_767), .Y(n_786) );
INVx1_ASAP7_75t_L g782 ( .A(n_768), .Y(n_782) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_776), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_773), .B(n_782), .C(n_783), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_777), .B(n_785), .C(n_786), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_784), .Y(n_780) );
OAI221xp5_ASAP7_75t_L g931 ( .A1(n_783), .A2(n_847), .B1(n_857), .B2(n_932), .C(n_933), .Y(n_931) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
XNOR2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g790 ( .A(n_791), .Y(n_790) );
NOR2x1_ASAP7_75t_L g792 ( .A(n_793), .B(n_806), .Y(n_792) );
NAND4xp25_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .C(n_798), .D(n_803), .Y(n_793) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx3_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g1101 ( .A(n_802), .Y(n_1101) );
NAND4xp25_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .C(n_810), .D(n_812), .Y(n_806) );
INVx1_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
BUFx4_ASAP7_75t_R g815 ( .A(n_816), .Y(n_815) );
OAI221xp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_1056), .B1(n_1058), .B2(n_1077), .C(n_1082), .Y(n_817) );
NOR3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_979), .C(n_1022), .Y(n_818) );
NAND5xp2_ASAP7_75t_L g819 ( .A(n_820), .B(n_920), .C(n_949), .D(n_958), .E(n_974), .Y(n_819) );
OAI31xp33_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_873), .A3(n_894), .B(n_910), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_840), .Y(n_821) );
INVx1_ASAP7_75t_L g997 ( .A(n_822), .Y(n_997) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_837), .Y(n_822) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_823), .Y(n_881) );
AND2x2_ASAP7_75t_L g905 ( .A(n_823), .B(n_877), .Y(n_905) );
AND2x2_ASAP7_75t_L g925 ( .A(n_823), .B(n_884), .Y(n_925) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_823), .B(n_837), .Y(n_1021) );
AND2x4_ASAP7_75t_SL g823 ( .A(n_824), .B(n_831), .Y(n_823) );
INVx1_ASAP7_75t_L g845 ( .A(n_825), .Y(n_845) );
AND2x4_ASAP7_75t_L g829 ( .A(n_826), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_826), .B(n_830), .Y(n_847) );
AND2x4_ASAP7_75t_L g858 ( .A(n_826), .B(n_833), .Y(n_858) );
AND2x4_ASAP7_75t_L g872 ( .A(n_826), .B(n_830), .Y(n_872) );
INVx2_ASAP7_75t_SL g919 ( .A(n_829), .Y(n_919) );
AND2x2_ASAP7_75t_L g836 ( .A(n_830), .B(n_835), .Y(n_836) );
AND2x4_ASAP7_75t_L g867 ( .A(n_830), .B(n_835), .Y(n_867) );
AND2x2_ASAP7_75t_L g870 ( .A(n_830), .B(n_835), .Y(n_870) );
INVx1_ASAP7_75t_L g853 ( .A(n_832), .Y(n_853) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
AND2x4_ASAP7_75t_L g864 ( .A(n_833), .B(n_835), .Y(n_864) );
AND2x2_ASAP7_75t_L g879 ( .A(n_833), .B(n_835), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g1107 ( .A(n_835), .Y(n_1107) );
INVx1_ASAP7_75t_L g851 ( .A(n_836), .Y(n_851) );
AND2x2_ASAP7_75t_L g875 ( .A(n_837), .B(n_876), .Y(n_875) );
CKINVDCx6p67_ASAP7_75t_R g886 ( .A(n_837), .Y(n_886) );
INVx1_ASAP7_75t_L g900 ( .A(n_837), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_837), .B(n_881), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_837), .B(n_883), .Y(n_987) );
AND2x2_ASAP7_75t_L g998 ( .A(n_837), .B(n_989), .Y(n_998) );
AND2x2_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_854), .Y(n_841) );
AND2x2_ASAP7_75t_L g885 ( .A(n_842), .B(n_886), .Y(n_885) );
AND2x2_ASAP7_75t_L g898 ( .A(n_842), .B(n_899), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_842), .B(n_924), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g939 ( .A(n_842), .B(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_842), .B(n_945), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_842), .B(n_905), .Y(n_1012) );
NOR2x1p5_ASAP7_75t_L g1020 ( .A(n_842), .B(n_1021), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1031 ( .A(n_842), .B(n_892), .Y(n_1031) );
INVx1_ASAP7_75t_L g1040 ( .A(n_842), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_842), .B(n_895), .Y(n_1048) );
CKINVDCx6p67_ASAP7_75t_R g842 ( .A(n_843), .Y(n_842) );
AND2x2_ASAP7_75t_L g891 ( .A(n_843), .B(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g908 ( .A(n_843), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_843), .B(n_929), .Y(n_928) );
AND2x2_ASAP7_75t_L g964 ( .A(n_843), .B(n_883), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_843), .B(n_855), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_843), .B(n_969), .Y(n_968) );
AND2x2_ASAP7_75t_L g989 ( .A(n_843), .B(n_905), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_843), .B(n_886), .Y(n_1055) );
OR2x6_ASAP7_75t_SL g843 ( .A(n_844), .B(n_849), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_847), .B2(n_848), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_847), .A2(n_857), .B1(n_859), .B2(n_860), .Y(n_856) );
OAI22xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B1(n_852), .B2(n_853), .Y(n_849) );
OAI221xp5_ASAP7_75t_L g937 ( .A1(n_854), .A2(n_938), .B1(n_944), .B2(n_946), .C(n_947), .Y(n_937) );
INVx1_ASAP7_75t_L g957 ( .A(n_854), .Y(n_957) );
OR2x2_ASAP7_75t_L g854 ( .A(n_855), .B(n_868), .Y(n_854) );
AND2x2_ASAP7_75t_L g888 ( .A(n_855), .B(n_889), .Y(n_888) );
INVx3_ASAP7_75t_L g892 ( .A(n_855), .Y(n_892) );
INVx2_ASAP7_75t_L g903 ( .A(n_855), .Y(n_903) );
AND2x2_ASAP7_75t_L g945 ( .A(n_855), .B(n_868), .Y(n_945) );
OR2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_861), .Y(n_855) );
INVx3_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_865), .B2(n_866), .Y(n_861) );
INVx3_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_867), .Y(n_1057) );
INVx2_ASAP7_75t_L g889 ( .A(n_868), .Y(n_889) );
AND2x2_ASAP7_75t_L g973 ( .A(n_868), .B(n_892), .Y(n_973) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_868), .B(n_915), .Y(n_1037) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_871), .Y(n_868) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_882), .B(n_887), .C(n_890), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
AND2x2_ASAP7_75t_SL g893 ( .A(n_876), .B(n_886), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_876), .B(n_907), .Y(n_946) );
AND2x2_ASAP7_75t_L g990 ( .A(n_876), .B(n_898), .Y(n_990) );
AND2x2_ASAP7_75t_L g876 ( .A(n_877), .B(n_881), .Y(n_876) );
INVx1_ASAP7_75t_L g884 ( .A(n_877), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_880), .Y(n_877) );
AND2x2_ASAP7_75t_L g883 ( .A(n_881), .B(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_881), .B(n_899), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_881), .B(n_898), .Y(n_1034) );
INVx1_ASAP7_75t_L g955 ( .A(n_882), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_885), .Y(n_882) );
AND2x2_ASAP7_75t_L g897 ( .A(n_883), .B(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g953 ( .A(n_883), .Y(n_953) );
O2A1O1Ixp33_ASAP7_75t_L g983 ( .A1(n_883), .A2(n_984), .B(n_985), .C(n_986), .Y(n_983) );
OAI211xp5_ASAP7_75t_L g1009 ( .A1(n_883), .A2(n_1010), .B(n_1011), .C(n_1012), .Y(n_1009) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_884), .B(n_899), .Y(n_929) );
AND2x2_ASAP7_75t_L g943 ( .A(n_884), .B(n_899), .Y(n_943) );
AND2x2_ASAP7_75t_L g969 ( .A(n_884), .B(n_886), .Y(n_969) );
INVx1_ASAP7_75t_L g1008 ( .A(n_884), .Y(n_1008) );
AND2x2_ASAP7_75t_L g924 ( .A(n_886), .B(n_925), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_886), .B(n_905), .Y(n_952) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_886), .B(n_935), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_886), .B(n_964), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_887), .B(n_911), .Y(n_994) );
AOI21xp33_ASAP7_75t_L g1033 ( .A1(n_887), .A2(n_906), .B(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_888), .B(n_907), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_888), .B(n_924), .Y(n_1051) );
INVx3_ASAP7_75t_L g895 ( .A(n_889), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_889), .B(n_915), .Y(n_960) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_889), .B(n_914), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_889), .B(n_915), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_893), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g1011 ( .A(n_891), .B(n_925), .Y(n_1011) );
INVx1_ASAP7_75t_L g927 ( .A(n_892), .Y(n_927) );
AOI21xp33_ASAP7_75t_L g986 ( .A1(n_892), .A2(n_942), .B(n_987), .Y(n_986) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_892), .B(n_913), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_892), .B(n_914), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_893), .B(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g1046 ( .A(n_893), .Y(n_1046) );
AOI32xp33_ASAP7_75t_SL g894 ( .A1(n_895), .A2(n_896), .A3(n_901), .B1(n_906), .B2(n_909), .Y(n_894) );
INVx3_ASAP7_75t_L g909 ( .A(n_895), .Y(n_909) );
AOI31xp33_ASAP7_75t_L g979 ( .A1(n_895), .A2(n_980), .A3(n_991), .B(n_992), .Y(n_979) );
INVx1_ASAP7_75t_L g1049 ( .A(n_895), .Y(n_1049) );
OAI211xp5_ASAP7_75t_L g1050 ( .A1(n_896), .A2(n_961), .B(n_1051), .C(n_1052), .Y(n_1050) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
AND2x2_ASAP7_75t_L g904 ( .A(n_898), .B(n_905), .Y(n_904) );
INVxp67_ASAP7_75t_SL g1010 ( .A(n_898), .Y(n_1010) );
AND2x2_ASAP7_75t_L g963 ( .A(n_899), .B(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
INVx1_ASAP7_75t_L g921 ( .A(n_901), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_904), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g1052 ( .A(n_902), .B(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx2_ASAP7_75t_L g962 ( .A(n_903), .Y(n_962) );
INVx1_ASAP7_75t_L g935 ( .A(n_905), .Y(n_935) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_905), .B(n_1054), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_907), .B(n_943), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_907), .B(n_973), .Y(n_1005) );
INVx3_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g948 ( .A(n_909), .B(n_930), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_909), .A2(n_956), .B1(n_997), .B2(n_998), .Y(n_996) );
AOI32xp33_ASAP7_75t_L g1003 ( .A1(n_910), .A2(n_1004), .A3(n_1006), .B1(n_1009), .B2(n_1013), .Y(n_1003) );
INVx3_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g992 ( .A1(n_911), .A2(n_981), .B1(n_993), .B2(n_1002), .Y(n_992) );
INVx3_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx3_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_914), .B(n_950), .Y(n_991) );
NOR3xp33_ASAP7_75t_L g1029 ( .A(n_914), .B(n_1030), .C(n_1032), .Y(n_1029) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_914), .B(n_950), .Y(n_1042) );
INVx3_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
AND2x2_ASAP7_75t_L g956 ( .A(n_915), .B(n_957), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_915), .B(n_945), .Y(n_1027) );
AND2x4_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .Y(n_915) );
INVx2_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
OAI321xp33_ASAP7_75t_L g920 ( .A1(n_921), .A2(n_922), .A3(n_926), .B1(n_934), .B2(n_937), .C(n_948), .Y(n_920) );
AOI221xp5_ASAP7_75t_L g1043 ( .A1(n_922), .A2(n_1044), .B1(n_1047), .B2(n_1049), .C(n_1050), .Y(n_1043) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_925), .B(n_1026), .Y(n_1025) );
INVx1_ASAP7_75t_L g1032 ( .A(n_925), .Y(n_1032) );
OAI21xp33_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B(n_930), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_929), .B(n_967), .Y(n_966) );
CKINVDCx16_ASAP7_75t_R g947 ( .A(n_930), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_930), .B(n_972), .Y(n_971) );
AOI221xp5_ASAP7_75t_SL g999 ( .A1(n_930), .A2(n_959), .B1(n_977), .B2(n_990), .C(n_1000), .Y(n_999) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx3_ASAP7_75t_L g950 ( .A(n_931), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_939), .B(n_941), .Y(n_938) );
INVx1_ASAP7_75t_L g982 ( .A(n_939), .Y(n_982) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
OAI21xp33_ASAP7_75t_L g1035 ( .A1(n_942), .A2(n_1036), .B(n_1038), .Y(n_1035) );
INVx1_ASAP7_75t_L g1045 ( .A(n_943), .Y(n_1045) );
OAI211xp5_ASAP7_75t_L g981 ( .A1(n_944), .A2(n_982), .B(n_983), .C(n_988), .Y(n_981) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
O2A1O1Ixp33_ASAP7_75t_L g1016 ( .A1(n_947), .A2(n_1017), .B(n_1019), .C(n_1020), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g965 ( .A1(n_948), .A2(n_966), .B1(n_968), .B2(n_970), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_951), .B1(n_955), .B2(n_956), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g1022 ( .A1(n_950), .A2(n_1023), .B1(n_1042), .B2(n_1043), .Y(n_1022) );
AOI21xp33_ASAP7_75t_L g951 ( .A1(n_952), .A2(n_953), .B(n_954), .Y(n_951) );
INVx1_ASAP7_75t_L g1041 ( .A(n_952), .Y(n_1041) );
INVx1_ASAP7_75t_L g985 ( .A(n_954), .Y(n_985) );
INVx1_ASAP7_75t_L g978 ( .A(n_956), .Y(n_978) );
O2A1O1Ixp33_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_961), .B(n_963), .C(n_965), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
OAI211xp5_ASAP7_75t_L g1024 ( .A1(n_960), .A2(n_987), .B(n_1025), .C(n_1028), .Y(n_1024) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVxp67_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_973), .A2(n_989), .B(n_990), .Y(n_988) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
INVxp67_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
A2O1A1Ixp33_ASAP7_75t_L g1038 ( .A1(n_984), .A2(n_1000), .B(n_1039), .C(n_1041), .Y(n_1038) );
OAI211xp5_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_995), .B(n_996), .C(n_999), .Y(n_993) );
INVx1_ASAP7_75t_L g1015 ( .A(n_998), .Y(n_1015) );
INVx1_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
NAND3xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1015), .C(n_1016), .Y(n_1002) );
INVxp67_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
NOR3xp33_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1033), .C(n_1035), .Y(n_1023) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
CKINVDCx14_ASAP7_75t_R g1039 ( .A(n_1040), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1046), .Y(n_1044) );
INVx1_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g1056 ( .A(n_1057), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
XOR2x2_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1076), .Y(n_1060) );
NOR2x1_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1067), .Y(n_1061) );
NAND4xp25_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .C(n_1065), .D(n_1066), .Y(n_1062) );
NAND4xp25_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1070), .C(n_1071), .D(n_1074), .Y(n_1067) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1078), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
HB1xp67_ASAP7_75t_SL g1086 ( .A(n_1087), .Y(n_1086) );
NOR3xp33_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1091), .C(n_1095), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1090), .Y(n_1088) );
NAND2xp5_ASAP7_75t_SL g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
NAND4xp25_ASAP7_75t_SL g1095 ( .A(n_1096), .B(n_1097), .C(n_1100), .D(n_1102), .Y(n_1095) );
BUFx2_ASAP7_75t_SL g1103 ( .A(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
endmodule