module fake_jpeg_28869_n_115 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_115);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_3),
.B(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_1),
.Y(n_49)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_39),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_17),
.A2(n_1),
.B1(n_10),
.B2(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_52),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_56),
.Y(n_59)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_22),
.B1(n_21),
.B2(n_16),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_12),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_14),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_21),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_65),
.B1(n_69),
.B2(n_44),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_16),
.Y(n_60)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_68),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_51),
.B(n_48),
.Y(n_62)
);

XNOR2x1_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_47),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_28),
.B(n_23),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

BUFx12f_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_66),
.B(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_72),
.Y(n_83)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_23),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_38),
.B(n_53),
.C(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_80),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_73),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_90),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_70),
.B1(n_61),
.B2(n_72),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_84),
.B(n_78),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_91),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_85),
.C(n_77),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_77),
.C(n_74),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_96),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

BUFx12f_ASAP7_75t_SL g103 ( 
.A(n_94),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_88),
.B1(n_99),
.B2(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_102),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_110),
.A2(n_106),
.B(n_107),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_111),
.C(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_100),
.Y(n_115)
);


endmodule