module fake_jpeg_27184_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx8_ASAP7_75t_SL g15 ( 
.A(n_10),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_23),
.Y(n_35)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

AO22x2_ASAP7_75t_L g32 ( 
.A1(n_15),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_14),
.B1(n_22),
.B2(n_15),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_42),
.B1(n_33),
.B2(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_40),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_22),
.B1(n_13),
.B2(n_19),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_57),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_60),
.B1(n_39),
.B2(n_41),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_31),
.B(n_25),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_53),
.B(n_18),
.Y(n_72)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_58),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_59),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_2),
.B(n_3),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_25),
.C(n_21),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_56),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_21),
.C(n_12),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_35),
.B(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_40),
.B1(n_34),
.B2(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_70),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_38),
.C(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_38),
.C(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_67),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_52),
.B1(n_60),
.B2(n_39),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_74),
.B1(n_57),
.B2(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_43),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_12),
.B(n_18),
.C(n_13),
.Y(n_69)
);

XOR2x1_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_17),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_87),
.B1(n_41),
.B2(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_59),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_90),
.B(n_69),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_67),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_20),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_44),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_41),
.B1(n_36),
.B2(n_37),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_95),
.B(n_90),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_66),
.C(n_70),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_86),
.C(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_65),
.B(n_8),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_44),
.Y(n_97)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_84),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_89),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_104),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_91),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_84),
.C(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_97),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_77),
.B(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_113),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_104),
.B(n_98),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_108),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_105),
.B(n_106),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_37),
.C(n_65),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_95),
.B1(n_99),
.B2(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_118),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_101),
.A3(n_93),
.B1(n_87),
.B2(n_20),
.C(n_81),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_36),
.C(n_41),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_120),
.A3(n_20),
.B1(n_9),
.B2(n_10),
.C1(n_5),
.C2(n_8),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_126),
.B(n_8),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_129),
.B(n_9),
.Y(n_130)
);

AOI21x1_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_9),
.B(n_11),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_11),
.Y(n_131)
);


endmodule