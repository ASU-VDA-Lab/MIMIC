module fake_jpeg_23101_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx3_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_21),
.A2(n_19),
.B1(n_15),
.B2(n_20),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_13),
.C(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_26),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

NAND2xp67_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_39),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_3),
.B1(n_9),
.B2(n_38),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_15),
.B1(n_11),
.B2(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_49),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_31),
.Y(n_57)
);

AO22x2_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_29),
.C(n_34),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_31),
.C(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_48),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_48),
.B1(n_42),
.B2(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_61),
.B(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_49),
.B1(n_54),
.B2(n_52),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_63),
.A2(n_64),
.B(n_62),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_65),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_58),
.B(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_36),
.Y(n_72)
);


endmodule