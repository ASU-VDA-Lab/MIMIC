module fake_ariane_3238_n_7517 (n_913, n_1681, n_1486, n_1507, n_589, n_1174, n_1469, n_691, n_1353, n_1355, n_423, n_1383, n_603, n_373, n_1250, n_1169, n_789, n_850, n_610, n_245, n_1713, n_96, n_319, n_49, n_1436, n_690, n_416, n_1109, n_1430, n_525, n_187, n_1463, n_1238, n_1515, n_817, n_1837, n_924, n_781, n_1566, n_189, n_717, n_72, n_952, n_864, n_1096, n_1379, n_57, n_1706, n_117, n_524, n_1214, n_634, n_1839, n_1246, n_1138, n_214, n_1853, n_764, n_1503, n_462, n_1196, n_1181, n_32, n_410, n_1187, n_1131, n_1225, n_737, n_137, n_1298, n_1745, n_1366, n_232, n_52, n_568, n_1088, n_77, n_1424, n_766, n_1835, n_1457, n_377, n_1682, n_1836, n_520, n_870, n_1453, n_279, n_945, n_958, n_813, n_419, n_146, n_270, n_338, n_995, n_285, n_1184, n_202, n_1535, n_500, n_665, n_754, n_903, n_871, n_1073, n_239, n_402, n_1277, n_1746, n_54, n_829, n_1761, n_1062, n_339, n_738, n_1690, n_672, n_740, n_1283, n_167, n_1736, n_1018, n_69, n_259, n_953, n_1364, n_143, n_1224, n_1425, n_625, n_557, n_1107, n_1688, n_989, n_242, n_645, n_331, n_559, n_267, n_495, n_350, n_381, n_795, n_721, n_1084, n_1718, n_1276, n_200, n_1428, n_1284, n_1241, n_821, n_561, n_770, n_1514, n_1528, n_507, n_486, n_901, n_569, n_1145, n_971, n_787, n_1650, n_31, n_1519, n_1195, n_1522, n_518, n_1207, n_222, n_786, n_1404, n_868, n_1847, n_1542, n_1314, n_1512, n_1539, n_884, n_1851, n_1415, n_1034, n_1652, n_1676, n_1085, n_277, n_1636, n_432, n_293, n_823, n_620, n_93, n_1074, n_859, n_1765, n_108, n_587, n_693, n_863, n_303, n_1254, n_929, n_206, n_352, n_899, n_1703, n_611, n_1295, n_1850, n_238, n_365, n_1013, n_1495, n_1637, n_136, n_334, n_192, n_661, n_1751, n_300, n_533, n_104, n_438, n_1560, n_1654, n_1548, n_16, n_1811, n_440, n_273, n_1396, n_1230, n_612, n_333, n_1840, n_376, n_512, n_1597, n_1771, n_1544, n_579, n_844, n_1012, n_1267, n_1354, n_1790, n_149, n_1213, n_237, n_780, n_1021, n_1443, n_491, n_1465, n_1595, n_1142, n_1140, n_705, n_570, n_260, n_942, n_1437, n_7, n_1378, n_461, n_1121, n_1416, n_209, n_490, n_1461, n_17, n_1391, n_225, n_1599, n_1876, n_1006, n_1830, n_575, n_546, n_503, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_1669, n_1675, n_676, n_42, n_1838, n_1594, n_680, n_287, n_1716, n_302, n_1872, n_380, n_1585, n_1432, n_94, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_1590, n_1351, n_1274, n_257, n_652, n_1819, n_475, n_135, n_947, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_1442, n_482, n_798, n_577, n_1833, n_407, n_1691, n_27, n_916, n_1386, n_912, n_460, n_1555, n_1842, n_366, n_762, n_1253, n_1468, n_1661, n_555, n_804, n_1656, n_1382, n_966, n_992, n_955, n_1182, n_794, n_78, n_1692, n_1562, n_514, n_418, n_1376, n_513, n_288, n_179, n_1292, n_1178, n_1435, n_1750, n_1026, n_1506, n_1610, n_306, n_92, n_203, n_436, n_150, n_324, n_669, n_931, n_1491, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_1418, n_746, n_1357, n_292, n_1079, n_1787, n_1389, n_615, n_1139, n_76, n_517, n_1312, n_1717, n_0, n_1812, n_824, n_428, n_159, n_892, n_1880, n_959, n_30, n_1399, n_1101, n_1567, n_1343, n_563, n_1855, n_144, n_990, n_1623, n_867, n_1226, n_944, n_749, n_1780, n_815, n_542, n_1340, n_470, n_1240, n_1087, n_632, n_477, n_650, n_425, n_1433, n_1825, n_1155, n_1071, n_712, n_976, n_909, n_1392, n_767, n_1832, n_1841, n_1680, n_964, n_1627, n_382, n_489, n_80, n_251, n_974, n_506, n_1731, n_799, n_1147, n_397, n_471, n_351, n_965, n_155, n_934, n_1447, n_1220, n_356, n_698, n_1674, n_124, n_307, n_1209, n_1020, n_1563, n_646, n_1633, n_34, n_404, n_172, n_1058, n_347, n_1042, n_183, n_1234, n_479, n_1578, n_1455, n_299, n_836, n_1279, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_1568, n_20, n_1483, n_1363, n_367, n_1111, n_970, n_1689, n_713, n_1255, n_1646, n_598, n_345, n_1237, n_927, n_261, n_1095, n_1728, n_370, n_706, n_286, n_1401, n_1419, n_1531, n_776, n_424, n_1651, n_85, n_130, n_1387, n_466, n_1263, n_346, n_1817, n_348, n_552, n_670, n_1826, n_379, n_138, n_162, n_264, n_441, n_1032, n_1217, n_1496, n_637, n_1592, n_73, n_327, n_1259, n_1177, n_1231, n_980, n_1618, n_1869, n_1743, n_905, n_207, n_720, n_926, n_41, n_194, n_1802, n_1163, n_186, n_1795, n_1384, n_145, n_1868, n_59, n_1501, n_1173, n_1068, n_1198, n_1570, n_487, n_1518, n_1456, n_90, n_1879, n_1648, n_1413, n_855, n_158, n_808, n_1365, n_553, n_1439, n_814, n_578, n_1665, n_1287, n_405, n_1611, n_120, n_320, n_1414, n_1134, n_1484, n_647, n_1423, n_481, n_600, n_1053, n_1609, n_529, n_502, n_218, n_1467, n_247, n_1828, n_1798, n_1304, n_1608, n_1744, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1349, n_1709, n_1061, n_326, n_681, n_227, n_874, n_1278, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_1726, n_545, n_1015, n_1377, n_1162, n_536, n_1614, n_325, n_1740, n_1602, n_688, n_636, n_427, n_1098, n_1490, n_442, n_777, n_1553, n_1080, n_920, n_1760, n_1086, n_1092, n_986, n_1104, n_729, n_887, n_1122, n_1205, n_1408, n_163, n_1693, n_1132, n_390, n_1156, n_501, n_314, n_1823, n_1120, n_1202, n_627, n_1188, n_1498, n_1371, n_233, n_957, n_388, n_1402, n_1242, n_1607, n_1489, n_1218, n_221, n_321, n_86, n_1586, n_861, n_1543, n_1431, n_877, n_1119, n_1863, n_1763, n_1666, n_1500, n_616, n_1055, n_1395, n_1346, n_1189, n_1089, n_281, n_1859, n_262, n_1502, n_1523, n_1478, n_735, n_297, n_1005, n_527, n_46, n_84, n_1294, n_1667, n_845, n_888, n_1649, n_1677, n_1297, n_178, n_551, n_417, n_1708, n_70, n_343, n_1222, n_1844, n_582, n_755, n_1097, n_1219, n_1711, n_710, n_534, n_1791, n_1460, n_1239, n_278, n_560, n_890, n_842, n_148, n_451, n_745, n_1741, n_1572, n_1793, n_61, n_742, n_1081, n_1373, n_1388, n_1266, n_1540, n_1719, n_769, n_1797, n_13, n_1753, n_1372, n_476, n_832, n_55, n_535, n_744, n_982, n_1800, n_915, n_215, n_1075, n_454, n_298, n_1331, n_1529, n_1227, n_655, n_1734, n_1860, n_403, n_1007, n_1580, n_1319, n_657, n_837, n_812, n_606, n_951, n_862, n_1700, n_659, n_1332, n_509, n_1854, n_666, n_1747, n_430, n_1206, n_1729, n_722, n_1508, n_1532, n_1171, n_1030, n_785, n_1309, n_999, n_1766, n_1338, n_1342, n_456, n_1867, n_852, n_1394, n_704, n_1060, n_1044, n_1714, n_521, n_873, n_1301, n_1748, n_1243, n_1400, n_342, n_1466, n_1513, n_1527, n_358, n_1783, n_608, n_1538, n_1037, n_1329, n_317, n_1545, n_134, n_1257, n_1480, n_1668, n_1878, n_1605, n_1078, n_266, n_157, n_1161, n_811, n_624, n_791, n_876, n_618, n_1191, n_736, n_1025, n_1215, n_241, n_1449, n_687, n_797, n_1786, n_480, n_1327, n_1475, n_211, n_642, n_1804, n_97, n_408, n_1406, n_595, n_1405, n_602, n_1757, n_592, n_1499, n_854, n_1318, n_393, n_1632, n_1769, n_474, n_805, n_295, n_1658, n_190, n_1072, n_695, n_1526, n_1305, n_64, n_180, n_730, n_386, n_1596, n_1281, n_516, n_1137, n_1873, n_1258, n_197, n_640, n_463, n_1476, n_1524, n_1733, n_1856, n_943, n_1118, n_678, n_651, n_1874, n_1293, n_961, n_469, n_1046, n_1807, n_726, n_1123, n_1657, n_878, n_1784, n_771, n_1321, n_752, n_71, n_1488, n_985, n_421, n_1330, n_906, n_1180, n_1697, n_283, n_806, n_1350, n_1556, n_649, n_1561, n_374, n_1352, n_1824, n_643, n_1492, n_226, n_1441, n_1822, n_682, n_36, n_1616, n_819, n_586, n_1324, n_1429, n_1778, n_1776, n_686, n_605, n_1154, n_584, n_1557, n_1759, n_1829, n_1130, n_1450, n_349, n_756, n_1016, n_1149, n_1505, n_979, n_1642, n_2, n_1815, n_897, n_949, n_1493, n_515, n_807, n_891, n_885, n_1659, n_198, n_1864, n_1208, n_396, n_802, n_23, n_1151, n_554, n_960, n_1256, n_87, n_714, n_790, n_354, n_140, n_725, n_1577, n_151, n_1448, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_1852, n_801, n_1286, n_818, n_1685, n_779, n_594, n_1877, n_1397, n_35, n_1052, n_272, n_1333, n_1306, n_1849, n_833, n_1426, n_879, n_1117, n_38, n_422, n_1269, n_1303, n_1547, n_1438, n_1541, n_597, n_75, n_1047, n_95, n_1472, n_1593, n_1050, n_566, n_152, n_169, n_106, n_1201, n_1288, n_173, n_858, n_1185, n_335, n_1035, n_1143, n_344, n_426, n_433, n_398, n_62, n_210, n_1090, n_1367, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1565, n_1192, n_128, n_224, n_82, n_894, n_1380, n_1624, n_1801, n_420, n_1291, n_562, n_748, n_510, n_1045, n_256, n_1160, n_1882, n_1023, n_1881, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_467, n_1511, n_1422, n_644, n_1197, n_276, n_497, n_1165, n_1641, n_168, n_81, n_538, n_1517, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_1307, n_1128, n_1671, n_1417, n_1048, n_775, n_667, n_1049, n_14, n_869, n_141, n_846, n_1398, n_1356, n_1341, n_1504, n_1773, n_1440, n_1370, n_1603, n_305, n_312, n_56, n_60, n_728, n_413, n_715, n_889, n_1066, n_1549, n_935, n_685, n_911, n_361, n_89, n_623, n_1712, n_1403, n_1065, n_453, n_1534, n_74, n_810, n_19, n_40, n_1290, n_181, n_617, n_543, n_1362, n_1559, n_236, n_601, n_683, n_565, n_628, n_1300, n_743, n_1194, n_1647, n_1546, n_1420, n_907, n_1454, n_660, n_464, n_962, n_941, n_1210, n_847, n_747, n_1622, n_1135, n_918, n_107, n_639, n_452, n_673, n_1038, n_414, n_571, n_1521, n_1694, n_6, n_284, n_593, n_1695, n_1164, n_37, n_58, n_609, n_1193, n_1345, n_613, n_1022, n_1336, n_1033, n_1774, n_409, n_171, n_519, n_384, n_1166, n_1056, n_526, n_1767, n_1040, n_674, n_1158, n_316, n_125, n_1444, n_1803, n_820, n_1749, n_43, n_872, n_1653, n_254, n_1157, n_1584, n_234, n_848, n_1664, n_280, n_629, n_1739, n_161, n_1814, n_532, n_1789, n_763, n_99, n_540, n_216, n_692, n_5, n_1857, n_984, n_1687, n_223, n_1552, n_750, n_834, n_1612, n_800, n_1816, n_1756, n_1606, n_395, n_621, n_1587, n_213, n_1772, n_67, n_1014, n_724, n_1427, n_1481, n_493, n_1311, n_1589, n_114, n_1100, n_585, n_875, n_1617, n_827, n_697, n_622, n_1626, n_1335, n_1715, n_296, n_880, n_793, n_1175, n_132, n_751, n_1027, n_1070, n_1621, n_739, n_1485, n_1028, n_1221, n_530, n_1785, n_792, n_1262, n_580, n_1579, n_494, n_434, n_975, n_229, n_394, n_923, n_1645, n_1124, n_1381, n_1494, n_932, n_1183, n_1326, n_1805, n_981, n_1110, n_1758, n_243, n_1407, n_185, n_1204, n_1554, n_994, n_1360, n_973, n_268, n_972, n_164, n_184, n_856, n_1248, n_1176, n_1564, n_1054, n_508, n_118, n_121, n_1679, n_1858, n_353, n_1678, n_1482, n_1361, n_1601, n_1057, n_191, n_1834, n_978, n_1011, n_1520, n_1509, n_828, n_322, n_1411, n_1359, n_558, n_1721, n_116, n_39, n_653, n_1445, n_1317, n_783, n_556, n_1127, n_170, n_1536, n_1471, n_160, n_119, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_987, n_936, n_1620, n_1385, n_1525, n_541, n_499, n_1775, n_788, n_12, n_908, n_1036, n_341, n_1270, n_109, n_1167, n_1272, n_549, n_591, n_969, n_919, n_1663, n_50, n_1625, n_318, n_1458, n_103, n_244, n_679, n_1630, n_220, n_663, n_1720, n_443, n_1412, n_1738, n_1550, n_528, n_1358, n_1200, n_387, n_406, n_826, n_139, n_1735, n_1788, n_391, n_940, n_1537, n_1077, n_607, n_956, n_445, n_765, n_1809, n_1843, n_122, n_1268, n_385, n_917, n_1271, n_372, n_15, n_1530, n_631, n_399, n_1170, n_1261, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1323, n_1462, n_1064, n_633, n_900, n_1446, n_1282, n_1701, n_1093, n_1551, n_1755, n_1285, n_193, n_733, n_761, n_731, n_336, n_1813, n_315, n_311, n_1452, n_1573, n_8, n_668, n_758, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_1322, n_1473, n_835, n_446, n_1076, n_1348, n_753, n_1770, n_701, n_1003, n_1125, n_1710, n_1865, n_309, n_1344, n_115, n_1390, n_401, n_485, n_1792, n_504, n_483, n_435, n_1141, n_1629, n_291, n_1640, n_822, n_1094, n_840, n_1459, n_1510, n_1099, n_839, n_79, n_1754, n_3, n_759, n_567, n_91, n_240, n_369, n_1727, n_44, n_1575, n_1848, n_1172, n_614, n_1212, n_831, n_778, n_48, n_1619, n_188, n_323, n_550, n_1315, n_1660, n_997, n_635, n_694, n_1643, n_1320, n_1113, n_248, n_1152, n_1845, n_921, n_1615, n_1236, n_228, n_1265, n_1576, n_1470, n_671, n_1533, n_1806, n_1, n_1409, n_1148, n_1588, n_1684, n_1673, n_1334, n_654, n_1275, n_488, n_904, n_505, n_88, n_1696, n_498, n_1875, n_1059, n_684, n_1039, n_539, n_1150, n_977, n_449, n_392, n_1628, n_1289, n_1831, n_1497, n_1866, n_459, n_1136, n_1782, n_458, n_1190, n_1600, n_1144, n_383, n_838, n_1558, n_1316, n_175, n_950, n_1017, n_711, n_734, n_723, n_1393, n_658, n_630, n_1369, n_53, n_362, n_310, n_1781, n_709, n_24, n_809, n_1686, n_235, n_881, n_1019, n_1477, n_1777, n_662, n_641, n_910, n_290, n_741, n_939, n_1410, n_371, n_199, n_217, n_1114, n_1325, n_1742, n_708, n_308, n_1223, n_201, n_1768, n_572, n_1199, n_865, n_10, n_1273, n_1041, n_993, n_1862, n_948, n_922, n_1004, n_1810, n_448, n_1347, n_860, n_1043, n_255, n_450, n_1764, n_896, n_1737, n_1479, n_1613, n_902, n_1031, n_1723, n_1638, n_853, n_716, n_1571, n_1698, n_196, n_1337, n_774, n_933, n_1779, n_596, n_954, n_1168, n_1821, n_219, n_1310, n_231, n_656, n_492, n_574, n_252, n_664, n_1591, n_1229, n_1683, n_68, n_1732, n_415, n_63, n_1280, n_544, n_1516, n_1186, n_1705, n_599, n_768, n_1091, n_537, n_1063, n_25, n_991, n_83, n_389, n_1724, n_1670, n_1707, n_1799, n_1126, n_195, n_1846, n_938, n_1328, n_895, n_110, n_304, n_1639, n_583, n_1302, n_1000, n_313, n_626, n_378, n_1581, n_98, n_946, n_757, n_375, n_113, n_1655, n_1818, n_33, n_1146, n_1634, n_1203, n_998, n_1699, n_1598, n_472, n_937, n_1474, n_265, n_1583, n_1604, n_208, n_1631, n_1702, n_156, n_174, n_275, n_100, n_1794, n_1375, n_147, n_204, n_1232, n_996, n_1211, n_1368, n_963, n_1264, n_51, n_1082, n_1725, n_496, n_1827, n_866, n_26, n_246, n_925, n_1752, n_1313, n_1001, n_1722, n_1115, n_1339, n_1002, n_1644, n_105, n_1051, n_719, n_131, n_263, n_1102, n_360, n_1129, n_1252, n_250, n_1464, n_1296, n_773, n_165, n_1010, n_882, n_1249, n_101, n_803, n_1871, n_329, n_718, n_1434, n_340, n_1569, n_289, n_9, n_112, n_45, n_548, n_523, n_1662, n_457, n_1299, n_1870, n_177, n_782, n_364, n_258, n_431, n_1861, n_1228, n_1244, n_1796, n_411, n_484, n_849, n_22, n_1820, n_29, n_357, n_412, n_1251, n_447, n_1421, n_1762, n_1233, n_1808, n_1574, n_1672, n_1635, n_1704, n_893, n_1582, n_841, n_886, n_1069, n_359, n_1308, n_573, n_796, n_127, n_531, n_1730, n_1374, n_1451, n_1487, n_675, n_7517);

input n_913;
input n_1681;
input n_1486;
input n_1507;
input n_589;
input n_1174;
input n_1469;
input n_691;
input n_1353;
input n_1355;
input n_423;
input n_1383;
input n_603;
input n_373;
input n_1250;
input n_1169;
input n_789;
input n_850;
input n_610;
input n_245;
input n_1713;
input n_96;
input n_319;
input n_49;
input n_1436;
input n_690;
input n_416;
input n_1109;
input n_1430;
input n_525;
input n_187;
input n_1463;
input n_1238;
input n_1515;
input n_817;
input n_1837;
input n_924;
input n_781;
input n_1566;
input n_189;
input n_717;
input n_72;
input n_952;
input n_864;
input n_1096;
input n_1379;
input n_57;
input n_1706;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1839;
input n_1246;
input n_1138;
input n_214;
input n_1853;
input n_764;
input n_1503;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_410;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_1298;
input n_1745;
input n_1366;
input n_232;
input n_52;
input n_568;
input n_1088;
input n_77;
input n_1424;
input n_766;
input n_1835;
input n_1457;
input n_377;
input n_1682;
input n_1836;
input n_520;
input n_870;
input n_1453;
input n_279;
input n_945;
input n_958;
input n_813;
input n_419;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1184;
input n_202;
input n_1535;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_1073;
input n_239;
input n_402;
input n_1277;
input n_1746;
input n_54;
input n_829;
input n_1761;
input n_1062;
input n_339;
input n_738;
input n_1690;
input n_672;
input n_740;
input n_1283;
input n_167;
input n_1736;
input n_1018;
input n_69;
input n_259;
input n_953;
input n_1364;
input n_143;
input n_1224;
input n_1425;
input n_625;
input n_557;
input n_1107;
input n_1688;
input n_989;
input n_242;
input n_645;
input n_331;
input n_559;
input n_267;
input n_495;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_1718;
input n_1276;
input n_200;
input n_1428;
input n_1284;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_1514;
input n_1528;
input n_507;
input n_486;
input n_901;
input n_569;
input n_1145;
input n_971;
input n_787;
input n_1650;
input n_31;
input n_1519;
input n_1195;
input n_1522;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_1404;
input n_868;
input n_1847;
input n_1542;
input n_1314;
input n_1512;
input n_1539;
input n_884;
input n_1851;
input n_1415;
input n_1034;
input n_1652;
input n_1676;
input n_1085;
input n_277;
input n_1636;
input n_432;
input n_293;
input n_823;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_1765;
input n_108;
input n_587;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_206;
input n_352;
input n_899;
input n_1703;
input n_611;
input n_1295;
input n_1850;
input n_238;
input n_365;
input n_1013;
input n_1495;
input n_1637;
input n_136;
input n_334;
input n_192;
input n_661;
input n_1751;
input n_300;
input n_533;
input n_104;
input n_438;
input n_1560;
input n_1654;
input n_1548;
input n_16;
input n_1811;
input n_440;
input n_273;
input n_1396;
input n_1230;
input n_612;
input n_333;
input n_1840;
input n_376;
input n_512;
input n_1597;
input n_1771;
input n_1544;
input n_579;
input n_844;
input n_1012;
input n_1267;
input n_1354;
input n_1790;
input n_149;
input n_1213;
input n_237;
input n_780;
input n_1021;
input n_1443;
input n_491;
input n_1465;
input n_1595;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_1437;
input n_7;
input n_1378;
input n_461;
input n_1121;
input n_1416;
input n_209;
input n_490;
input n_1461;
input n_17;
input n_1391;
input n_225;
input n_1599;
input n_1876;
input n_1006;
input n_1830;
input n_575;
input n_546;
input n_503;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_1669;
input n_1675;
input n_676;
input n_42;
input n_1838;
input n_1594;
input n_680;
input n_287;
input n_1716;
input n_302;
input n_1872;
input n_380;
input n_1585;
input n_1432;
input n_94;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_1590;
input n_1351;
input n_1274;
input n_257;
input n_652;
input n_1819;
input n_475;
input n_135;
input n_947;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_1442;
input n_482;
input n_798;
input n_577;
input n_1833;
input n_407;
input n_1691;
input n_27;
input n_916;
input n_1386;
input n_912;
input n_460;
input n_1555;
input n_1842;
input n_366;
input n_762;
input n_1253;
input n_1468;
input n_1661;
input n_555;
input n_804;
input n_1656;
input n_1382;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_1692;
input n_1562;
input n_514;
input n_418;
input n_1376;
input n_513;
input n_288;
input n_179;
input n_1292;
input n_1178;
input n_1435;
input n_1750;
input n_1026;
input n_1506;
input n_1610;
input n_306;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_669;
input n_931;
input n_1491;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_1418;
input n_746;
input n_1357;
input n_292;
input n_1079;
input n_1787;
input n_1389;
input n_615;
input n_1139;
input n_76;
input n_517;
input n_1312;
input n_1717;
input n_0;
input n_1812;
input n_824;
input n_428;
input n_159;
input n_892;
input n_1880;
input n_959;
input n_30;
input n_1399;
input n_1101;
input n_1567;
input n_1343;
input n_563;
input n_1855;
input n_144;
input n_990;
input n_1623;
input n_867;
input n_1226;
input n_944;
input n_749;
input n_1780;
input n_815;
input n_542;
input n_1340;
input n_470;
input n_1240;
input n_1087;
input n_632;
input n_477;
input n_650;
input n_425;
input n_1433;
input n_1825;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_1392;
input n_767;
input n_1832;
input n_1841;
input n_1680;
input n_964;
input n_1627;
input n_382;
input n_489;
input n_80;
input n_251;
input n_974;
input n_506;
input n_1731;
input n_799;
input n_1147;
input n_397;
input n_471;
input n_351;
input n_965;
input n_155;
input n_934;
input n_1447;
input n_1220;
input n_356;
input n_698;
input n_1674;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_1563;
input n_646;
input n_1633;
input n_34;
input n_404;
input n_172;
input n_1058;
input n_347;
input n_1042;
input n_183;
input n_1234;
input n_479;
input n_1578;
input n_1455;
input n_299;
input n_836;
input n_1279;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_1568;
input n_20;
input n_1483;
input n_1363;
input n_367;
input n_1111;
input n_970;
input n_1689;
input n_713;
input n_1255;
input n_1646;
input n_598;
input n_345;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_1728;
input n_370;
input n_706;
input n_286;
input n_1401;
input n_1419;
input n_1531;
input n_776;
input n_424;
input n_1651;
input n_85;
input n_130;
input n_1387;
input n_466;
input n_1263;
input n_346;
input n_1817;
input n_348;
input n_552;
input n_670;
input n_1826;
input n_379;
input n_138;
input n_162;
input n_264;
input n_441;
input n_1032;
input n_1217;
input n_1496;
input n_637;
input n_1592;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_980;
input n_1618;
input n_1869;
input n_1743;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_194;
input n_1802;
input n_1163;
input n_186;
input n_1795;
input n_1384;
input n_145;
input n_1868;
input n_59;
input n_1501;
input n_1173;
input n_1068;
input n_1198;
input n_1570;
input n_487;
input n_1518;
input n_1456;
input n_90;
input n_1879;
input n_1648;
input n_1413;
input n_855;
input n_158;
input n_808;
input n_1365;
input n_553;
input n_1439;
input n_814;
input n_578;
input n_1665;
input n_1287;
input n_405;
input n_1611;
input n_120;
input n_320;
input n_1414;
input n_1134;
input n_1484;
input n_647;
input n_1423;
input n_481;
input n_600;
input n_1053;
input n_1609;
input n_529;
input n_502;
input n_218;
input n_1467;
input n_247;
input n_1828;
input n_1798;
input n_1304;
input n_1608;
input n_1744;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1349;
input n_1709;
input n_1061;
input n_326;
input n_681;
input n_227;
input n_874;
input n_1278;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_1726;
input n_545;
input n_1015;
input n_1377;
input n_1162;
input n_536;
input n_1614;
input n_325;
input n_1740;
input n_1602;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_1490;
input n_442;
input n_777;
input n_1553;
input n_1080;
input n_920;
input n_1760;
input n_1086;
input n_1092;
input n_986;
input n_1104;
input n_729;
input n_887;
input n_1122;
input n_1205;
input n_1408;
input n_163;
input n_1693;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_314;
input n_1823;
input n_1120;
input n_1202;
input n_627;
input n_1188;
input n_1498;
input n_1371;
input n_233;
input n_957;
input n_388;
input n_1402;
input n_1242;
input n_1607;
input n_1489;
input n_1218;
input n_221;
input n_321;
input n_86;
input n_1586;
input n_861;
input n_1543;
input n_1431;
input n_877;
input n_1119;
input n_1863;
input n_1763;
input n_1666;
input n_1500;
input n_616;
input n_1055;
input n_1395;
input n_1346;
input n_1189;
input n_1089;
input n_281;
input n_1859;
input n_262;
input n_1502;
input n_1523;
input n_1478;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_46;
input n_84;
input n_1294;
input n_1667;
input n_845;
input n_888;
input n_1649;
input n_1677;
input n_1297;
input n_178;
input n_551;
input n_417;
input n_1708;
input n_70;
input n_343;
input n_1222;
input n_1844;
input n_582;
input n_755;
input n_1097;
input n_1219;
input n_1711;
input n_710;
input n_534;
input n_1791;
input n_1460;
input n_1239;
input n_278;
input n_560;
input n_890;
input n_842;
input n_148;
input n_451;
input n_745;
input n_1741;
input n_1572;
input n_1793;
input n_61;
input n_742;
input n_1081;
input n_1373;
input n_1388;
input n_1266;
input n_1540;
input n_1719;
input n_769;
input n_1797;
input n_13;
input n_1753;
input n_1372;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_982;
input n_1800;
input n_915;
input n_215;
input n_1075;
input n_454;
input n_298;
input n_1331;
input n_1529;
input n_1227;
input n_655;
input n_1734;
input n_1860;
input n_403;
input n_1007;
input n_1580;
input n_1319;
input n_657;
input n_837;
input n_812;
input n_606;
input n_951;
input n_862;
input n_1700;
input n_659;
input n_1332;
input n_509;
input n_1854;
input n_666;
input n_1747;
input n_430;
input n_1206;
input n_1729;
input n_722;
input n_1508;
input n_1532;
input n_1171;
input n_1030;
input n_785;
input n_1309;
input n_999;
input n_1766;
input n_1338;
input n_1342;
input n_456;
input n_1867;
input n_852;
input n_1394;
input n_704;
input n_1060;
input n_1044;
input n_1714;
input n_521;
input n_873;
input n_1301;
input n_1748;
input n_1243;
input n_1400;
input n_342;
input n_1466;
input n_1513;
input n_1527;
input n_358;
input n_1783;
input n_608;
input n_1538;
input n_1037;
input n_1329;
input n_317;
input n_1545;
input n_134;
input n_1257;
input n_1480;
input n_1668;
input n_1878;
input n_1605;
input n_1078;
input n_266;
input n_157;
input n_1161;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_1449;
input n_687;
input n_797;
input n_1786;
input n_480;
input n_1327;
input n_1475;
input n_211;
input n_642;
input n_1804;
input n_97;
input n_408;
input n_1406;
input n_595;
input n_1405;
input n_602;
input n_1757;
input n_592;
input n_1499;
input n_854;
input n_1318;
input n_393;
input n_1632;
input n_1769;
input n_474;
input n_805;
input n_295;
input n_1658;
input n_190;
input n_1072;
input n_695;
input n_1526;
input n_1305;
input n_64;
input n_180;
input n_730;
input n_386;
input n_1596;
input n_1281;
input n_516;
input n_1137;
input n_1873;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_1476;
input n_1524;
input n_1733;
input n_1856;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_1874;
input n_1293;
input n_961;
input n_469;
input n_1046;
input n_1807;
input n_726;
input n_1123;
input n_1657;
input n_878;
input n_1784;
input n_771;
input n_1321;
input n_752;
input n_71;
input n_1488;
input n_985;
input n_421;
input n_1330;
input n_906;
input n_1180;
input n_1697;
input n_283;
input n_806;
input n_1350;
input n_1556;
input n_649;
input n_1561;
input n_374;
input n_1352;
input n_1824;
input n_643;
input n_1492;
input n_226;
input n_1441;
input n_1822;
input n_682;
input n_36;
input n_1616;
input n_819;
input n_586;
input n_1324;
input n_1429;
input n_1778;
input n_1776;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1557;
input n_1759;
input n_1829;
input n_1130;
input n_1450;
input n_349;
input n_756;
input n_1016;
input n_1149;
input n_1505;
input n_979;
input n_1642;
input n_2;
input n_1815;
input n_897;
input n_949;
input n_1493;
input n_515;
input n_807;
input n_891;
input n_885;
input n_1659;
input n_198;
input n_1864;
input n_1208;
input n_396;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_1256;
input n_87;
input n_714;
input n_790;
input n_354;
input n_140;
input n_725;
input n_1577;
input n_151;
input n_1448;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_1852;
input n_801;
input n_1286;
input n_818;
input n_1685;
input n_779;
input n_594;
input n_1877;
input n_1397;
input n_35;
input n_1052;
input n_272;
input n_1333;
input n_1306;
input n_1849;
input n_833;
input n_1426;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_1269;
input n_1303;
input n_1547;
input n_1438;
input n_1541;
input n_597;
input n_75;
input n_1047;
input n_95;
input n_1472;
input n_1593;
input n_1050;
input n_566;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_1288;
input n_173;
input n_858;
input n_1185;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_1367;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1565;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_1380;
input n_1624;
input n_1801;
input n_420;
input n_1291;
input n_562;
input n_748;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1882;
input n_1023;
input n_1881;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_467;
input n_1511;
input n_1422;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_1641;
input n_168;
input n_81;
input n_538;
input n_1517;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_1307;
input n_1128;
input n_1671;
input n_1417;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_14;
input n_869;
input n_141;
input n_846;
input n_1398;
input n_1356;
input n_1341;
input n_1504;
input n_1773;
input n_1440;
input n_1370;
input n_1603;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_715;
input n_889;
input n_1066;
input n_1549;
input n_935;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1712;
input n_1403;
input n_1065;
input n_453;
input n_1534;
input n_74;
input n_810;
input n_19;
input n_40;
input n_1290;
input n_181;
input n_617;
input n_543;
input n_1362;
input n_1559;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_1300;
input n_743;
input n_1194;
input n_1647;
input n_1546;
input n_1420;
input n_907;
input n_1454;
input n_660;
input n_464;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1622;
input n_1135;
input n_918;
input n_107;
input n_639;
input n_452;
input n_673;
input n_1038;
input n_414;
input n_571;
input n_1521;
input n_1694;
input n_6;
input n_284;
input n_593;
input n_1695;
input n_1164;
input n_37;
input n_58;
input n_609;
input n_1193;
input n_1345;
input n_613;
input n_1022;
input n_1336;
input n_1033;
input n_1774;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_526;
input n_1767;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_1444;
input n_1803;
input n_820;
input n_1749;
input n_43;
input n_872;
input n_1653;
input n_254;
input n_1157;
input n_1584;
input n_234;
input n_848;
input n_1664;
input n_280;
input n_629;
input n_1739;
input n_161;
input n_1814;
input n_532;
input n_1789;
input n_763;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_1857;
input n_984;
input n_1687;
input n_223;
input n_1552;
input n_750;
input n_834;
input n_1612;
input n_800;
input n_1816;
input n_1756;
input n_1606;
input n_395;
input n_621;
input n_1587;
input n_213;
input n_1772;
input n_67;
input n_1014;
input n_724;
input n_1427;
input n_1481;
input n_493;
input n_1311;
input n_1589;
input n_114;
input n_1100;
input n_585;
input n_875;
input n_1617;
input n_827;
input n_697;
input n_622;
input n_1626;
input n_1335;
input n_1715;
input n_296;
input n_880;
input n_793;
input n_1175;
input n_132;
input n_751;
input n_1027;
input n_1070;
input n_1621;
input n_739;
input n_1485;
input n_1028;
input n_1221;
input n_530;
input n_1785;
input n_792;
input n_1262;
input n_580;
input n_1579;
input n_494;
input n_434;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1645;
input n_1124;
input n_1381;
input n_1494;
input n_932;
input n_1183;
input n_1326;
input n_1805;
input n_981;
input n_1110;
input n_1758;
input n_243;
input n_1407;
input n_185;
input n_1204;
input n_1554;
input n_994;
input n_1360;
input n_973;
input n_268;
input n_972;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1564;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_1679;
input n_1858;
input n_353;
input n_1678;
input n_1482;
input n_1361;
input n_1601;
input n_1057;
input n_191;
input n_1834;
input n_978;
input n_1011;
input n_1520;
input n_1509;
input n_828;
input n_322;
input n_1411;
input n_1359;
input n_558;
input n_1721;
input n_116;
input n_39;
input n_653;
input n_1445;
input n_1317;
input n_783;
input n_556;
input n_1127;
input n_170;
input n_1536;
input n_1471;
input n_160;
input n_119;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_987;
input n_936;
input n_1620;
input n_1385;
input n_1525;
input n_541;
input n_499;
input n_1775;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_341;
input n_1270;
input n_109;
input n_1167;
input n_1272;
input n_549;
input n_591;
input n_969;
input n_919;
input n_1663;
input n_50;
input n_1625;
input n_318;
input n_1458;
input n_103;
input n_244;
input n_679;
input n_1630;
input n_220;
input n_663;
input n_1720;
input n_443;
input n_1412;
input n_1738;
input n_1550;
input n_528;
input n_1358;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_1735;
input n_1788;
input n_391;
input n_940;
input n_1537;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_765;
input n_1809;
input n_1843;
input n_122;
input n_1268;
input n_385;
input n_917;
input n_1271;
input n_372;
input n_15;
input n_1530;
input n_631;
input n_399;
input n_1170;
input n_1261;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1323;
input n_1462;
input n_1064;
input n_633;
input n_900;
input n_1446;
input n_1282;
input n_1701;
input n_1093;
input n_1551;
input n_1755;
input n_1285;
input n_193;
input n_733;
input n_761;
input n_731;
input n_336;
input n_1813;
input n_315;
input n_311;
input n_1452;
input n_1573;
input n_8;
input n_668;
input n_758;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_1322;
input n_1473;
input n_835;
input n_446;
input n_1076;
input n_1348;
input n_753;
input n_1770;
input n_701;
input n_1003;
input n_1125;
input n_1710;
input n_1865;
input n_309;
input n_1344;
input n_115;
input n_1390;
input n_401;
input n_485;
input n_1792;
input n_504;
input n_483;
input n_435;
input n_1141;
input n_1629;
input n_291;
input n_1640;
input n_822;
input n_1094;
input n_840;
input n_1459;
input n_1510;
input n_1099;
input n_839;
input n_79;
input n_1754;
input n_3;
input n_759;
input n_567;
input n_91;
input n_240;
input n_369;
input n_1727;
input n_44;
input n_1575;
input n_1848;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_1619;
input n_188;
input n_323;
input n_550;
input n_1315;
input n_1660;
input n_997;
input n_635;
input n_694;
input n_1643;
input n_1320;
input n_1113;
input n_248;
input n_1152;
input n_1845;
input n_921;
input n_1615;
input n_1236;
input n_228;
input n_1265;
input n_1576;
input n_1470;
input n_671;
input n_1533;
input n_1806;
input n_1;
input n_1409;
input n_1148;
input n_1588;
input n_1684;
input n_1673;
input n_1334;
input n_654;
input n_1275;
input n_488;
input n_904;
input n_505;
input n_88;
input n_1696;
input n_498;
input n_1875;
input n_1059;
input n_684;
input n_1039;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_392;
input n_1628;
input n_1289;
input n_1831;
input n_1497;
input n_1866;
input n_459;
input n_1136;
input n_1782;
input n_458;
input n_1190;
input n_1600;
input n_1144;
input n_383;
input n_838;
input n_1558;
input n_1316;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_723;
input n_1393;
input n_658;
input n_630;
input n_1369;
input n_53;
input n_362;
input n_310;
input n_1781;
input n_709;
input n_24;
input n_809;
input n_1686;
input n_235;
input n_881;
input n_1019;
input n_1477;
input n_1777;
input n_662;
input n_641;
input n_910;
input n_290;
input n_741;
input n_939;
input n_1410;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_1325;
input n_1742;
input n_708;
input n_308;
input n_1223;
input n_201;
input n_1768;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1273;
input n_1041;
input n_993;
input n_1862;
input n_948;
input n_922;
input n_1004;
input n_1810;
input n_448;
input n_1347;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_1764;
input n_896;
input n_1737;
input n_1479;
input n_1613;
input n_902;
input n_1031;
input n_1723;
input n_1638;
input n_853;
input n_716;
input n_1571;
input n_1698;
input n_196;
input n_1337;
input n_774;
input n_933;
input n_1779;
input n_596;
input n_954;
input n_1168;
input n_1821;
input n_219;
input n_1310;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1591;
input n_1229;
input n_1683;
input n_68;
input n_1732;
input n_415;
input n_63;
input n_1280;
input n_544;
input n_1516;
input n_1186;
input n_1705;
input n_599;
input n_768;
input n_1091;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_83;
input n_389;
input n_1724;
input n_1670;
input n_1707;
input n_1799;
input n_1126;
input n_195;
input n_1846;
input n_938;
input n_1328;
input n_895;
input n_110;
input n_304;
input n_1639;
input n_583;
input n_1302;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_1581;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_1655;
input n_1818;
input n_33;
input n_1146;
input n_1634;
input n_1203;
input n_998;
input n_1699;
input n_1598;
input n_472;
input n_937;
input n_1474;
input n_265;
input n_1583;
input n_1604;
input n_208;
input n_1631;
input n_1702;
input n_156;
input n_174;
input n_275;
input n_100;
input n_1794;
input n_1375;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_1368;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_1725;
input n_496;
input n_1827;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1752;
input n_1313;
input n_1001;
input n_1722;
input n_1115;
input n_1339;
input n_1002;
input n_1644;
input n_105;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_1129;
input n_1252;
input n_250;
input n_1464;
input n_1296;
input n_773;
input n_165;
input n_1010;
input n_882;
input n_1249;
input n_101;
input n_803;
input n_1871;
input n_329;
input n_718;
input n_1434;
input n_340;
input n_1569;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_523;
input n_1662;
input n_457;
input n_1299;
input n_1870;
input n_177;
input n_782;
input n_364;
input n_258;
input n_431;
input n_1861;
input n_1228;
input n_1244;
input n_1796;
input n_411;
input n_484;
input n_849;
input n_22;
input n_1820;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_447;
input n_1421;
input n_1762;
input n_1233;
input n_1808;
input n_1574;
input n_1672;
input n_1635;
input n_1704;
input n_893;
input n_1582;
input n_841;
input n_886;
input n_1069;
input n_359;
input n_1308;
input n_573;
input n_796;
input n_127;
input n_531;
input n_1730;
input n_1374;
input n_1451;
input n_1487;
input n_675;

output n_7517;

wire n_3527;
wire n_2752;
wire n_4474;
wire n_7329;
wire n_4030;
wire n_7029;
wire n_6790;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_6603;
wire n_2679;
wire n_6557;
wire n_5402;
wire n_6581;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_7277;
wire n_2680;
wire n_3264;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_2002;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_7127;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_5302;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_7053;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_5479;
wire n_2646;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6358;
wire n_6293;
wire n_2482;
wire n_7001;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_6524;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_7464;
wire n_4260;
wire n_3348;
wire n_3261;
wire n_7368;
wire n_2807;
wire n_6664;
wire n_7428;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_7373;
wire n_2390;
wire n_6891;
wire n_4500;
wire n_2322;
wire n_2663;
wire n_5481;
wire n_6539;
wire n_4824;
wire n_7467;
wire n_5340;
wire n_3545;
wire n_6797;
wire n_7392;
wire n_4741;
wire n_4143;
wire n_4273;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_5896;
wire n_7338;
wire n_4567;
wire n_5833;
wire n_6249;
wire n_6887;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_7200;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_6808;
wire n_3749;
wire n_5691;
wire n_3482;
wire n_7490;
wire n_6295;
wire n_5403;
wire n_1900;
wire n_6096;
wire n_4268;
wire n_6338;
wire n_6992;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_3325;
wire n_6681;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_6542;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_6452;
wire n_5247;
wire n_5464;
wire n_7306;
wire n_4476;
wire n_6740;
wire n_6978;
wire n_7507;
wire n_2956;
wire n_5210;
wire n_7215;
wire n_2382;
wire n_7379;
wire n_7441;
wire n_5292;
wire n_1918;
wire n_7438;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_3458;
wire n_5843;
wire n_7108;
wire n_3511;
wire n_2077;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_6156;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_7162;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_7331;
wire n_5913;
wire n_4530;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_6872;
wire n_6644;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_6236;
wire n_7104;
wire n_3506;
wire n_4827;
wire n_6801;
wire n_4993;
wire n_7397;
wire n_3678;
wire n_7205;
wire n_2791;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_6563;
wire n_5968;
wire n_3549;
wire n_3914;
wire n_6398;
wire n_5586;
wire n_7461;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_7224;
wire n_6966;
wire n_5056;
wire n_2015;
wire n_7259;
wire n_5984;
wire n_5204;
wire n_6705;
wire n_6724;
wire n_2877;
wire n_7307;
wire n_6776;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_6624;
wire n_6710;
wire n_6883;
wire n_3172;
wire n_4033;
wire n_2659;
wire n_3747;
wire n_6553;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_6261;
wire n_6659;
wire n_7351;
wire n_3614;
wire n_7256;
wire n_2257;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_6893;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_3559;
wire n_5778;
wire n_7021;
wire n_5179;
wire n_2435;
wire n_6337;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_6378;
wire n_5549;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_7488;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_6206;
wire n_2954;
wire n_4438;
wire n_6538;
wire n_3814;
wire n_6996;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_7231;
wire n_4195;
wire n_7007;
wire n_6579;
wire n_5091;
wire n_4866;
wire n_7230;
wire n_2019;
wire n_5708;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_7403;
wire n_6665;
wire n_3147;
wire n_3661;
wire n_7168;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2649;
wire n_6033;
wire n_6461;
wire n_6860;
wire n_2919;
wire n_7322;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_6709;
wire n_2632;
wire n_5557;
wire n_6914;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_7287;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_3087;
wire n_6009;
wire n_7221;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_3704;
wire n_6382;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_6615;
wire n_7294;
wire n_6192;
wire n_5773;
wire n_7414;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_6418;
wire n_6263;
wire n_1943;
wire n_6731;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_7185;
wire n_5149;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_7141;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_6619;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_6759;
wire n_6903;
wire n_3466;
wire n_7416;
wire n_2074;
wire n_5031;
wire n_6768;
wire n_7092;
wire n_7233;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_7191;
wire n_2117;
wire n_6189;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_6761;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_7202;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_7445;
wire n_5858;
wire n_5985;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_6366;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_7176;
wire n_5552;
wire n_6074;
wire n_3764;
wire n_4773;
wire n_5028;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_2125;
wire n_4974;
wire n_5123;
wire n_6689;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_4856;
wire n_2618;
wire n_7096;
wire n_4216;
wire n_2707;
wire n_5596;
wire n_6482;
wire n_2849;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_6335;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_3713;
wire n_6229;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_7293;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_7144;
wire n_3931;
wire n_2190;
wire n_2516;
wire n_4991;
wire n_7316;
wire n_7508;
wire n_3070;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_6943;
wire n_1957;
wire n_1953;
wire n_6631;
wire n_5889;
wire n_7151;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_6728;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_7472;
wire n_4800;
wire n_7075;
wire n_5427;
wire n_4440;
wire n_4425;
wire n_6770;
wire n_5450;
wire n_6508;
wire n_2821;
wire n_3696;
wire n_4781;
wire n_6031;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_7105;
wire n_7013;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_7254;
wire n_2448;
wire n_2211;
wire n_5904;
wire n_6628;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_6456;
wire n_7407;
wire n_3277;
wire n_4863;
wire n_5463;
wire n_2978;
wire n_6328;
wire n_6929;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_2958;
wire n_7481;
wire n_4429;
wire n_6484;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_7182;
wire n_5476;
wire n_5483;
wire n_5511;
wire n_3486;
wire n_6639;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_7423;
wire n_3256;
wire n_7375;
wire n_7076;
wire n_6344;
wire n_6435;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_7419;
wire n_6600;
wire n_7010;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_5073;
wire n_6555;
wire n_4306;
wire n_6360;
wire n_6735;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_6803;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_5419;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_6036;
wire n_7346;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_6650;
wire n_6573;
wire n_6904;
wire n_3753;
wire n_6329;
wire n_7385;
wire n_6244;
wire n_4846;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_7295;
wire n_4076;
wire n_7148;
wire n_3142;
wire n_7169;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_6756;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_6946;
wire n_5931;
wire n_4635;
wire n_5532;
wire n_7311;
wire n_3740;
wire n_6804;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_7039;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_6427;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6442;
wire n_6188;
wire n_3421;
wire n_3548;
wire n_4906;
wire n_6846;
wire n_4630;
wire n_6840;
wire n_6645;
wire n_4829;
wire n_6749;
wire n_6915;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_7455;
wire n_6247;
wire n_5921;
wire n_4966;
wire n_2250;
wire n_6104;
wire n_3321;
wire n_4188;
wire n_2001;
wire n_7509;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_3715;
wire n_2610;
wire n_2626;
wire n_7497;
wire n_7315;
wire n_2892;
wire n_6939;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_6706;
wire n_7431;
wire n_3842;
wire n_4202;
wire n_6909;
wire n_2044;
wire n_5679;
wire n_6487;
wire n_3886;
wire n_2619;
wire n_5141;
wire n_3098;
wire n_6627;
wire n_4503;
wire n_7253;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_2968;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_7452;
wire n_6551;
wire n_3386;
wire n_7505;
wire n_3921;
wire n_2177;
wire n_6516;
wire n_2766;
wire n_4196;
wire n_7318;
wire n_2613;
wire n_7411;
wire n_7326;
wire n_5667;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_6500;
wire n_5027;
wire n_2343;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_1921;
wire n_6630;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_6798;
wire n_5999;
wire n_2110;
wire n_7498;
wire n_6421;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_4355;
wire n_7453;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_6652;
wire n_7183;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_6395;
wire n_3497;
wire n_6403;
wire n_4542;
wire n_5451;
wire n_6578;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_6350;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_2068;
wire n_3595;
wire n_6875;
wire n_7189;
wire n_4060;
wire n_6194;
wire n_2459;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_6475;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1940;
wire n_3683;
wire n_6502;
wire n_6944;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_6805;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_7240;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_7499;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_6075;
wire n_6559;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_6248;
wire n_6541;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_4733;
wire n_7219;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_6638;
wire n_7063;
wire n_7402;
wire n_6351;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_7382;
wire n_4004;
wire n_5238;
wire n_3630;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_6474;
wire n_5743;
wire n_6481;
wire n_1956;
wire n_4111;
wire n_5633;
wire n_7510;
wire n_3786;
wire n_6022;
wire n_6991;
wire n_2828;
wire n_7434;
wire n_5950;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_6744;
wire n_3645;
wire n_5705;
wire n_6927;
wire n_7335;
wire n_4996;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_7495;
wire n_4785;
wire n_2870;
wire n_1893;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_3610;
wire n_2443;
wire n_5011;
wire n_6757;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_6485;
wire n_5848;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6495;
wire n_6209;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_7413;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_4628;
wire n_6802;
wire n_7343;
wire n_5982;
wire n_7109;
wire n_4083;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_7506;
wire n_3940;
wire n_6809;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_6349;
wire n_3680;
wire n_6716;
wire n_3565;
wire n_6905;
wire n_5388;
wire n_7470;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_6203;
wire n_2138;
wire n_6407;
wire n_3040;
wire n_4230;
wire n_6899;
wire n_6413;
wire n_3360;
wire n_1930;
wire n_3585;
wire n_7070;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_7299;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_6960;
wire n_4073;
wire n_7249;
wire n_5763;
wire n_3633;
wire n_6061;
wire n_2584;
wire n_4001;
wire n_5701;
wire n_7002;
wire n_6273;
wire n_7094;
wire n_7396;
wire n_3111;
wire n_2997;
wire n_7018;
wire n_6746;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_6545;
wire n_6763;
wire n_1996;
wire n_2009;
wire n_5907;
wire n_4339;
wire n_7297;
wire n_6013;
wire n_6182;
wire n_6754;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_5895;
wire n_2651;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_3632;
wire n_2522;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_3457;
wire n_5384;
wire n_6477;
wire n_7486;
wire n_2324;
wire n_6575;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_6391;
wire n_2740;
wire n_1991;
wire n_7140;
wire n_4066;
wire n_6252;
wire n_6426;
wire n_4681;
wire n_3303;
wire n_6592;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_3768;
wire n_4295;
wire n_4100;
wire n_6668;
wire n_2372;
wire n_3445;
wire n_2105;
wire n_4087;
wire n_4473;
wire n_4619;
wire n_6670;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_6962;
wire n_2429;
wire n_6779;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_6901;
wire n_4266;
wire n_6336;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_6503;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_7100;
wire n_4777;
wire n_7243;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_7415;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_3366;
wire n_6998;
wire n_7395;
wire n_5844;
wire n_6298;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_6609;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_4976;
wire n_6525;
wire n_3555;
wire n_5938;
wire n_7274;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_6494;
wire n_3556;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_2148;
wire n_5548;
wire n_6974;
wire n_4663;
wire n_5840;
wire n_6882;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_6498;
wire n_6562;
wire n_3293;
wire n_4902;
wire n_4686;
wire n_2384;
wire n_3707;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_6965;
wire n_2058;
wire n_3231;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_6963;
wire n_6951;
wire n_3058;
wire n_5355;
wire n_2047;
wire n_3398;
wire n_3709;
wire n_6284;
wire n_3592;
wire n_5321;
wire n_7454;
wire n_2536;
wire n_3399;
wire n_4772;
wire n_6931;
wire n_6521;
wire n_5915;
wire n_7276;
wire n_6379;
wire n_7085;
wire n_6306;
wire n_4120;
wire n_6834;
wire n_2880;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_5116;
wire n_3771;
wire n_7225;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_6471;
wire n_6949;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_6760;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_6589;
wire n_3083;
wire n_4570;
wire n_7014;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_5059;
wire n_4655;
wire n_7459;
wire n_7160;
wire n_7324;
wire n_6046;
wire n_7054;
wire n_4493;
wire n_6055;
wire n_7161;
wire n_6364;
wire n_6091;
wire n_6348;
wire n_4896;
wire n_4851;
wire n_6848;
wire n_2479;
wire n_6788;
wire n_6144;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_6896;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_4901;
wire n_3480;
wire n_7201;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_7241;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_4602;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_2537;
wire n_3745;
wire n_6748;
wire n_7430;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_5901;
wire n_2837;
wire n_2446;
wire n_6582;
wire n_4116;
wire n_5360;
wire n_7269;
wire n_7047;
wire n_2671;
wire n_2702;
wire n_6937;
wire n_4363;
wire n_3561;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_3154;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_7067;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_6607;
wire n_4439;
wire n_4985;
wire n_3382;
wire n_7117;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_4660;
wire n_3081;
wire n_6446;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_2579;
wire n_1961;
wire n_6849;
wire n_2960;
wire n_3270;
wire n_6807;
wire n_2844;
wire n_1979;
wire n_6616;
wire n_6719;
wire n_4814;
wire n_6178;
wire n_6677;
wire n_2221;
wire n_5502;
wire n_2317;
wire n_2838;
wire n_2200;
wire n_7302;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_7238;
wire n_6862;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_7292;
wire n_5098;
wire n_6000;
wire n_6774;
wire n_6443;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_7248;
wire n_3830;
wire n_3252;
wire n_6647;
wire n_5466;
wire n_6941;
wire n_7239;
wire n_6552;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_7112;
wire n_3420;
wire n_3859;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_4831;
wire n_4782;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_2162;
wire n_5953;
wire n_5703;
wire n_6886;
wire n_7078;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_7006;
wire n_4031;
wire n_5119;
wire n_4147;
wire n_3073;
wire n_6531;
wire n_3571;
wire n_4576;
wire n_7354;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_6726;
wire n_6983;
wire n_7513;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_6935;
wire n_2899;
wire n_6984;
wire n_6778;
wire n_6897;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_6345;
wire n_6386;
wire n_3728;
wire n_2722;
wire n_6596;
wire n_5107;
wire n_7165;
wire n_4680;
wire n_5067;
wire n_6830;
wire n_2061;
wire n_2685;
wire n_5987;
wire n_2512;
wire n_2788;
wire n_6642;
wire n_6291;
wire n_6510;
wire n_5264;
wire n_2595;
wire n_3084;
wire n_6781;
wire n_4593;
wire n_7123;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_6509;
wire n_2717;
wire n_6376;
wire n_2981;
wire n_4995;
wire n_5873;
wire n_6514;
wire n_4498;
wire n_6741;
wire n_6434;
wire n_5741;
wire n_2743;
wire n_2969;
wire n_3429;
wire n_2466;
wire n_6593;
wire n_3758;
wire n_6690;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_6947;
wire n_4850;
wire n_3716;
wire n_7157;
wire n_2926;
wire n_4937;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_6375;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_7091;
wire n_4354;
wire n_6429;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_2855;
wire n_2848;
wire n_6775;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_6970;
wire n_6948;
wire n_3460;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_6920;
wire n_2693;
wire n_7409;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_7381;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_7087;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_2365;
wire n_5684;
wire n_7228;
wire n_5981;
wire n_6632;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_6623;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_2224;
wire n_6933;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_3046;
wire n_2293;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_6908;
wire n_5097;
wire n_2695;
wire n_7084;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_6537;
wire n_4003;
wire n_6390;
wire n_2302;
wire n_6799;
wire n_3014;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_7195;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_7298;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_7115;
wire n_2495;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_6412;
wire n_6271;
wire n_7235;
wire n_2511;
wire n_6572;
wire n_3981;
wire n_7271;
wire n_2681;
wire n_7222;
wire n_2535;
wire n_3031;
wire n_6930;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_3138;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_6584;
wire n_4494;
wire n_6387;
wire n_4201;
wire n_6470;
wire n_7206;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_6625;
wire n_4074;
wire n_7383;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_6826;
wire n_2662;
wire n_4386;
wire n_6341;
wire n_6374;
wire n_3917;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_2296;
wire n_5735;
wire n_6363;
wire n_6588;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_6811;
wire n_6687;
wire n_4658;
wire n_7135;
wire n_6037;
wire n_4186;
wire n_2241;
wire n_6865;
wire n_7211;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_7132;
wire n_3377;
wire n_6722;
wire n_6420;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_6911;
wire n_7129;
wire n_7080;
wire n_3374;
wire n_4870;
wire n_6981;
wire n_4818;
wire n_7436;
wire n_7020;
wire n_5935;
wire n_6696;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_6653;
wire n_6372;
wire n_4129;
wire n_7120;
wire n_5488;
wire n_6900;
wire n_5727;
wire n_3599;
wire n_6660;
wire n_5988;
wire n_6424;
wire n_5646;
wire n_7448;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_6787;
wire n_5832;
wire n_6254;
wire n_7460;
wire n_3401;
wire n_7142;
wire n_6423;
wire n_6526;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_7465;
wire n_5470;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_6222;
wire n_2218;
wire n_2593;
wire n_6969;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_6587;
wire n_6688;
wire n_6505;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_6762;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_6987;
wire n_3995;
wire n_3908;
wire n_6453;
wire n_6308;
wire n_3892;
wire n_7449;
wire n_3501;
wire n_3216;
wire n_3568;
wire n_2555;
wire n_2708;
wire n_6187;
wire n_6597;
wire n_4844;
wire n_6220;
wire n_4049;
wire n_2661;
wire n_7479;
wire n_2470;
wire n_3551;
wire n_5037;
wire n_7305;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_6439;
wire n_4324;
wire n_1898;
wire n_1907;
wire n_6547;
wire n_7177;
wire n_5160;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_5484;
wire n_1895;
wire n_7353;
wire n_4104;
wire n_3791;
wire n_6478;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_7050;
wire n_3151;
wire n_6906;
wire n_3016;
wire n_2460;
wire n_6739;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_5385;
wire n_7482;
wire n_3990;
wire n_5622;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_3735;
wire n_7410;
wire n_6422;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_6604;
wire n_3964;
wire n_6611;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_6999;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_6440;
wire n_4977;
wire n_2492;
wire n_6976;
wire n_7234;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_2900;
wire n_2912;
wire n_5936;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_6784;
wire n_1950;
wire n_2264;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_2928;
wire n_5505;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_5504;
wire n_7348;
wire n_4118;
wire n_6829;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_2730;
wire n_6464;
wire n_5129;
wire n_7320;
wire n_4704;
wire n_2720;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_6838;
wire n_2700;
wire n_6368;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_7155;
wire n_6640;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_6850;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_2454;
wire n_6550;
wire n_6656;
wire n_6972;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_7043;
wire n_3317;
wire n_7266;
wire n_5653;
wire n_4835;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_4790;
wire n_7035;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_7442;
wire n_4727;
wire n_6568;
wire n_3654;
wire n_5627;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_7153;
wire n_6258;
wire n_2173;
wire n_3982;
wire n_7350;
wire n_3647;
wire n_7314;
wire n_6026;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_6700;
wire n_7136;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_5697;
wire n_2020;
wire n_5606;
wire n_6727;
wire n_2310;
wire n_5911;
wire n_7340;
wire n_3600;
wire n_7303;
wire n_6139;
wire n_7399;
wire n_5382;
wire n_4327;
wire n_7387;
wire n_3190;
wire n_3027;
wire n_6454;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_3967;
wire n_6333;
wire n_7004;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_3096;
wire n_7207;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_7167;
wire n_2234;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_5841;
wire n_7146;
wire n_7030;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_3344;
wire n_4754;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_3117;
wire n_4684;
wire n_3384;
wire n_5279;
wire n_7159;
wire n_2592;
wire n_3490;
wire n_7280;
wire n_5043;
wire n_7339;
wire n_4241;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_6455;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_6476;
wire n_5232;
wire n_4256;
wire n_2560;
wire n_5035;
wire n_3037;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_2007;
wire n_3363;
wire n_6636;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_6554;
wire n_5631;
wire n_3481;
wire n_6994;
wire n_7401;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_7321;
wire n_4457;
wire n_2150;
wire n_6785;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_6870;
wire n_3305;
wire n_6643;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_6695;
wire n_3354;
wire n_5608;
wire n_6501;
wire n_2204;
wire n_2040;
wire n_6466;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_6467;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_7188;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_4217;
wire n_5277;
wire n_6507;
wire n_1942;
wire n_6618;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_3969;
wire n_6873;
wire n_2282;
wire n_4605;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_7101;
wire n_2428;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_7261;
wire n_4592;
wire n_4999;
wire n_6993;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_2589;
wire n_4086;
wire n_6767;
wire n_4656;
wire n_4862;
wire n_5687;
wire n_6558;
wire n_6755;
wire n_6153;
wire n_3536;
wire n_7263;
wire n_3782;
wire n_6608;
wire n_6202;
wire n_6780;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_6635;
wire n_7245;
wire n_7310;
wire n_6359;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_7093;
wire n_4177;
wire n_2501;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_7418;
wire n_6353;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_6577;
wire n_2028;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_7312;
wire n_7514;
wire n_6105;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_7113;
wire n_6548;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_6657;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_2676;
wire n_7282;
wire n_4550;
wire n_2770;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_3278;
wire n_2375;
wire n_5579;
wire n_4167;
wire n_6380;
wire n_3608;
wire n_4895;
wire n_6163;
wire n_7170;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_5188;
wire n_6674;
wire n_5049;
wire n_2212;
wire n_7489;
wire n_6331;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_6493;
wire n_7363;
wire n_7281;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_2358;
wire n_3546;
wire n_2355;
wire n_5887;
wire n_3068;
wire n_6321;
wire n_5683;
wire n_3002;
wire n_7192;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_2351;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_6824;
wire n_6954;
wire n_6450;
wire n_6995;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_6347;
wire n_6496;
wire n_4776;
wire n_2704;
wire n_6745;
wire n_3729;
wire n_6698;
wire n_4471;
wire n_6968;
wire n_7377;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_7296;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_6743;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_6330;
wire n_7178;
wire n_1941;
wire n_7045;
wire n_3637;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_6015;
wire n_6408;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_7300;
wire n_2297;
wire n_6861;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_6528;
wire n_3820;
wire n_5144;
wire n_6895;
wire n_3072;
wire n_2961;
wire n_5509;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_7400;
wire n_3631;
wire n_7393;
wire n_6590;
wire n_6523;
wire n_5169;
wire n_4885;
wire n_7475;
wire n_4698;
wire n_3674;
wire n_5349;
wire n_6472;
wire n_3763;
wire n_6389;
wire n_3499;
wire n_5534;
wire n_3947;
wire n_3910;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_2678;
wire n_6869;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_3088;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_2421;
wire n_3295;
wire n_5751;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_6885;
wire n_5039;
wire n_6580;
wire n_6613;
wire n_4265;
wire n_6404;
wire n_6120;
wire n_3557;
wire n_2269;
wire n_7491;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_7150;
wire n_6530;
wire n_6602;
wire n_4149;
wire n_4958;
wire n_6135;
wire n_5563;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_2239;
wire n_6942;
wire n_6892;
wire n_4730;
wire n_7357;
wire n_6782;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_2304;
wire n_2514;
wire n_6977;
wire n_7229;
wire n_7336;
wire n_5932;
wire n_6598;
wire n_6795;
wire n_6121;
wire n_3430;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_6614;
wire n_6506;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_7493;
wire n_5664;
wire n_2738;
wire n_6406;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_3041;
wire n_2797;
wire n_5823;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_6989;
wire n_6299;
wire n_7424;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_7273;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_4834;
wire n_5332;
wire n_7149;
wire n_2866;
wire n_7116;
wire n_3153;
wire n_2346;
wire n_4692;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_6758;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_6629;
wire n_5288;
wire n_2694;
wire n_6356;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_7033;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_7147;
wire n_5294;
wire n_5570;
wire n_6411;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4802;
wire n_4793;
wire n_6032;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_6918;
wire n_4674;
wire n_4796;
wire n_7138;
wire n_6401;
wire n_7279;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_7137;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_7474;
wire n_4589;
wire n_7124;
wire n_5978;
wire n_6853;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_4625;
wire n_7098;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_5575;
wire n_6654;
wire n_4968;
wire n_6907;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_2109;
wire n_2709;
wire n_3419;
wire n_7323;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_6517;
wire n_4892;
wire n_6339;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_7247;
wire n_6394;
wire n_5607;
wire n_2782;
wire n_3929;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_6504;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_6814;
wire n_7216;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_6691;
wire n_3948;
wire n_4839;
wire n_5969;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6343;
wire n_6005;
wire n_2060;
wire n_3883;
wire n_6686;
wire n_4032;
wire n_2571;
wire n_6437;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_6536;
wire n_6684;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_6697;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_5140;
wire n_2942;
wire n_6062;
wire n_4541;
wire n_6715;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_6771;
wire n_4171;
wire n_5847;
wire n_7204;
wire n_7022;
wire n_6383;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_6877;
wire n_7308;
wire n_7476;
wire n_4884;
wire n_3580;
wire n_4276;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_5718;
wire n_7208;
wire n_5001;
wire n_6567;
wire n_5658;
wire n_4174;
wire n_6868;
wire n_7290;
wire n_5131;
wire n_6813;
wire n_5546;
wire n_6294;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_6520;
wire n_3119;
wire n_6671;
wire n_4740;
wire n_4394;
wire n_5544;
wire n_6444;
wire n_6637;
wire n_6729;
wire n_5660;
wire n_6958;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_2810;
wire n_6703;
wire n_1884;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_7265;
wire n_4180;
wire n_4459;
wire n_6878;
wire n_3624;
wire n_6725;
wire n_5808;
wire n_6527;
wire n_4594;
wire n_7289;
wire n_2748;
wire n_4642;
wire n_6913;
wire n_7473;
wire n_7242;
wire n_6533;
wire n_7164;
wire n_2925;
wire n_3544;
wire n_6845;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_7483;
wire n_5710;
wire n_2628;
wire n_7389;
wire n_3219;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_7046;
wire n_4587;
wire n_3688;
wire n_5008;
wire n_3871;
wire n_3757;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_6357;
wire n_3479;
wire n_5499;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_6522;
wire n_4285;
wire n_7097;
wire n_7000;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_2755;
wire n_5109;
wire n_6713;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_2220;
wire n_7342;
wire n_7044;
wire n_6108;
wire n_6100;
wire n_6800;
wire n_7364;
wire n_6866;
wire n_7114;
wire n_6373;
wire n_4433;
wire n_2829;
wire n_7332;
wire n_5862;
wire n_7477;
wire n_1914;
wire n_2253;
wire n_7468;
wire n_5886;
wire n_6415;
wire n_6783;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_6340;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_6392;
wire n_6513;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_6720;
wire n_5883;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_5630;
wire n_6666;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_2113;
wire n_6815;
wire n_6207;
wire n_6381;
wire n_3711;
wire n_5054;
wire n_6571;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_2812;
wire n_3300;
wire n_7061;
wire n_7066;
wire n_5496;
wire n_7485;
wire n_3104;
wire n_7174;
wire n_4122;
wire n_6661;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_6967;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_5132;
wire n_3498;
wire n_2350;
wire n_6414;
wire n_5535;
wire n_4506;
wire n_6097;
wire n_6057;
wire n_6936;
wire n_4728;
wire n_7171;
wire n_1886;
wire n_4346;
wire n_7003;
wire n_2187;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_6922;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_7501;
wire n_6432;
wire n_2055;
wire n_2998;
wire n_7366;
wire n_4359;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_6880;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_6926;
wire n_3057;
wire n_5761;
wire n_6699;
wire n_3983;
wire n_3318;
wire n_7232;
wire n_3385;
wire n_7511;
wire n_3773;
wire n_3494;
wire n_6957;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_6694;
wire n_3260;
wire n_2496;
wire n_3349;
wire n_6449;
wire n_4348;
wire n_7422;
wire n_3139;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_3636;
wire n_6591;
wire n_7466;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_6594;
wire n_6342;
wire n_6195;
wire n_2716;
wire n_6441;
wire n_7158;
wire n_2944;
wire n_3439;
wire n_2780;
wire n_7500;
wire n_4084;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_6354;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_6662;
wire n_7494;
wire n_3984;
wire n_4389;
wire n_6433;
wire n_6200;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_2660;
wire n_3426;
wire n_6902;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_7197;
wire n_3737;
wire n_6369;
wire n_5657;
wire n_3579;
wire n_2379;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_6956;
wire n_2284;
wire n_6451;
wire n_3005;
wire n_5420;
wire n_6497;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_4387;
wire n_3186;
wire n_2508;
wire n_6701;
wire n_2594;
wire n_5298;
wire n_3417;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_7032;
wire n_3392;
wire n_7198;
wire n_6884;
wire n_5081;
wire n_6921;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_6876;
wire n_3512;
wire n_4552;
wire n_7193;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_5957;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_6362;
wire n_4328;
wire n_5191;
wire n_6067;
wire n_2893;
wire n_6833;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_2280;
wire n_7126;
wire n_5867;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_7496;
wire n_6430;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_7196;
wire n_2614;
wire n_7360;
wire n_5428;
wire n_6325;
wire n_2494;
wire n_4865;
wire n_6678;
wire n_2128;
wire n_4071;
wire n_6564;
wire n_7268;
wire n_4436;
wire n_5786;
wire n_5822;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_6385;
wire n_5798;
wire n_4137;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_4535;
wire n_4385;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_7073;
wire n_6309;
wire n_3732;
wire n_6519;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_7349;
wire n_1929;
wire n_4319;
wire n_6585;
wire n_2929;
wire n_4358;
wire n_7122;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_6490;
wire n_4651;
wire n_3167;
wire n_4748;
wire n_2857;
wire n_4618;
wire n_6721;
wire n_3787;
wire n_4025;
wire n_3050;
wire n_3919;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_7019;
wire n_5315;
wire n_3708;
wire n_2633;
wire n_5752;
wire n_2907;
wire n_2353;
wire n_2528;
wire n_5746;
wire n_4910;
wire n_2325;
wire n_4724;
wire n_3718;
wire n_6685;
wire n_3390;
wire n_2298;
wire n_4666;
wire n_3140;
wire n_4082;
wire n_2320;
wire n_3976;
wire n_3381;
wire n_2546;
wire n_2813;
wire n_7347;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_6971;
wire n_3336;
wire n_5903;
wire n_7199;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_6549;
wire n_5003;
wire n_3840;
wire n_6540;
wire n_7166;
wire n_2198;
wire n_6658;
wire n_5369;
wire n_6683;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_6327;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_7213;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_6820;
wire n_2497;
wire n_5446;
wire n_7107;
wire n_4561;
wire n_3291;
wire n_7456;
wire n_7369;
wire n_2578;
wire n_2475;
wire n_7250;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_6676;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_5024;
wire n_7012;
wire n_3043;
wire n_2747;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_4412;
wire n_2845;
wire n_2036;
wire n_6923;
wire n_3358;
wire n_6704;
wire n_2003;
wire n_2533;
wire n_7406;
wire n_4682;
wire n_6673;
wire n_2419;
wire n_2330;
wire n_6534;
wire n_5078;
wire n_4810;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_6246;
wire n_5005;
wire n_6126;
wire n_7372;
wire n_7427;
wire n_6151;
wire n_6828;
wire n_6841;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_5474;
wire n_2767;
wire n_7009;
wire n_3376;
wire n_7371;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_7463;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_6889;
wire n_2749;
wire n_5962;
wire n_4413;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_6723;
wire n_7398;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_7011;
wire n_3405;
wire n_2313;
wire n_6393;
wire n_7074;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_3131;
wire n_4138;
wire n_7083;
wire n_1973;
wire n_2882;
wire n_7143;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_4577;
wire n_6312;
wire n_2154;
wire n_1986;
wire n_6711;
wire n_2624;
wire n_6818;
wire n_6438;
wire n_2054;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_2938;
wire n_7209;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_7330;
wire n_6007;
wire n_6734;
wire n_6535;
wire n_6879;
wire n_3106;
wire n_6208;
wire n_7190;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_4620;
wire n_5397;
wire n_6457;
wire n_6255;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_5566;
wire n_3304;
wire n_7288;
wire n_4388;
wire n_7362;
wire n_7082;
wire n_7237;
wire n_3247;
wire n_7131;
wire n_6276;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_7042;
wire n_2809;
wire n_5652;
wire n_5805;
wire n_7304;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_6934;
wire n_7386;
wire n_2972;
wire n_7391;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_7023;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_7404;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_6765;
wire n_4973;
wire n_4792;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_2534;
wire n_6352;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_6093;
wire n_5370;
wire n_7378;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_5902;
wire n_2510;
wire n_6402;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_6764;
wire n_2639;
wire n_7016;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_6215;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_6955;
wire n_5952;
wire n_7180;
wire n_2086;
wire n_1926;
wire n_6569;
wire n_2966;
wire n_2409;
wire n_3431;
wire n_3355;
wire n_7031;
wire n_5716;
wire n_3897;
wire n_7103;
wire n_6605;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2597;
wire n_2321;
wire n_6832;
wire n_5980;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_6544;
wire n_6469;
wire n_5036;
wire n_6332;
wire n_2186;
wire n_5790;
wire n_7130;
wire n_6680;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_7134;
wire n_3042;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_5485;
wire n_5525;
wire n_7102;
wire n_6259;
wire n_3004;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_7133;
wire n_3838;
wire n_6289;
wire n_6651;
wire n_4059;
wire n_6565;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_7227;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_6836;
wire n_3273;
wire n_2918;
wire n_6595;
wire n_6186;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_7236;
wire n_4833;
wire n_3394;
wire n_6405;
wire n_2235;
wire n_5850;
wire n_6786;
wire n_4564;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_6769;
wire n_6844;
wire n_4322;
wire n_6361;
wire n_2260;
wire n_4080;
wire n_2206;
wire n_6766;
wire n_4185;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_6751;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_7457;
wire n_5372;
wire n_6736;
wire n_4507;
wire n_4756;
wire n_5860;
wire n_2422;
wire n_6416;
wire n_2933;
wire n_7515;
wire n_3387;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_7049;
wire n_6945;
wire n_6143;
wire n_2736;
wire n_6491;
wire n_3825;
wire n_4198;
wire n_7172;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_2664;
wire n_4154;
wire n_7344;
wire n_5859;
wire n_6447;
wire n_4390;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_7325;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_6175;
wire n_6445;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_6499;
wire n_1982;
wire n_5311;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_6842;
wire n_4002;
wire n_7361;
wire n_4679;
wire n_6397;
wire n_3815;
wire n_6827;
wire n_2193;
wire n_2369;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_3504;
wire n_2587;
wire n_5547;
wire n_4693;
wire n_6822;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_7079;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_7309;
wire n_7119;
wire n_3026;
wire n_7184;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_3112;
wire n_2562;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_5301;
wire n_5126;
wire n_6732;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_6817;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_3779;
wire n_6982;
wire n_7291;
wire n_2275;
wire n_7435;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_1891;
wire n_6560;
wire n_6634;
wire n_5348;
wire n_4868;
wire n_7017;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_5654;
wire n_2318;
wire n_2819;
wire n_2229;
wire n_6400;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_3045;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_6655;
wire n_1905;
wire n_5448;
wire n_2573;
wire n_6480;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_3249;
wire n_3483;
wire n_6621;
wire n_6851;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_7420;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_3033;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_2089;
wire n_6283;
wire n_4688;
wire n_7156;
wire n_4939;
wire n_5900;
wire n_7319;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_6819;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_6898;
wire n_6570;
wire n_5486;
wire n_2135;
wire n_7260;
wire n_6894;
wire n_4475;
wire n_6843;
wire n_5432;
wire n_5851;
wire n_7516;
wire n_6317;
wire n_6928;
wire n_6707;
wire n_7244;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_6806;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_6835;
wire n_7286;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_2461;
wire n_3719;
wire n_7154;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_5295;
wire n_6088;
wire n_1999;
wire n_7194;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_5855;
wire n_7175;
wire n_3965;
wire n_3905;
wire n_7163;
wire n_3797;
wire n_7027;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_6964;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_7068;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_2323;
wire n_4549;
wire n_7327;
wire n_6610;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6752;
wire n_6959;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_7317;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_6675;
wire n_2832;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_7384;
wire n_2914;
wire n_5656;
wire n_7218;
wire n_1988;
wire n_5678;
wire n_6561;
wire n_6858;
wire n_5865;
wire n_6050;
wire n_7512;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_4809;
wire n_7152;
wire n_4012;
wire n_2049;
wire n_5212;
wire n_4760;
wire n_6823;
wire n_3606;
wire n_7062;
wire n_7090;
wire n_2232;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_7223;
wire n_5251;
wire n_5965;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_6796;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_5042;
wire n_7055;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_5368;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_3183;
wire n_3607;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_7388;
wire n_7056;
wire n_7437;
wire n_6489;
wire n_5310;
wire n_2769;
wire n_4987;
wire n_6714;
wire n_3013;
wire n_4572;
wire n_7417;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_7446;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_6620;
wire n_6791;
wire n_4540;
wire n_6821;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_6583;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_3089;
wire n_4854;
wire n_5477;
wire n_2727;
wire n_5234;
wire n_6890;
wire n_6988;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_7257;
wire n_3126;
wire n_2759;
wire n_6973;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_6488;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_7005;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_7081;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_6399;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_3095;
wire n_7341;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_4775;
wire n_6256;
wire n_2620;
wire n_7264;
wire n_2499;
wire n_2549;
wire n_6648;
wire n_7492;
wire n_6649;
wire n_3093;
wire n_2970;
wire n_6910;
wire n_3885;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_6431;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_7285;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_6512;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_7051;
wire n_6773;
wire n_2155;
wire n_6231;
wire n_7503;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_5659;
wire n_6859;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_5598;
wire n_2753;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_6912;
wire n_3567;
wire n_7425;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_5783;
wire n_6837;
wire n_6747;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_6916;
wire n_2378;
wire n_5530;
wire n_6718;
wire n_5809;
wire n_2213;
wire n_7121;
wire n_6410;
wire n_6473;
wire n_4056;
wire n_4806;
wire n_5993;
wire n_4015;
wire n_6574;
wire n_2924;
wire n_6492;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_3170;
wire n_2311;
wire n_6857;
wire n_2287;
wire n_3415;
wire n_6975;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_6646;
wire n_4234;
wire n_3467;
wire n_5821;
wire n_3179;
wire n_6622;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_7469;
wire n_3699;
wire n_6118;
wire n_2120;
wire n_7125;
wire n_6028;
wire n_6663;
wire n_6532;
wire n_3816;
wire n_3528;
wire n_6267;
wire n_6682;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_7203;
wire n_5943;
wire n_6556;
wire n_4880;
wire n_4051;
wire n_2834;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_7128;
wire n_5335;
wire n_6365;
wire n_7111;
wire n_2801;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_3623;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_6950;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_7284;
wire n_3615;
wire n_7057;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_7064;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_7278;
wire n_6772;
wire n_7088;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_7048;
wire n_6617;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_3471;
wire n_4075;
wire n_2932;
wire n_2027;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_6777;
wire n_6742;
wire n_7447;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_6479;
wire n_5099;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_7365;
wire n_3443;
wire n_3988;
wire n_2599;
wire n_5022;
wire n_6370;
wire n_2075;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_7275;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_6856;
wire n_3009;
wire n_7095;
wire n_7390;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_7037;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_6693;
wire n_6712;
wire n_3957;
wire n_3418;
wire n_7471;
wire n_6465;
wire n_5673;
wire n_5814;
wire n_6586;
wire n_7058;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_6730;
wire n_6367;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_6515;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_7429;
wire n_6940;
wire n_2949;
wire n_7008;
wire n_6468;
wire n_4269;
wire n_1927;
wire n_7139;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_7432;
wire n_2124;
wire n_1894;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_6483;
wire n_4463;
wire n_5357;
wire n_7173;
wire n_3648;
wire n_6576;
wire n_6810;
wire n_1975;
wire n_5421;
wire n_4396;
wire n_1990;
wire n_6708;
wire n_6667;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_6040;
wire n_1890;
wire n_6847;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_7251;
wire n_3166;
wire n_7356;
wire n_3649;
wire n_7412;
wire n_3065;
wire n_7212;
wire n_5045;
wire n_5237;
wire n_7060;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_5769;
wire n_2637;
wire n_6750;
wire n_7444;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_7426;
wire n_3953;
wire n_4400;
wire n_7502;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_6855;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_2916;
wire n_7252;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_6543;
wire n_4192;
wire n_6789;
wire n_5972;
wire n_3400;
wire n_7065;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_5146;
wire n_7367;
wire n_7267;
wire n_7405;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_6825;
wire n_1993;
wire n_6460;
wire n_4035;
wire n_6952;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_3060;
wire n_6218;
wire n_6486;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_6852;
wire n_5577;
wire n_5872;
wire n_6692;
wire n_5017;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_7220;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_6888;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_7270;
wire n_4750;
wire n_2348;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_6626;
wire n_4537;
wire n_5838;
wire n_7034;
wire n_3694;
wire n_6854;
wire n_6793;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_6980;
wire n_7040;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_7458;
wire n_4065;
wire n_4705;
wire n_6794;
wire n_1971;
wire n_2945;
wire n_3543;
wire n_7179;
wire n_3448;
wire n_7433;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6334;
wire n_6257;
wire n_4152;
wire n_6874;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_6355;
wire n_7015;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_7226;
wire n_1987;
wire n_7217;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_6377;
wire n_5401;
wire n_4595;
wire n_7272;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_6021;
wire n_4617;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_6511;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_5942;
wire n_5764;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_6867;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_7255;
wire n_3309;
wire n_7181;
wire n_2796;
wire n_5393;
wire n_4817;
wire n_6863;
wire n_7352;
wire n_7355;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_7328;
wire n_2771;
wire n_6322;
wire n_7359;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_3769;
wire n_4437;
wire n_6419;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_7283;
wire n_7089;
wire n_2635;
wire n_2999;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_6417;
wire n_7145;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_6979;
wire n_5986;
wire n_6932;
wire n_2934;
wire n_7258;
wire n_5104;
wire n_6961;
wire n_6792;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_6919;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_7440;
wire n_6831;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_7072;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_3509;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_6458;
wire n_6986;
wire n_3456;
wire n_4532;
wire n_5863;
wire n_6633;
wire n_3790;
wire n_7118;
wire n_6152;
wire n_5734;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_7069;
wire n_5199;
wire n_6546;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_6925;
wire n_7186;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_6428;
wire n_6924;
wire n_3077;
wire n_4944;
wire n_6425;
wire n_3478;
wire n_3062;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_7246;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_7301;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_7262;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_3310;
wire n_2642;
wire n_4423;
wire n_3689;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_6282;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_7059;
wire n_6985;
wire n_4350;
wire n_5600;
wire n_6737;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_5767;
wire n_6459;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_6384;
wire n_4669;
wire n_5228;
wire n_2600;
wire n_7443;
wire n_3436;
wire n_5973;
wire n_7484;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_6753;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_6448;
wire n_5186;
wire n_7487;
wire n_4585;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_7077;
wire n_3686;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_7024;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_6529;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_7214;
wire n_2572;
wire n_4490;
wire n_3677;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_2488;
wire n_6134;
wire n_4158;
wire n_6812;
wire n_3079;
wire n_5190;
wire n_6733;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_6938;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_6212;
wire n_3440;
wire n_6816;
wire n_3658;
wire n_7374;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_7110;
wire n_5714;
wire n_2169;
wire n_6953;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_7086;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_4877;
wire n_2065;
wire n_7038;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_7345;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_2724;
wire n_2258;
wire n_7041;
wire n_6717;
wire n_6881;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_6871;
wire n_2967;
wire n_5343;
wire n_6672;
wire n_6518;
wire n_7334;
wire n_4021;
wire n_6396;
wire n_7028;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_6601;
wire n_2268;
wire n_3469;
wire n_2835;
wire n_5835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_6606;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_6092;
wire n_6462;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_7333;
wire n_3878;
wire n_4197;
wire n_6669;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_7337;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_7439;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_7210;
wire n_3898;
wire n_6228;
wire n_6702;
wire n_7358;
wire n_4749;
wire n_5924;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_6997;
wire n_4238;
wire n_6371;
wire n_2005;
wire n_7187;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_7313;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_6641;
wire n_3845;
wire n_6463;
wire n_3203;
wire n_4986;
wire n_4668;
wire n_6264;
wire n_5782;
wire n_4168;
wire n_7036;
wire n_4298;
wire n_7370;
wire n_4743;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_7480;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_6990;
wire n_5034;
wire n_3312;
wire n_7071;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_3752;
wire n_3672;
wire n_7380;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_7376;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_6409;
wire n_4095;
wire n_5927;
wire n_4485;
wire n_6388;
wire n_3593;
wire n_6839;
wire n_5163;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_6864;
wire n_4890;
wire n_2485;
wire n_6679;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_5507;
wire n_4573;
wire n_4943;
wire n_2875;
wire n_6599;
wire n_3519;
wire n_2209;
wire n_7504;
wire n_4042;
wire n_7099;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_7052;
wire n_6738;
wire n_5226;
wire n_2081;
wire n_6566;
wire n_5696;
wire n_3053;
wire n_5014;
wire n_7106;
wire n_6346;
wire n_3772;
wire n_7408;
wire n_2891;
wire n_4335;
wire n_7026;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_7394;
wire n_4516;
wire n_5235;
wire n_6436;
wire n_2798;
wire n_7450;
wire n_3217;
wire n_6081;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_7462;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_7421;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_6238;
wire n_7025;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_7478;
wire n_3308;
wire n_6326;
wire n_3204;
wire n_7451;
wire n_4134;
wire n_5018;
wire n_6917;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_6612;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_350),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_338),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_707),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_496),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_1328),
.Y(n_1887)
);

CKINVDCx5p33_ASAP7_75t_R g1888 ( 
.A(n_1652),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1593),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1612),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_229),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1575),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1421),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1180),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1047),
.Y(n_1895)
);

BUFx2_ASAP7_75t_L g1896 ( 
.A(n_779),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1595),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_794),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1774),
.Y(n_1899)
);

CKINVDCx5p33_ASAP7_75t_R g1900 ( 
.A(n_1706),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1802),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_23),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1657),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_119),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1598),
.Y(n_1905)
);

BUFx10_ASAP7_75t_L g1906 ( 
.A(n_1297),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_291),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_311),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_80),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_737),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1040),
.Y(n_1911)
);

INVx2_ASAP7_75t_SL g1912 ( 
.A(n_1850),
.Y(n_1912)
);

CKINVDCx5p33_ASAP7_75t_R g1913 ( 
.A(n_1150),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_774),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1779),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1040),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_284),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1681),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1751),
.Y(n_1919)
);

BUFx3_ASAP7_75t_L g1920 ( 
.A(n_1640),
.Y(n_1920)
);

BUFx3_ASAP7_75t_L g1921 ( 
.A(n_1369),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_66),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1678),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1037),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_686),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1251),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1237),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1056),
.Y(n_1928)
);

INVx1_ASAP7_75t_SL g1929 ( 
.A(n_546),
.Y(n_1929)
);

INVx2_ASAP7_75t_SL g1930 ( 
.A(n_1727),
.Y(n_1930)
);

INVx1_ASAP7_75t_SL g1931 ( 
.A(n_848),
.Y(n_1931)
);

CKINVDCx20_ASAP7_75t_R g1932 ( 
.A(n_379),
.Y(n_1932)
);

BUFx8_ASAP7_75t_SL g1933 ( 
.A(n_1336),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1041),
.Y(n_1934)
);

INVx2_ASAP7_75t_SL g1935 ( 
.A(n_1452),
.Y(n_1935)
);

INVxp67_ASAP7_75t_SL g1936 ( 
.A(n_1816),
.Y(n_1936)
);

CKINVDCx5p33_ASAP7_75t_R g1937 ( 
.A(n_1870),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1240),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_800),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1583),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1879),
.Y(n_1941)
);

INVxp67_ASAP7_75t_L g1942 ( 
.A(n_652),
.Y(n_1942)
);

CKINVDCx20_ASAP7_75t_R g1943 ( 
.A(n_1671),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_646),
.Y(n_1944)
);

BUFx10_ASAP7_75t_L g1945 ( 
.A(n_1799),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_998),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1267),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_806),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1632),
.Y(n_1949)
);

CKINVDCx20_ASAP7_75t_R g1950 ( 
.A(n_1385),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1227),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1507),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_810),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_594),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_370),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1513),
.Y(n_1956)
);

BUFx10_ASAP7_75t_L g1957 ( 
.A(n_1182),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_414),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1618),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_917),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_883),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1122),
.Y(n_1962)
);

CKINVDCx20_ASAP7_75t_R g1963 ( 
.A(n_806),
.Y(n_1963)
);

BUFx2_ASAP7_75t_L g1964 ( 
.A(n_1124),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1041),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_422),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_666),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_1634),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1),
.Y(n_1969)
);

BUFx6f_ASAP7_75t_L g1970 ( 
.A(n_1515),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1516),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1704),
.Y(n_1972)
);

CKINVDCx20_ASAP7_75t_R g1973 ( 
.A(n_539),
.Y(n_1973)
);

CKINVDCx5p33_ASAP7_75t_R g1974 ( 
.A(n_1154),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_526),
.Y(n_1975)
);

BUFx10_ASAP7_75t_L g1976 ( 
.A(n_304),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1716),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_624),
.Y(n_1978)
);

BUFx6f_ASAP7_75t_L g1979 ( 
.A(n_1465),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1129),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1189),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1317),
.Y(n_1982)
);

CKINVDCx20_ASAP7_75t_R g1983 ( 
.A(n_243),
.Y(n_1983)
);

HB1xp67_ASAP7_75t_L g1984 ( 
.A(n_515),
.Y(n_1984)
);

CKINVDCx5p33_ASAP7_75t_R g1985 ( 
.A(n_353),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_559),
.Y(n_1986)
);

BUFx3_ASAP7_75t_L g1987 ( 
.A(n_1741),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1812),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1400),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_960),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1509),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1032),
.Y(n_1992)
);

CKINVDCx5p33_ASAP7_75t_R g1993 ( 
.A(n_1819),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_108),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1344),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1839),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1380),
.Y(n_1997)
);

CKINVDCx5p33_ASAP7_75t_R g1998 ( 
.A(n_112),
.Y(n_1998)
);

INVx1_ASAP7_75t_SL g1999 ( 
.A(n_905),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1371),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1471),
.Y(n_2001)
);

CKINVDCx5p33_ASAP7_75t_R g2002 ( 
.A(n_1587),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1693),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1674),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1630),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_575),
.Y(n_2006)
);

CKINVDCx20_ASAP7_75t_R g2007 ( 
.A(n_1164),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1279),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_64),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_351),
.Y(n_2010)
);

CKINVDCx5p33_ASAP7_75t_R g2011 ( 
.A(n_710),
.Y(n_2011)
);

BUFx5_ASAP7_75t_L g2012 ( 
.A(n_766),
.Y(n_2012)
);

CKINVDCx5p33_ASAP7_75t_R g2013 ( 
.A(n_1758),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1361),
.Y(n_2014)
);

CKINVDCx5p33_ASAP7_75t_R g2015 ( 
.A(n_1588),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1212),
.Y(n_2016)
);

BUFx10_ASAP7_75t_L g2017 ( 
.A(n_1178),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1661),
.Y(n_2018)
);

CKINVDCx5p33_ASAP7_75t_R g2019 ( 
.A(n_1455),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_226),
.Y(n_2020)
);

CKINVDCx16_ASAP7_75t_R g2021 ( 
.A(n_1148),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1662),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_998),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1130),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_1732),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_198),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_1661),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_955),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_610),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1719),
.Y(n_2030)
);

CKINVDCx20_ASAP7_75t_R g2031 ( 
.A(n_1517),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_674),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_42),
.Y(n_2033)
);

CKINVDCx20_ASAP7_75t_R g2034 ( 
.A(n_1231),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1167),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_1769),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_1551),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1537),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1339),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_577),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_1319),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1294),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_68),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_596),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1477),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_1682),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_222),
.Y(n_2047)
);

CKINVDCx5p33_ASAP7_75t_R g2048 ( 
.A(n_745),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1538),
.Y(n_2049)
);

CKINVDCx5p33_ASAP7_75t_R g2050 ( 
.A(n_531),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_133),
.Y(n_2051)
);

CKINVDCx5p33_ASAP7_75t_R g2052 ( 
.A(n_1170),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_650),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_762),
.Y(n_2054)
);

BUFx2_ASAP7_75t_L g2055 ( 
.A(n_1468),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1234),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1246),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_130),
.Y(n_2058)
);

BUFx10_ASAP7_75t_L g2059 ( 
.A(n_1338),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_1781),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1840),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1604),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1781),
.Y(n_2063)
);

CKINVDCx20_ASAP7_75t_R g2064 ( 
.A(n_924),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_89),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1080),
.Y(n_2066)
);

CKINVDCx5p33_ASAP7_75t_R g2067 ( 
.A(n_506),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_174),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1806),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1453),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1129),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1221),
.Y(n_2072)
);

CKINVDCx5p33_ASAP7_75t_R g2073 ( 
.A(n_1518),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1846),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_290),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_1191),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_827),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_945),
.Y(n_2078)
);

CKINVDCx5p33_ASAP7_75t_R g2079 ( 
.A(n_1708),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1852),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1363),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1687),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_1286),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_643),
.Y(n_2084)
);

CKINVDCx5p33_ASAP7_75t_R g2085 ( 
.A(n_1559),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_1686),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_22),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_26),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_469),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1790),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1408),
.Y(n_2091)
);

CKINVDCx5p33_ASAP7_75t_R g2092 ( 
.A(n_1035),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_983),
.Y(n_2093)
);

CKINVDCx5p33_ASAP7_75t_R g2094 ( 
.A(n_1106),
.Y(n_2094)
);

CKINVDCx20_ASAP7_75t_R g2095 ( 
.A(n_1388),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1729),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1872),
.Y(n_2097)
);

CKINVDCx5p33_ASAP7_75t_R g2098 ( 
.A(n_803),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1295),
.Y(n_2099)
);

CKINVDCx16_ASAP7_75t_R g2100 ( 
.A(n_241),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1180),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_539),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1120),
.Y(n_2103)
);

CKINVDCx20_ASAP7_75t_R g2104 ( 
.A(n_1406),
.Y(n_2104)
);

CKINVDCx5p33_ASAP7_75t_R g2105 ( 
.A(n_641),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_957),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1598),
.Y(n_2107)
);

CKINVDCx5p33_ASAP7_75t_R g2108 ( 
.A(n_1361),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1725),
.Y(n_2109)
);

CKINVDCx5p33_ASAP7_75t_R g2110 ( 
.A(n_1202),
.Y(n_2110)
);

CKINVDCx5p33_ASAP7_75t_R g2111 ( 
.A(n_612),
.Y(n_2111)
);

INVx1_ASAP7_75t_SL g2112 ( 
.A(n_1163),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_157),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1705),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1721),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1756),
.Y(n_2116)
);

CKINVDCx5p33_ASAP7_75t_R g2117 ( 
.A(n_546),
.Y(n_2117)
);

CKINVDCx5p33_ASAP7_75t_R g2118 ( 
.A(n_1808),
.Y(n_2118)
);

CKINVDCx20_ASAP7_75t_R g2119 ( 
.A(n_1167),
.Y(n_2119)
);

CKINVDCx5p33_ASAP7_75t_R g2120 ( 
.A(n_1214),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_631),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1552),
.Y(n_2122)
);

CKINVDCx5p33_ASAP7_75t_R g2123 ( 
.A(n_1702),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_352),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_108),
.Y(n_2125)
);

CKINVDCx5p33_ASAP7_75t_R g2126 ( 
.A(n_1855),
.Y(n_2126)
);

CKINVDCx5p33_ASAP7_75t_R g2127 ( 
.A(n_475),
.Y(n_2127)
);

INVx1_ASAP7_75t_SL g2128 ( 
.A(n_703),
.Y(n_2128)
);

CKINVDCx5p33_ASAP7_75t_R g2129 ( 
.A(n_132),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1668),
.Y(n_2130)
);

CKINVDCx5p33_ASAP7_75t_R g2131 ( 
.A(n_1734),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1172),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1085),
.Y(n_2133)
);

CKINVDCx5p33_ASAP7_75t_R g2134 ( 
.A(n_1643),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1777),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_82),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_838),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_730),
.Y(n_2138)
);

CKINVDCx5p33_ASAP7_75t_R g2139 ( 
.A(n_1711),
.Y(n_2139)
);

CKINVDCx20_ASAP7_75t_R g2140 ( 
.A(n_1770),
.Y(n_2140)
);

BUFx8_ASAP7_75t_SL g2141 ( 
.A(n_1701),
.Y(n_2141)
);

CKINVDCx14_ASAP7_75t_R g2142 ( 
.A(n_1281),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_202),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1736),
.Y(n_2144)
);

CKINVDCx14_ASAP7_75t_R g2145 ( 
.A(n_1079),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_757),
.Y(n_2146)
);

CKINVDCx5p33_ASAP7_75t_R g2147 ( 
.A(n_1309),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1714),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_142),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_23),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_832),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_472),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_224),
.Y(n_2153)
);

BUFx2_ASAP7_75t_L g2154 ( 
.A(n_565),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1127),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1719),
.Y(n_2156)
);

CKINVDCx5p33_ASAP7_75t_R g2157 ( 
.A(n_1603),
.Y(n_2157)
);

CKINVDCx20_ASAP7_75t_R g2158 ( 
.A(n_991),
.Y(n_2158)
);

CKINVDCx5p33_ASAP7_75t_R g2159 ( 
.A(n_1645),
.Y(n_2159)
);

BUFx3_ASAP7_75t_L g2160 ( 
.A(n_1152),
.Y(n_2160)
);

CKINVDCx5p33_ASAP7_75t_R g2161 ( 
.A(n_1760),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_139),
.Y(n_2162)
);

CKINVDCx5p33_ASAP7_75t_R g2163 ( 
.A(n_944),
.Y(n_2163)
);

BUFx10_ASAP7_75t_L g2164 ( 
.A(n_359),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_709),
.Y(n_2165)
);

INVx1_ASAP7_75t_SL g2166 ( 
.A(n_406),
.Y(n_2166)
);

CKINVDCx5p33_ASAP7_75t_R g2167 ( 
.A(n_241),
.Y(n_2167)
);

BUFx2_ASAP7_75t_L g2168 ( 
.A(n_552),
.Y(n_2168)
);

CKINVDCx20_ASAP7_75t_R g2169 ( 
.A(n_1825),
.Y(n_2169)
);

CKINVDCx5p33_ASAP7_75t_R g2170 ( 
.A(n_764),
.Y(n_2170)
);

INVx1_ASAP7_75t_SL g2171 ( 
.A(n_717),
.Y(n_2171)
);

INVx1_ASAP7_75t_SL g2172 ( 
.A(n_648),
.Y(n_2172)
);

CKINVDCx5p33_ASAP7_75t_R g2173 ( 
.A(n_761),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_163),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_906),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_228),
.Y(n_2176)
);

INVx1_ASAP7_75t_SL g2177 ( 
.A(n_28),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1132),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_372),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_1754),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1196),
.Y(n_2181)
);

CKINVDCx5p33_ASAP7_75t_R g2182 ( 
.A(n_798),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1408),
.Y(n_2183)
);

INVxp33_ASAP7_75t_SL g2184 ( 
.A(n_238),
.Y(n_2184)
);

CKINVDCx20_ASAP7_75t_R g2185 ( 
.A(n_1665),
.Y(n_2185)
);

CKINVDCx20_ASAP7_75t_R g2186 ( 
.A(n_688),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1021),
.Y(n_2187)
);

CKINVDCx5p33_ASAP7_75t_R g2188 ( 
.A(n_1747),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_109),
.Y(n_2189)
);

CKINVDCx5p33_ASAP7_75t_R g2190 ( 
.A(n_1853),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_518),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1223),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1680),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_349),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_1094),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1755),
.Y(n_2196)
);

CKINVDCx5p33_ASAP7_75t_R g2197 ( 
.A(n_8),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_607),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_778),
.Y(n_2199)
);

CKINVDCx5p33_ASAP7_75t_R g2200 ( 
.A(n_809),
.Y(n_2200)
);

CKINVDCx5p33_ASAP7_75t_R g2201 ( 
.A(n_1345),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1031),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1321),
.Y(n_2203)
);

CKINVDCx5p33_ASAP7_75t_R g2204 ( 
.A(n_580),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1601),
.Y(n_2205)
);

CKINVDCx16_ASAP7_75t_R g2206 ( 
.A(n_612),
.Y(n_2206)
);

CKINVDCx5p33_ASAP7_75t_R g2207 ( 
.A(n_1284),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_245),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_1228),
.Y(n_2209)
);

CKINVDCx5p33_ASAP7_75t_R g2210 ( 
.A(n_1269),
.Y(n_2210)
);

CKINVDCx5p33_ASAP7_75t_R g2211 ( 
.A(n_1432),
.Y(n_2211)
);

BUFx2_ASAP7_75t_L g2212 ( 
.A(n_419),
.Y(n_2212)
);

CKINVDCx5p33_ASAP7_75t_R g2213 ( 
.A(n_1214),
.Y(n_2213)
);

BUFx2_ASAP7_75t_L g2214 ( 
.A(n_1608),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_611),
.Y(n_2215)
);

CKINVDCx5p33_ASAP7_75t_R g2216 ( 
.A(n_1316),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1061),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_409),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_417),
.Y(n_2219)
);

BUFx10_ASAP7_75t_L g2220 ( 
.A(n_1725),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1160),
.Y(n_2221)
);

BUFx3_ASAP7_75t_L g2222 ( 
.A(n_421),
.Y(n_2222)
);

CKINVDCx20_ASAP7_75t_R g2223 ( 
.A(n_26),
.Y(n_2223)
);

CKINVDCx5p33_ASAP7_75t_R g2224 ( 
.A(n_1700),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_1337),
.Y(n_2225)
);

CKINVDCx16_ASAP7_75t_R g2226 ( 
.A(n_500),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_371),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1012),
.Y(n_2228)
);

HB1xp67_ASAP7_75t_L g2229 ( 
.A(n_1843),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_1241),
.Y(n_2230)
);

BUFx5_ASAP7_75t_L g2231 ( 
.A(n_782),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_301),
.Y(n_2232)
);

CKINVDCx5p33_ASAP7_75t_R g2233 ( 
.A(n_870),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_877),
.Y(n_2234)
);

CKINVDCx20_ASAP7_75t_R g2235 ( 
.A(n_1481),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_526),
.Y(n_2236)
);

CKINVDCx5p33_ASAP7_75t_R g2237 ( 
.A(n_1717),
.Y(n_2237)
);

INVx1_ASAP7_75t_SL g2238 ( 
.A(n_754),
.Y(n_2238)
);

CKINVDCx20_ASAP7_75t_R g2239 ( 
.A(n_984),
.Y(n_2239)
);

HB1xp67_ASAP7_75t_L g2240 ( 
.A(n_550),
.Y(n_2240)
);

CKINVDCx5p33_ASAP7_75t_R g2241 ( 
.A(n_1679),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_304),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1763),
.Y(n_2243)
);

BUFx3_ASAP7_75t_L g2244 ( 
.A(n_1629),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_182),
.Y(n_2245)
);

CKINVDCx5p33_ASAP7_75t_R g2246 ( 
.A(n_1628),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_837),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1256),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_306),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1740),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_1689),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_1307),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_1221),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_877),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1375),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_655),
.Y(n_2256)
);

BUFx10_ASAP7_75t_L g2257 ( 
.A(n_874),
.Y(n_2257)
);

CKINVDCx5p33_ASAP7_75t_R g2258 ( 
.A(n_1847),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_626),
.Y(n_2259)
);

CKINVDCx5p33_ASAP7_75t_R g2260 ( 
.A(n_98),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_880),
.Y(n_2261)
);

INVxp67_ASAP7_75t_SL g2262 ( 
.A(n_1777),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_188),
.Y(n_2263)
);

CKINVDCx5p33_ASAP7_75t_R g2264 ( 
.A(n_613),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1366),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_1215),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_445),
.Y(n_2267)
);

INVx1_ASAP7_75t_SL g2268 ( 
.A(n_1782),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_734),
.Y(n_2269)
);

CKINVDCx5p33_ASAP7_75t_R g2270 ( 
.A(n_1762),
.Y(n_2270)
);

CKINVDCx5p33_ASAP7_75t_R g2271 ( 
.A(n_27),
.Y(n_2271)
);

CKINVDCx5p33_ASAP7_75t_R g2272 ( 
.A(n_190),
.Y(n_2272)
);

CKINVDCx20_ASAP7_75t_R g2273 ( 
.A(n_952),
.Y(n_2273)
);

CKINVDCx14_ASAP7_75t_R g2274 ( 
.A(n_1267),
.Y(n_2274)
);

CKINVDCx5p33_ASAP7_75t_R g2275 ( 
.A(n_1739),
.Y(n_2275)
);

CKINVDCx5p33_ASAP7_75t_R g2276 ( 
.A(n_838),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1627),
.Y(n_2277)
);

CKINVDCx5p33_ASAP7_75t_R g2278 ( 
.A(n_520),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_1060),
.Y(n_2279)
);

BUFx3_ASAP7_75t_L g2280 ( 
.A(n_336),
.Y(n_2280)
);

CKINVDCx5p33_ASAP7_75t_R g2281 ( 
.A(n_1471),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_459),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1454),
.Y(n_2283)
);

CKINVDCx16_ASAP7_75t_R g2284 ( 
.A(n_1624),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_39),
.Y(n_2285)
);

CKINVDCx5p33_ASAP7_75t_R g2286 ( 
.A(n_1132),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_1035),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_1304),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_143),
.Y(n_2289)
);

CKINVDCx5p33_ASAP7_75t_R g2290 ( 
.A(n_1001),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_1505),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1791),
.Y(n_2292)
);

CKINVDCx20_ASAP7_75t_R g2293 ( 
.A(n_1477),
.Y(n_2293)
);

INVx1_ASAP7_75t_SL g2294 ( 
.A(n_1858),
.Y(n_2294)
);

CKINVDCx5p33_ASAP7_75t_R g2295 ( 
.A(n_1555),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1280),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1583),
.Y(n_2297)
);

CKINVDCx14_ASAP7_75t_R g2298 ( 
.A(n_1742),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_214),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_1106),
.Y(n_2300)
);

CKINVDCx5p33_ASAP7_75t_R g2301 ( 
.A(n_904),
.Y(n_2301)
);

CKINVDCx5p33_ASAP7_75t_R g2302 ( 
.A(n_1666),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_472),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1856),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_185),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_441),
.Y(n_2306)
);

CKINVDCx5p33_ASAP7_75t_R g2307 ( 
.A(n_62),
.Y(n_2307)
);

BUFx2_ASAP7_75t_L g2308 ( 
.A(n_1192),
.Y(n_2308)
);

CKINVDCx5p33_ASAP7_75t_R g2309 ( 
.A(n_586),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1535),
.Y(n_2310)
);

INVx1_ASAP7_75t_SL g2311 ( 
.A(n_1094),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_557),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1382),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_1312),
.Y(n_2314)
);

BUFx5_ASAP7_75t_L g2315 ( 
.A(n_1808),
.Y(n_2315)
);

CKINVDCx5p33_ASAP7_75t_R g2316 ( 
.A(n_1723),
.Y(n_2316)
);

CKINVDCx5p33_ASAP7_75t_R g2317 ( 
.A(n_1654),
.Y(n_2317)
);

CKINVDCx20_ASAP7_75t_R g2318 ( 
.A(n_296),
.Y(n_2318)
);

CKINVDCx5p33_ASAP7_75t_R g2319 ( 
.A(n_209),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_940),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_876),
.Y(n_2321)
);

CKINVDCx5p33_ASAP7_75t_R g2322 ( 
.A(n_1712),
.Y(n_2322)
);

CKINVDCx5p33_ASAP7_75t_R g2323 ( 
.A(n_1849),
.Y(n_2323)
);

CKINVDCx5p33_ASAP7_75t_R g2324 ( 
.A(n_469),
.Y(n_2324)
);

CKINVDCx5p33_ASAP7_75t_R g2325 ( 
.A(n_1746),
.Y(n_2325)
);

CKINVDCx5p33_ASAP7_75t_R g2326 ( 
.A(n_1633),
.Y(n_2326)
);

BUFx10_ASAP7_75t_L g2327 ( 
.A(n_1090),
.Y(n_2327)
);

CKINVDCx20_ASAP7_75t_R g2328 ( 
.A(n_1213),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_1343),
.Y(n_2329)
);

BUFx10_ASAP7_75t_L g2330 ( 
.A(n_433),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1096),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_1754),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1333),
.Y(n_2333)
);

CKINVDCx5p33_ASAP7_75t_R g2334 ( 
.A(n_1735),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_950),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_345),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_1823),
.Y(n_2337)
);

CKINVDCx5p33_ASAP7_75t_R g2338 ( 
.A(n_129),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1177),
.Y(n_2339)
);

BUFx2_ASAP7_75t_L g2340 ( 
.A(n_281),
.Y(n_2340)
);

CKINVDCx20_ASAP7_75t_R g2341 ( 
.A(n_46),
.Y(n_2341)
);

CKINVDCx5p33_ASAP7_75t_R g2342 ( 
.A(n_1196),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_1734),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_396),
.Y(n_2344)
);

CKINVDCx5p33_ASAP7_75t_R g2345 ( 
.A(n_786),
.Y(n_2345)
);

CKINVDCx5p33_ASAP7_75t_R g2346 ( 
.A(n_122),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_455),
.Y(n_2347)
);

CKINVDCx5p33_ASAP7_75t_R g2348 ( 
.A(n_1100),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1768),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1062),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_28),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_1761),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_979),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_663),
.Y(n_2354)
);

INVx1_ASAP7_75t_SL g2355 ( 
.A(n_740),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_1113),
.Y(n_2356)
);

CKINVDCx5p33_ASAP7_75t_R g2357 ( 
.A(n_986),
.Y(n_2357)
);

CKINVDCx5p33_ASAP7_75t_R g2358 ( 
.A(n_693),
.Y(n_2358)
);

CKINVDCx5p33_ASAP7_75t_R g2359 ( 
.A(n_497),
.Y(n_2359)
);

CKINVDCx5p33_ASAP7_75t_R g2360 ( 
.A(n_759),
.Y(n_2360)
);

INVxp67_ASAP7_75t_L g2361 ( 
.A(n_409),
.Y(n_2361)
);

CKINVDCx5p33_ASAP7_75t_R g2362 ( 
.A(n_99),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_1339),
.Y(n_2363)
);

CKINVDCx5p33_ASAP7_75t_R g2364 ( 
.A(n_234),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_1650),
.Y(n_2365)
);

CKINVDCx20_ASAP7_75t_R g2366 ( 
.A(n_1818),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_770),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_198),
.Y(n_2368)
);

CKINVDCx5p33_ASAP7_75t_R g2369 ( 
.A(n_182),
.Y(n_2369)
);

CKINVDCx5p33_ASAP7_75t_R g2370 ( 
.A(n_375),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_1104),
.Y(n_2371)
);

CKINVDCx5p33_ASAP7_75t_R g2372 ( 
.A(n_449),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_459),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_566),
.Y(n_2374)
);

CKINVDCx5p33_ASAP7_75t_R g2375 ( 
.A(n_1574),
.Y(n_2375)
);

CKINVDCx5p33_ASAP7_75t_R g2376 ( 
.A(n_307),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1349),
.Y(n_2377)
);

CKINVDCx5p33_ASAP7_75t_R g2378 ( 
.A(n_1204),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_1706),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_826),
.Y(n_2380)
);

CKINVDCx5p33_ASAP7_75t_R g2381 ( 
.A(n_1629),
.Y(n_2381)
);

BUFx3_ASAP7_75t_L g2382 ( 
.A(n_1234),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_474),
.Y(n_2383)
);

HB1xp67_ASAP7_75t_L g2384 ( 
.A(n_348),
.Y(n_2384)
);

CKINVDCx5p33_ASAP7_75t_R g2385 ( 
.A(n_1),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1744),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_687),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1056),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1694),
.Y(n_2389)
);

CKINVDCx5p33_ASAP7_75t_R g2390 ( 
.A(n_1519),
.Y(n_2390)
);

CKINVDCx5p33_ASAP7_75t_R g2391 ( 
.A(n_525),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_72),
.Y(n_2392)
);

BUFx10_ASAP7_75t_L g2393 ( 
.A(n_967),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_239),
.Y(n_2394)
);

INVx1_ASAP7_75t_SL g2395 ( 
.A(n_1053),
.Y(n_2395)
);

CKINVDCx5p33_ASAP7_75t_R g2396 ( 
.A(n_684),
.Y(n_2396)
);

CKINVDCx5p33_ASAP7_75t_R g2397 ( 
.A(n_1690),
.Y(n_2397)
);

CKINVDCx5p33_ASAP7_75t_R g2398 ( 
.A(n_1421),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_865),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_959),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_358),
.Y(n_2401)
);

INVxp33_ASAP7_75t_L g2402 ( 
.A(n_142),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_227),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_333),
.Y(n_2404)
);

CKINVDCx5p33_ASAP7_75t_R g2405 ( 
.A(n_498),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_572),
.Y(n_2406)
);

CKINVDCx5p33_ASAP7_75t_R g2407 ( 
.A(n_624),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_78),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_79),
.Y(n_2409)
);

CKINVDCx5p33_ASAP7_75t_R g2410 ( 
.A(n_225),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_1036),
.Y(n_2411)
);

CKINVDCx20_ASAP7_75t_R g2412 ( 
.A(n_1857),
.Y(n_2412)
);

CKINVDCx5p33_ASAP7_75t_R g2413 ( 
.A(n_1575),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_1685),
.Y(n_2414)
);

INVx1_ASAP7_75t_SL g2415 ( 
.A(n_1362),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_1248),
.Y(n_2416)
);

BUFx5_ASAP7_75t_L g2417 ( 
.A(n_870),
.Y(n_2417)
);

CKINVDCx20_ASAP7_75t_R g2418 ( 
.A(n_1183),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_458),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_1619),
.Y(n_2420)
);

CKINVDCx5p33_ASAP7_75t_R g2421 ( 
.A(n_1696),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1465),
.Y(n_2422)
);

CKINVDCx5p33_ASAP7_75t_R g2423 ( 
.A(n_130),
.Y(n_2423)
);

CKINVDCx16_ASAP7_75t_R g2424 ( 
.A(n_622),
.Y(n_2424)
);

CKINVDCx5p33_ASAP7_75t_R g2425 ( 
.A(n_1332),
.Y(n_2425)
);

CKINVDCx5p33_ASAP7_75t_R g2426 ( 
.A(n_1329),
.Y(n_2426)
);

BUFx10_ASAP7_75t_L g2427 ( 
.A(n_118),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_99),
.Y(n_2428)
);

CKINVDCx5p33_ASAP7_75t_R g2429 ( 
.A(n_1703),
.Y(n_2429)
);

INVx2_ASAP7_75t_SL g2430 ( 
.A(n_448),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_1811),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1144),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_380),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_934),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_355),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_603),
.Y(n_2436)
);

CKINVDCx20_ASAP7_75t_R g2437 ( 
.A(n_654),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_1493),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1347),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_66),
.Y(n_2440)
);

CKINVDCx5p33_ASAP7_75t_R g2441 ( 
.A(n_904),
.Y(n_2441)
);

CKINVDCx5p33_ASAP7_75t_R g2442 ( 
.A(n_323),
.Y(n_2442)
);

CKINVDCx5p33_ASAP7_75t_R g2443 ( 
.A(n_449),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_674),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_962),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_1547),
.Y(n_2446)
);

CKINVDCx5p33_ASAP7_75t_R g2447 ( 
.A(n_1769),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1426),
.Y(n_2448)
);

CKINVDCx5p33_ASAP7_75t_R g2449 ( 
.A(n_36),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_1677),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_557),
.Y(n_2451)
);

INVx2_ASAP7_75t_SL g2452 ( 
.A(n_852),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_981),
.Y(n_2453)
);

CKINVDCx5p33_ASAP7_75t_R g2454 ( 
.A(n_1788),
.Y(n_2454)
);

INVx2_ASAP7_75t_SL g2455 ( 
.A(n_599),
.Y(n_2455)
);

CKINVDCx5p33_ASAP7_75t_R g2456 ( 
.A(n_166),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_248),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_919),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_1154),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_1684),
.Y(n_2460)
);

CKINVDCx5p33_ASAP7_75t_R g2461 ( 
.A(n_625),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_301),
.Y(n_2462)
);

CKINVDCx5p33_ASAP7_75t_R g2463 ( 
.A(n_891),
.Y(n_2463)
);

BUFx3_ASAP7_75t_L g2464 ( 
.A(n_1767),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_59),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_1812),
.Y(n_2466)
);

CKINVDCx5p33_ASAP7_75t_R g2467 ( 
.A(n_1420),
.Y(n_2467)
);

CKINVDCx14_ASAP7_75t_R g2468 ( 
.A(n_1683),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_1710),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_1748),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_187),
.Y(n_2471)
);

BUFx3_ASAP7_75t_L g2472 ( 
.A(n_321),
.Y(n_2472)
);

CKINVDCx5p33_ASAP7_75t_R g2473 ( 
.A(n_1324),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_123),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_1564),
.Y(n_2475)
);

INVx3_ASAP7_75t_L g2476 ( 
.A(n_508),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_1282),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_51),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_1649),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_1730),
.Y(n_2480)
);

HB1xp67_ASAP7_75t_L g2481 ( 
.A(n_627),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_343),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_306),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_1656),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_842),
.Y(n_2485)
);

CKINVDCx5p33_ASAP7_75t_R g2486 ( 
.A(n_1663),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_437),
.Y(n_2487)
);

CKINVDCx5p33_ASAP7_75t_R g2488 ( 
.A(n_1723),
.Y(n_2488)
);

CKINVDCx5p33_ASAP7_75t_R g2489 ( 
.A(n_390),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_1220),
.Y(n_2490)
);

CKINVDCx5p33_ASAP7_75t_R g2491 ( 
.A(n_1750),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1655),
.Y(n_2492)
);

CKINVDCx20_ASAP7_75t_R g2493 ( 
.A(n_1869),
.Y(n_2493)
);

CKINVDCx20_ASAP7_75t_R g2494 ( 
.A(n_1715),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_621),
.Y(n_2495)
);

INVx1_ASAP7_75t_L g2496 ( 
.A(n_1311),
.Y(n_2496)
);

CKINVDCx20_ASAP7_75t_R g2497 ( 
.A(n_319),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_1435),
.Y(n_2498)
);

CKINVDCx5p33_ASAP7_75t_R g2499 ( 
.A(n_1775),
.Y(n_2499)
);

CKINVDCx20_ASAP7_75t_R g2500 ( 
.A(n_1673),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_1628),
.Y(n_2501)
);

CKINVDCx5p33_ASAP7_75t_R g2502 ( 
.A(n_1712),
.Y(n_2502)
);

CKINVDCx5p33_ASAP7_75t_R g2503 ( 
.A(n_1091),
.Y(n_2503)
);

BUFx4f_ASAP7_75t_SL g2504 ( 
.A(n_1260),
.Y(n_2504)
);

CKINVDCx5p33_ASAP7_75t_R g2505 ( 
.A(n_1743),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_1286),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_349),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_1618),
.Y(n_2508)
);

INVx1_ASAP7_75t_SL g2509 ( 
.A(n_1255),
.Y(n_2509)
);

CKINVDCx5p33_ASAP7_75t_R g2510 ( 
.A(n_1315),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_129),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_1244),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_1764),
.Y(n_2513)
);

CKINVDCx20_ASAP7_75t_R g2514 ( 
.A(n_822),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_618),
.Y(n_2515)
);

CKINVDCx5p33_ASAP7_75t_R g2516 ( 
.A(n_124),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_1336),
.Y(n_2517)
);

INVx1_ASAP7_75t_SL g2518 ( 
.A(n_504),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_1261),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_1561),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_1875),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_443),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_1255),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_215),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_91),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_1105),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_1658),
.Y(n_2527)
);

CKINVDCx5p33_ASAP7_75t_R g2528 ( 
.A(n_910),
.Y(n_2528)
);

CKINVDCx5p33_ASAP7_75t_R g2529 ( 
.A(n_746),
.Y(n_2529)
);

CKINVDCx16_ASAP7_75t_R g2530 ( 
.A(n_565),
.Y(n_2530)
);

CKINVDCx5p33_ASAP7_75t_R g2531 ( 
.A(n_1707),
.Y(n_2531)
);

CKINVDCx20_ASAP7_75t_R g2532 ( 
.A(n_1202),
.Y(n_2532)
);

CKINVDCx5p33_ASAP7_75t_R g2533 ( 
.A(n_649),
.Y(n_2533)
);

CKINVDCx20_ASAP7_75t_R g2534 ( 
.A(n_1881),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_1147),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_1638),
.Y(n_2536)
);

CKINVDCx20_ASAP7_75t_R g2537 ( 
.A(n_25),
.Y(n_2537)
);

INVx1_ASAP7_75t_SL g2538 ( 
.A(n_1692),
.Y(n_2538)
);

CKINVDCx5p33_ASAP7_75t_R g2539 ( 
.A(n_1697),
.Y(n_2539)
);

BUFx3_ASAP7_75t_L g2540 ( 
.A(n_1381),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_817),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_1617),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_208),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_1660),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_676),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_372),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_512),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_584),
.Y(n_2548)
);

CKINVDCx5p33_ASAP7_75t_R g2549 ( 
.A(n_1713),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_1659),
.Y(n_2550)
);

CKINVDCx20_ASAP7_75t_R g2551 ( 
.A(n_410),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_1728),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_1825),
.Y(n_2553)
);

CKINVDCx5p33_ASAP7_75t_R g2554 ( 
.A(n_1784),
.Y(n_2554)
);

CKINVDCx5p33_ASAP7_75t_R g2555 ( 
.A(n_225),
.Y(n_2555)
);

BUFx2_ASAP7_75t_L g2556 ( 
.A(n_276),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1824),
.Y(n_2557)
);

CKINVDCx5p33_ASAP7_75t_R g2558 ( 
.A(n_208),
.Y(n_2558)
);

CKINVDCx5p33_ASAP7_75t_R g2559 ( 
.A(n_1765),
.Y(n_2559)
);

CKINVDCx5p33_ASAP7_75t_R g2560 ( 
.A(n_718),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_1469),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_1183),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_638),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_749),
.Y(n_2564)
);

CKINVDCx16_ASAP7_75t_R g2565 ( 
.A(n_194),
.Y(n_2565)
);

CKINVDCx5p33_ASAP7_75t_R g2566 ( 
.A(n_1206),
.Y(n_2566)
);

CKINVDCx5p33_ASAP7_75t_R g2567 ( 
.A(n_809),
.Y(n_2567)
);

CKINVDCx5p33_ASAP7_75t_R g2568 ( 
.A(n_1757),
.Y(n_2568)
);

CKINVDCx5p33_ASAP7_75t_R g2569 ( 
.A(n_1228),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_1672),
.Y(n_2570)
);

CKINVDCx5p33_ASAP7_75t_R g2571 ( 
.A(n_589),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_423),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_582),
.Y(n_2573)
);

CKINVDCx5p33_ASAP7_75t_R g2574 ( 
.A(n_1177),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_243),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_1867),
.Y(n_2576)
);

BUFx10_ASAP7_75t_L g2577 ( 
.A(n_1508),
.Y(n_2577)
);

CKINVDCx5p33_ASAP7_75t_R g2578 ( 
.A(n_1491),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_1771),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_1637),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_1676),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_1220),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_295),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_1742),
.Y(n_2584)
);

CKINVDCx5p33_ASAP7_75t_R g2585 ( 
.A(n_958),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_67),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_1720),
.Y(n_2587)
);

CKINVDCx5p33_ASAP7_75t_R g2588 ( 
.A(n_1561),
.Y(n_2588)
);

CKINVDCx20_ASAP7_75t_R g2589 ( 
.A(n_491),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_650),
.Y(n_2590)
);

CKINVDCx5p33_ASAP7_75t_R g2591 ( 
.A(n_1245),
.Y(n_2591)
);

BUFx2_ASAP7_75t_L g2592 ( 
.A(n_1085),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_1142),
.Y(n_2593)
);

CKINVDCx16_ASAP7_75t_R g2594 ( 
.A(n_1092),
.Y(n_2594)
);

CKINVDCx5p33_ASAP7_75t_R g2595 ( 
.A(n_486),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1414),
.Y(n_2596)
);

BUFx3_ASAP7_75t_L g2597 ( 
.A(n_1726),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_413),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_731),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_1731),
.Y(n_2600)
);

INVx1_ASAP7_75t_SL g2601 ( 
.A(n_256),
.Y(n_2601)
);

BUFx6f_ASAP7_75t_L g2602 ( 
.A(n_1675),
.Y(n_2602)
);

INVx1_ASAP7_75t_SL g2603 ( 
.A(n_1378),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_968),
.Y(n_2604)
);

CKINVDCx5p33_ASAP7_75t_R g2605 ( 
.A(n_1445),
.Y(n_2605)
);

CKINVDCx5p33_ASAP7_75t_R g2606 ( 
.A(n_216),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_1688),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_1190),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_1880),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_567),
.Y(n_2610)
);

CKINVDCx5p33_ASAP7_75t_R g2611 ( 
.A(n_1759),
.Y(n_2611)
);

CKINVDCx5p33_ASAP7_75t_R g2612 ( 
.A(n_79),
.Y(n_2612)
);

CKINVDCx5p33_ASAP7_75t_R g2613 ( 
.A(n_978),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_447),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_489),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_793),
.Y(n_2616)
);

INVx3_ASAP7_75t_L g2617 ( 
.A(n_1815),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_327),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_561),
.Y(n_2619)
);

CKINVDCx5p33_ASAP7_75t_R g2620 ( 
.A(n_158),
.Y(n_2620)
);

CKINVDCx16_ASAP7_75t_R g2621 ( 
.A(n_20),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_1589),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_735),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_1547),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_1584),
.Y(n_2625)
);

CKINVDCx5p33_ASAP7_75t_R g2626 ( 
.A(n_1641),
.Y(n_2626)
);

CKINVDCx5p33_ASAP7_75t_R g2627 ( 
.A(n_1420),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_1653),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_711),
.Y(n_2629)
);

CKINVDCx20_ASAP7_75t_R g2630 ( 
.A(n_646),
.Y(n_2630)
);

CKINVDCx5p33_ASAP7_75t_R g2631 ( 
.A(n_1845),
.Y(n_2631)
);

CKINVDCx5p33_ASAP7_75t_R g2632 ( 
.A(n_1749),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_405),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_1046),
.Y(n_2634)
);

INVxp67_ASAP7_75t_SL g2635 ( 
.A(n_1069),
.Y(n_2635)
);

INVx2_ASAP7_75t_SL g2636 ( 
.A(n_1621),
.Y(n_2636)
);

CKINVDCx5p33_ASAP7_75t_R g2637 ( 
.A(n_608),
.Y(n_2637)
);

CKINVDCx5p33_ASAP7_75t_R g2638 ( 
.A(n_804),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_1580),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_1597),
.Y(n_2640)
);

BUFx10_ASAP7_75t_L g2641 ( 
.A(n_1038),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_1483),
.Y(n_2642)
);

BUFx3_ASAP7_75t_L g2643 ( 
.A(n_701),
.Y(n_2643)
);

INVx2_ASAP7_75t_SL g2644 ( 
.A(n_470),
.Y(n_2644)
);

CKINVDCx5p33_ASAP7_75t_R g2645 ( 
.A(n_354),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_1814),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_480),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_883),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_709),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_819),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_1745),
.Y(n_2651)
);

CKINVDCx5p33_ASAP7_75t_R g2652 ( 
.A(n_1640),
.Y(n_2652)
);

CKINVDCx5p33_ASAP7_75t_R g2653 ( 
.A(n_1749),
.Y(n_2653)
);

CKINVDCx20_ASAP7_75t_R g2654 ( 
.A(n_1452),
.Y(n_2654)
);

BUFx10_ASAP7_75t_L g2655 ( 
.A(n_1800),
.Y(n_2655)
);

CKINVDCx5p33_ASAP7_75t_R g2656 ( 
.A(n_1176),
.Y(n_2656)
);

CKINVDCx5p33_ASAP7_75t_R g2657 ( 
.A(n_371),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_778),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_1667),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_981),
.Y(n_2660)
);

CKINVDCx5p33_ASAP7_75t_R g2661 ( 
.A(n_496),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_869),
.Y(n_2662)
);

CKINVDCx5p33_ASAP7_75t_R g2663 ( 
.A(n_1644),
.Y(n_2663)
);

CKINVDCx5p33_ASAP7_75t_R g2664 ( 
.A(n_470),
.Y(n_2664)
);

CKINVDCx20_ASAP7_75t_R g2665 ( 
.A(n_1474),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_6),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_1635),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_1432),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_1766),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_1709),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_228),
.Y(n_2671)
);

CKINVDCx5p33_ASAP7_75t_R g2672 ( 
.A(n_1568),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_450),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_1484),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_1171),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_1705),
.Y(n_2676)
);

HB1xp67_ASAP7_75t_L g2677 ( 
.A(n_1698),
.Y(n_2677)
);

CKINVDCx5p33_ASAP7_75t_R g2678 ( 
.A(n_454),
.Y(n_2678)
);

CKINVDCx20_ASAP7_75t_R g2679 ( 
.A(n_1072),
.Y(n_2679)
);

BUFx2_ASAP7_75t_SL g2680 ( 
.A(n_773),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_1699),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_482),
.Y(n_2682)
);

BUFx10_ASAP7_75t_L g2683 ( 
.A(n_1096),
.Y(n_2683)
);

CKINVDCx5p33_ASAP7_75t_R g2684 ( 
.A(n_1738),
.Y(n_2684)
);

CKINVDCx5p33_ASAP7_75t_R g2685 ( 
.A(n_360),
.Y(n_2685)
);

CKINVDCx5p33_ASAP7_75t_R g2686 ( 
.A(n_1118),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_1020),
.Y(n_2687)
);

BUFx2_ASAP7_75t_L g2688 ( 
.A(n_1772),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_1860),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_1631),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_1837),
.Y(n_2691)
);

CKINVDCx5p33_ASAP7_75t_R g2692 ( 
.A(n_1304),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_139),
.Y(n_2693)
);

BUFx6f_ASAP7_75t_L g2694 ( 
.A(n_1727),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_623),
.Y(n_2695)
);

INVx1_ASAP7_75t_SL g2696 ( 
.A(n_1765),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_1359),
.Y(n_2697)
);

INVxp67_ASAP7_75t_L g2698 ( 
.A(n_226),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_519),
.Y(n_2699)
);

CKINVDCx20_ASAP7_75t_R g2700 ( 
.A(n_1232),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_249),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_445),
.Y(n_2702)
);

BUFx10_ASAP7_75t_L g2703 ( 
.A(n_1644),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_735),
.Y(n_2704)
);

BUFx8_ASAP7_75t_SL g2705 ( 
.A(n_1625),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_1753),
.Y(n_2706)
);

BUFx2_ASAP7_75t_L g2707 ( 
.A(n_1691),
.Y(n_2707)
);

INVx2_ASAP7_75t_SL g2708 ( 
.A(n_1093),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_374),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_714),
.Y(n_2710)
);

BUFx6f_ASAP7_75t_L g2711 ( 
.A(n_1088),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_1061),
.Y(n_2712)
);

CKINVDCx5p33_ASAP7_75t_R g2713 ( 
.A(n_1639),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_1469),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_346),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_267),
.Y(n_2716)
);

CKINVDCx20_ASAP7_75t_R g2717 ( 
.A(n_384),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_1595),
.Y(n_2718)
);

CKINVDCx5p33_ASAP7_75t_R g2719 ( 
.A(n_788),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_247),
.Y(n_2720)
);

BUFx2_ASAP7_75t_L g2721 ( 
.A(n_1684),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_1049),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_1755),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_697),
.Y(n_2724)
);

CKINVDCx5p33_ASAP7_75t_R g2725 ( 
.A(n_195),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_986),
.Y(n_2726)
);

CKINVDCx20_ASAP7_75t_R g2727 ( 
.A(n_1450),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_1774),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_1740),
.Y(n_2729)
);

CKINVDCx20_ASAP7_75t_R g2730 ( 
.A(n_587),
.Y(n_2730)
);

CKINVDCx5p33_ASAP7_75t_R g2731 ( 
.A(n_899),
.Y(n_2731)
);

BUFx6f_ASAP7_75t_L g2732 ( 
.A(n_178),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_1137),
.Y(n_2733)
);

CKINVDCx5p33_ASAP7_75t_R g2734 ( 
.A(n_1506),
.Y(n_2734)
);

CKINVDCx5p33_ASAP7_75t_R g2735 ( 
.A(n_1651),
.Y(n_2735)
);

INVx1_ASAP7_75t_SL g2736 ( 
.A(n_1851),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_1592),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_1485),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_1239),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_1728),
.Y(n_2740)
);

CKINVDCx5p33_ASAP7_75t_R g2741 ( 
.A(n_1647),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_1572),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_188),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_1589),
.Y(n_2744)
);

CKINVDCx5p33_ASAP7_75t_R g2745 ( 
.A(n_1722),
.Y(n_2745)
);

BUFx8_ASAP7_75t_SL g2746 ( 
.A(n_424),
.Y(n_2746)
);

CKINVDCx5p33_ASAP7_75t_R g2747 ( 
.A(n_1429),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_384),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_781),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_1476),
.Y(n_2750)
);

BUFx3_ASAP7_75t_L g2751 ( 
.A(n_767),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_1642),
.Y(n_2752)
);

INVx1_ASAP7_75t_SL g2753 ( 
.A(n_1554),
.Y(n_2753)
);

BUFx2_ASAP7_75t_SL g2754 ( 
.A(n_201),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_1545),
.Y(n_2755)
);

CKINVDCx5p33_ASAP7_75t_R g2756 ( 
.A(n_1632),
.Y(n_2756)
);

CKINVDCx20_ASAP7_75t_R g2757 ( 
.A(n_1257),
.Y(n_2757)
);

CKINVDCx16_ASAP7_75t_R g2758 ( 
.A(n_415),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_1099),
.Y(n_2759)
);

CKINVDCx5p33_ASAP7_75t_R g2760 ( 
.A(n_1773),
.Y(n_2760)
);

CKINVDCx5p33_ASAP7_75t_R g2761 ( 
.A(n_955),
.Y(n_2761)
);

CKINVDCx5p33_ASAP7_75t_R g2762 ( 
.A(n_1643),
.Y(n_2762)
);

CKINVDCx5p33_ASAP7_75t_R g2763 ( 
.A(n_410),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_635),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_1733),
.Y(n_2765)
);

BUFx10_ASAP7_75t_L g2766 ( 
.A(n_511),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_1775),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_1418),
.Y(n_2768)
);

BUFx5_ASAP7_75t_L g2769 ( 
.A(n_1636),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_192),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_1560),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_404),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_1507),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_1030),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_1498),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_1878),
.Y(n_2776)
);

CKINVDCx5p33_ASAP7_75t_R g2777 ( 
.A(n_1393),
.Y(n_2777)
);

INVx1_ASAP7_75t_SL g2778 ( 
.A(n_1352),
.Y(n_2778)
);

CKINVDCx20_ASAP7_75t_R g2779 ( 
.A(n_950),
.Y(n_2779)
);

CKINVDCx5p33_ASAP7_75t_R g2780 ( 
.A(n_321),
.Y(n_2780)
);

CKINVDCx5p33_ASAP7_75t_R g2781 ( 
.A(n_1370),
.Y(n_2781)
);

CKINVDCx20_ASAP7_75t_R g2782 ( 
.A(n_1103),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_1219),
.Y(n_2783)
);

CKINVDCx5p33_ASAP7_75t_R g2784 ( 
.A(n_516),
.Y(n_2784)
);

CKINVDCx5p33_ASAP7_75t_R g2785 ( 
.A(n_107),
.Y(n_2785)
);

CKINVDCx5p33_ASAP7_75t_R g2786 ( 
.A(n_428),
.Y(n_2786)
);

CKINVDCx20_ASAP7_75t_R g2787 ( 
.A(n_1455),
.Y(n_2787)
);

CKINVDCx14_ASAP7_75t_R g2788 ( 
.A(n_1084),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_117),
.Y(n_2789)
);

CKINVDCx5p33_ASAP7_75t_R g2790 ( 
.A(n_1303),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_1460),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_1752),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_324),
.Y(n_2793)
);

CKINVDCx5p33_ASAP7_75t_R g2794 ( 
.A(n_500),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_493),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_769),
.Y(n_2796)
);

CKINVDCx5p33_ASAP7_75t_R g2797 ( 
.A(n_569),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_1844),
.Y(n_2798)
);

CKINVDCx5p33_ASAP7_75t_R g2799 ( 
.A(n_1548),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_999),
.Y(n_2800)
);

CKINVDCx20_ASAP7_75t_R g2801 ( 
.A(n_821),
.Y(n_2801)
);

HB1xp67_ASAP7_75t_L g2802 ( 
.A(n_1466),
.Y(n_2802)
);

CKINVDCx20_ASAP7_75t_R g2803 ( 
.A(n_1656),
.Y(n_2803)
);

CKINVDCx5p33_ASAP7_75t_R g2804 ( 
.A(n_1192),
.Y(n_2804)
);

CKINVDCx20_ASAP7_75t_R g2805 ( 
.A(n_1223),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_1329),
.Y(n_2806)
);

CKINVDCx5p33_ASAP7_75t_R g2807 ( 
.A(n_427),
.Y(n_2807)
);

CKINVDCx5p33_ASAP7_75t_R g2808 ( 
.A(n_1313),
.Y(n_2808)
);

CKINVDCx5p33_ASAP7_75t_R g2809 ( 
.A(n_1077),
.Y(n_2809)
);

CKINVDCx5p33_ASAP7_75t_R g2810 ( 
.A(n_638),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_200),
.Y(n_2811)
);

CKINVDCx5p33_ASAP7_75t_R g2812 ( 
.A(n_330),
.Y(n_2812)
);

CKINVDCx5p33_ASAP7_75t_R g2813 ( 
.A(n_1416),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_1669),
.Y(n_2814)
);

INVx2_ASAP7_75t_L g2815 ( 
.A(n_1586),
.Y(n_2815)
);

CKINVDCx14_ASAP7_75t_R g2816 ( 
.A(n_177),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_1147),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_1635),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_1646),
.Y(n_2819)
);

BUFx5_ASAP7_75t_L g2820 ( 
.A(n_1670),
.Y(n_2820)
);

CKINVDCx5p33_ASAP7_75t_R g2821 ( 
.A(n_508),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_1232),
.Y(n_2822)
);

CKINVDCx5p33_ASAP7_75t_R g2823 ( 
.A(n_600),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_932),
.Y(n_2824)
);

CKINVDCx5p33_ASAP7_75t_R g2825 ( 
.A(n_1619),
.Y(n_2825)
);

CKINVDCx20_ASAP7_75t_R g2826 ( 
.A(n_1653),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_506),
.Y(n_2827)
);

BUFx2_ASAP7_75t_L g2828 ( 
.A(n_1078),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_938),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_493),
.Y(n_2830)
);

INVxp67_ASAP7_75t_SL g2831 ( 
.A(n_1718),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_1441),
.Y(n_2832)
);

CKINVDCx20_ASAP7_75t_R g2833 ( 
.A(n_1402),
.Y(n_2833)
);

CKINVDCx5p33_ASAP7_75t_R g2834 ( 
.A(n_338),
.Y(n_2834)
);

BUFx6f_ASAP7_75t_L g2835 ( 
.A(n_382),
.Y(n_2835)
);

CKINVDCx5p33_ASAP7_75t_R g2836 ( 
.A(n_1369),
.Y(n_2836)
);

BUFx6f_ASAP7_75t_L g2837 ( 
.A(n_1295),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_956),
.Y(n_2838)
);

CKINVDCx20_ASAP7_75t_R g2839 ( 
.A(n_567),
.Y(n_2839)
);

CKINVDCx5p33_ASAP7_75t_R g2840 ( 
.A(n_1679),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_1876),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_184),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_1737),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_151),
.Y(n_2844)
);

CKINVDCx5p33_ASAP7_75t_R g2845 ( 
.A(n_1823),
.Y(n_2845)
);

CKINVDCx5p33_ASAP7_75t_R g2846 ( 
.A(n_1648),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_209),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_1484),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_1093),
.Y(n_2849)
);

BUFx3_ASAP7_75t_L g2850 ( 
.A(n_1827),
.Y(n_2850)
);

CKINVDCx5p33_ASAP7_75t_R g2851 ( 
.A(n_340),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_554),
.Y(n_2852)
);

CKINVDCx16_ASAP7_75t_R g2853 ( 
.A(n_1119),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_1724),
.Y(n_2854)
);

CKINVDCx5p33_ASAP7_75t_R g2855 ( 
.A(n_1573),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_1627),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_522),
.Y(n_2857)
);

CKINVDCx5p33_ASAP7_75t_R g2858 ( 
.A(n_1010),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_602),
.Y(n_2859)
);

INVx2_ASAP7_75t_SL g2860 ( 
.A(n_178),
.Y(n_2860)
);

CKINVDCx16_ASAP7_75t_R g2861 ( 
.A(n_1274),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_258),
.Y(n_2862)
);

BUFx10_ASAP7_75t_L g2863 ( 
.A(n_1732),
.Y(n_2863)
);

CKINVDCx20_ASAP7_75t_R g2864 ( 
.A(n_1229),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_929),
.Y(n_2865)
);

CKINVDCx5p33_ASAP7_75t_R g2866 ( 
.A(n_1695),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_1664),
.Y(n_2867)
);

CKINVDCx5p33_ASAP7_75t_R g2868 ( 
.A(n_325),
.Y(n_2868)
);

BUFx10_ASAP7_75t_L g2869 ( 
.A(n_993),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2184),
.B(n_0),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2476),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2476),
.Y(n_2872)
);

INVx1_ASAP7_75t_SL g2873 ( 
.A(n_1933),
.Y(n_2873)
);

INVxp67_ASAP7_75t_L g2874 ( 
.A(n_1896),
.Y(n_2874)
);

INVxp67_ASAP7_75t_SL g2875 ( 
.A(n_2564),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2564),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2617),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2617),
.Y(n_2878)
);

INVxp33_ASAP7_75t_L g2879 ( 
.A(n_1984),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2141),
.Y(n_2880)
);

CKINVDCx16_ASAP7_75t_R g2881 ( 
.A(n_2142),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2012),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2012),
.Y(n_2883)
);

INVxp67_ASAP7_75t_SL g2884 ( 
.A(n_1893),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2012),
.Y(n_2885)
);

CKINVDCx5p33_ASAP7_75t_R g2886 ( 
.A(n_2705),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2012),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_1902),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2012),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2231),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2231),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2231),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2231),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2231),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2315),
.Y(n_2895)
);

NOR2xp67_ASAP7_75t_L g2896 ( 
.A(n_2004),
.B(n_0),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2315),
.Y(n_2897)
);

CKINVDCx20_ASAP7_75t_R g2898 ( 
.A(n_2145),
.Y(n_2898)
);

CKINVDCx16_ASAP7_75t_R g2899 ( 
.A(n_2274),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2315),
.Y(n_2900)
);

CKINVDCx5p33_ASAP7_75t_R g2901 ( 
.A(n_2746),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2315),
.Y(n_2902)
);

CKINVDCx5p33_ASAP7_75t_R g2903 ( 
.A(n_2021),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2315),
.Y(n_2904)
);

BUFx2_ASAP7_75t_L g2905 ( 
.A(n_1964),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2417),
.Y(n_2906)
);

INVxp33_ASAP7_75t_SL g2907 ( 
.A(n_2198),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2417),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2417),
.Y(n_2909)
);

CKINVDCx5p33_ASAP7_75t_R g2910 ( 
.A(n_2100),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2417),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2417),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2769),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2769),
.Y(n_2914)
);

CKINVDCx5p33_ASAP7_75t_R g2915 ( 
.A(n_2206),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2769),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2769),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_2226),
.Y(n_2918)
);

BUFx6f_ASAP7_75t_L g2919 ( 
.A(n_1893),
.Y(n_2919)
);

CKINVDCx20_ASAP7_75t_R g2920 ( 
.A(n_2298),
.Y(n_2920)
);

INVxp67_ASAP7_75t_SL g2921 ( 
.A(n_1893),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2769),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2820),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2820),
.Y(n_2924)
);

CKINVDCx20_ASAP7_75t_R g2925 ( 
.A(n_2468),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2820),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2820),
.Y(n_2927)
);

INVxp67_ASAP7_75t_SL g2928 ( 
.A(n_1970),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2820),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_1970),
.Y(n_2930)
);

BUFx3_ASAP7_75t_L g2931 ( 
.A(n_1920),
.Y(n_2931)
);

HB1xp67_ASAP7_75t_L g2932 ( 
.A(n_2240),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_1884),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_1897),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_1903),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_1910),
.Y(n_2936)
);

INVxp67_ASAP7_75t_SL g2937 ( 
.A(n_1970),
.Y(n_2937)
);

CKINVDCx5p33_ASAP7_75t_R g2938 ( 
.A(n_2284),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_1917),
.Y(n_2939)
);

BUFx6f_ASAP7_75t_L g2940 ( 
.A(n_1979),
.Y(n_2940)
);

HB1xp67_ASAP7_75t_L g2941 ( 
.A(n_2337),
.Y(n_2941)
);

NOR2xp67_ASAP7_75t_L g2942 ( 
.A(n_2384),
.B(n_2),
.Y(n_2942)
);

CKINVDCx16_ASAP7_75t_R g2943 ( 
.A(n_2788),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_1925),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_1927),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_1928),
.Y(n_2946)
);

CKINVDCx16_ASAP7_75t_R g2947 ( 
.A(n_2816),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_1934),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_1940),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_1944),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_1951),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_1955),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_1956),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_1959),
.Y(n_2954)
);

INVx2_ASAP7_75t_SL g2955 ( 
.A(n_2869),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_1961),
.Y(n_2956)
);

INVxp67_ASAP7_75t_L g2957 ( 
.A(n_2055),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_1962),
.Y(n_2958)
);

CKINVDCx5p33_ASAP7_75t_R g2959 ( 
.A(n_2424),
.Y(n_2959)
);

INVxp33_ASAP7_75t_L g2960 ( 
.A(n_2481),
.Y(n_2960)
);

OR2x2_ASAP7_75t_L g2961 ( 
.A(n_2154),
.B(n_2),
.Y(n_2961)
);

CKINVDCx5p33_ASAP7_75t_R g2962 ( 
.A(n_2530),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_1966),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_1971),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_1978),
.Y(n_2965)
);

CKINVDCx14_ASAP7_75t_R g2966 ( 
.A(n_2412),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_1991),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2000),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2001),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2008),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2009),
.Y(n_2971)
);

CKINVDCx20_ASAP7_75t_R g2972 ( 
.A(n_2493),
.Y(n_2972)
);

INVx2_ASAP7_75t_L g2973 ( 
.A(n_1979),
.Y(n_2973)
);

CKINVDCx5p33_ASAP7_75t_R g2974 ( 
.A(n_2565),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2010),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2018),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2026),
.Y(n_2977)
);

INVxp33_ASAP7_75t_SL g2978 ( 
.A(n_2673),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2029),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2030),
.Y(n_2980)
);

CKINVDCx20_ASAP7_75t_R g2981 ( 
.A(n_2534),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2032),
.Y(n_2982)
);

CKINVDCx5p33_ASAP7_75t_R g2983 ( 
.A(n_2594),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2035),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_1979),
.Y(n_2985)
);

CKINVDCx5p33_ASAP7_75t_R g2986 ( 
.A(n_2621),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2039),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2040),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2042),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2051),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2053),
.Y(n_2991)
);

INVxp33_ASAP7_75t_SL g2992 ( 
.A(n_2677),
.Y(n_2992)
);

INVx1_ASAP7_75t_L g2993 ( 
.A(n_2054),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2057),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2066),
.Y(n_2995)
);

INVxp67_ASAP7_75t_SL g2996 ( 
.A(n_1988),
.Y(n_2996)
);

CKINVDCx20_ASAP7_75t_R g2997 ( 
.A(n_2864),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_1988),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2068),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_1921),
.Y(n_3000)
);

CKINVDCx5p33_ASAP7_75t_R g3001 ( 
.A(n_2758),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2070),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2071),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2072),
.Y(n_3004)
);

CKINVDCx5p33_ASAP7_75t_R g3005 ( 
.A(n_2853),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_1988),
.Y(n_3006)
);

CKINVDCx20_ASAP7_75t_R g3007 ( 
.A(n_1932),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2078),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2090),
.Y(n_3009)
);

INVx2_ASAP7_75t_L g3010 ( 
.A(n_2249),
.Y(n_3010)
);

XNOR2xp5_ASAP7_75t_L g3011 ( 
.A(n_1938),
.B(n_3),
.Y(n_3011)
);

INVxp33_ASAP7_75t_SL g3012 ( 
.A(n_2774),
.Y(n_3012)
);

INVx1_ASAP7_75t_L g3013 ( 
.A(n_2101),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2103),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2106),
.Y(n_3015)
);

INVxp33_ASAP7_75t_SL g3016 ( 
.A(n_2802),
.Y(n_3016)
);

INVxp67_ASAP7_75t_SL g3017 ( 
.A(n_2249),
.Y(n_3017)
);

INVxp67_ASAP7_75t_SL g3018 ( 
.A(n_2249),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2107),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2114),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2122),
.Y(n_3021)
);

BUFx2_ASAP7_75t_L g3022 ( 
.A(n_2168),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2252),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2130),
.Y(n_3024)
);

INVxp33_ASAP7_75t_SL g3025 ( 
.A(n_2843),
.Y(n_3025)
);

CKINVDCx20_ASAP7_75t_R g3026 ( 
.A(n_1943),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2132),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2133),
.Y(n_3028)
);

NOR2xp67_ASAP7_75t_L g3029 ( 
.A(n_1942),
.B(n_3),
.Y(n_3029)
);

INVx1_ASAP7_75t_SL g3030 ( 
.A(n_1950),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2135),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2138),
.Y(n_3032)
);

CKINVDCx5p33_ASAP7_75t_R g3033 ( 
.A(n_2861),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2143),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2144),
.Y(n_3035)
);

CKINVDCx5p33_ASAP7_75t_R g3036 ( 
.A(n_2856),
.Y(n_3036)
);

CKINVDCx20_ASAP7_75t_R g3037 ( 
.A(n_1963),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2146),
.Y(n_3038)
);

BUFx3_ASAP7_75t_L g3039 ( 
.A(n_1987),
.Y(n_3039)
);

CKINVDCx16_ASAP7_75t_R g3040 ( 
.A(n_1906),
.Y(n_3040)
);

BUFx2_ASAP7_75t_L g3041 ( 
.A(n_2209),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2150),
.Y(n_3042)
);

INVxp33_ASAP7_75t_L g3043 ( 
.A(n_2212),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2152),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2153),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2175),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2176),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2178),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_1883),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2189),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2193),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2195),
.Y(n_3052)
);

HB1xp67_ASAP7_75t_L g3053 ( 
.A(n_2214),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2202),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2203),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2208),
.Y(n_3056)
);

INVxp33_ASAP7_75t_L g3057 ( 
.A(n_2308),
.Y(n_3057)
);

INVxp67_ASAP7_75t_L g3058 ( 
.A(n_2340),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2215),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2217),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2219),
.Y(n_3061)
);

INVxp33_ASAP7_75t_L g3062 ( 
.A(n_2556),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2227),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2234),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2243),
.Y(n_3065)
);

HB1xp67_ASAP7_75t_L g3066 ( 
.A(n_2592),
.Y(n_3066)
);

HB1xp67_ASAP7_75t_SL g3067 ( 
.A(n_2229),
.Y(n_3067)
);

CKINVDCx5p33_ASAP7_75t_R g3068 ( 
.A(n_2855),
.Y(n_3068)
);

INVx1_ASAP7_75t_SL g3069 ( 
.A(n_1965),
.Y(n_3069)
);

INVxp33_ASAP7_75t_SL g3070 ( 
.A(n_2688),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2250),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2254),
.Y(n_3072)
);

CKINVDCx20_ASAP7_75t_R g3073 ( 
.A(n_1973),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2255),
.Y(n_3074)
);

CKINVDCx20_ASAP7_75t_R g3075 ( 
.A(n_1983),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2256),
.Y(n_3076)
);

BUFx6f_ASAP7_75t_L g3077 ( 
.A(n_2252),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2259),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2261),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2269),
.Y(n_3080)
);

BUFx3_ASAP7_75t_L g3081 ( 
.A(n_2020),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2252),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2283),
.Y(n_3083)
);

BUFx3_ASAP7_75t_L g3084 ( 
.A(n_2160),
.Y(n_3084)
);

INVx1_ASAP7_75t_L g3085 ( 
.A(n_2297),
.Y(n_3085)
);

CKINVDCx5p33_ASAP7_75t_R g3086 ( 
.A(n_2858),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2303),
.Y(n_3087)
);

INVxp33_ASAP7_75t_SL g3088 ( 
.A(n_2707),
.Y(n_3088)
);

INVxp33_ASAP7_75t_L g3089 ( 
.A(n_2721),
.Y(n_3089)
);

OR2x2_ASAP7_75t_L g3090 ( 
.A(n_2828),
.B(n_4),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2875),
.B(n_2080),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2884),
.B(n_2097),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2919),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2955),
.B(n_2222),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_2881),
.B(n_2304),
.Y(n_3095)
);

BUFx12f_ASAP7_75t_L g3096 ( 
.A(n_2886),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_2919),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2921),
.B(n_2691),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2928),
.Y(n_3099)
);

INVx4_ASAP7_75t_L g3100 ( 
.A(n_3036),
.Y(n_3100)
);

NOR2x1_ASAP7_75t_L g3101 ( 
.A(n_2931),
.B(n_2294),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2899),
.B(n_2776),
.Y(n_3102)
);

INVx5_ASAP7_75t_L g3103 ( 
.A(n_3040),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2937),
.B(n_2798),
.Y(n_3104)
);

BUFx6f_ASAP7_75t_L g3105 ( 
.A(n_2919),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2943),
.B(n_2402),
.Y(n_3106)
);

INVx5_ASAP7_75t_L g3107 ( 
.A(n_2905),
.Y(n_3107)
);

INVx5_ASAP7_75t_L g3108 ( 
.A(n_3022),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2996),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3017),
.B(n_1912),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_3018),
.B(n_2074),
.Y(n_3111)
);

OR2x2_ASAP7_75t_L g3112 ( 
.A(n_3041),
.B(n_2305),
.Y(n_3112)
);

INVx3_ASAP7_75t_L g3113 ( 
.A(n_3000),
.Y(n_3113)
);

NOR2xp33_ASAP7_75t_L g3114 ( 
.A(n_2947),
.B(n_2736),
.Y(n_3114)
);

BUFx12f_ASAP7_75t_L g3115 ( 
.A(n_2901),
.Y(n_3115)
);

NOR2xp33_ASAP7_75t_L g3116 ( 
.A(n_3049),
.B(n_2609),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2940),
.Y(n_3117)
);

INVx5_ASAP7_75t_L g3118 ( 
.A(n_2940),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_3039),
.Y(n_3119)
);

HB1xp67_ASAP7_75t_L g3120 ( 
.A(n_2903),
.Y(n_3120)
);

INVx5_ASAP7_75t_L g3121 ( 
.A(n_2940),
.Y(n_3121)
);

INVx4_ASAP7_75t_L g3122 ( 
.A(n_3068),
.Y(n_3122)
);

BUFx2_ASAP7_75t_L g3123 ( 
.A(n_2910),
.Y(n_3123)
);

BUFx6f_ASAP7_75t_L g3124 ( 
.A(n_3077),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_3077),
.Y(n_3125)
);

BUFx12f_ASAP7_75t_L g3126 ( 
.A(n_2915),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2882),
.B(n_2689),
.Y(n_3127)
);

AND2x4_ASAP7_75t_L g3128 ( 
.A(n_2874),
.B(n_2244),
.Y(n_3128)
);

BUFx6f_ASAP7_75t_L g3129 ( 
.A(n_3077),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_3043),
.B(n_3057),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2871),
.Y(n_3131)
);

INVx4_ASAP7_75t_L g3132 ( 
.A(n_3086),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2872),
.Y(n_3133)
);

BUFx8_ASAP7_75t_SL g3134 ( 
.A(n_2997),
.Y(n_3134)
);

AND2x4_ASAP7_75t_L g3135 ( 
.A(n_2888),
.B(n_2280),
.Y(n_3135)
);

AND2x2_ASAP7_75t_L g3136 ( 
.A(n_3062),
.B(n_1906),
.Y(n_3136)
);

BUFx3_ASAP7_75t_L g3137 ( 
.A(n_3081),
.Y(n_3137)
);

BUFx3_ASAP7_75t_L g3138 ( 
.A(n_3084),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2883),
.B(n_2841),
.Y(n_3139)
);

BUFx6f_ASAP7_75t_L g3140 ( 
.A(n_2930),
.Y(n_3140)
);

INVx5_ASAP7_75t_L g3141 ( 
.A(n_2973),
.Y(n_3141)
);

NOR2x1_ASAP7_75t_L g3142 ( 
.A(n_2876),
.B(n_2877),
.Y(n_3142)
);

HB1xp67_ASAP7_75t_L g3143 ( 
.A(n_2918),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_L g3144 ( 
.A(n_3070),
.B(n_1937),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2878),
.Y(n_3145)
);

BUFx6f_ASAP7_75t_L g3146 ( 
.A(n_2985),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_3088),
.B(n_1941),
.Y(n_3147)
);

BUFx12f_ASAP7_75t_L g3148 ( 
.A(n_2938),
.Y(n_3148)
);

BUFx12f_ASAP7_75t_L g3149 ( 
.A(n_2959),
.Y(n_3149)
);

AND2x4_ASAP7_75t_L g3150 ( 
.A(n_2957),
.B(n_2288),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2885),
.B(n_2887),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2889),
.B(n_1996),
.Y(n_3152)
);

NOR2xp33_ASAP7_75t_L g3153 ( 
.A(n_2907),
.B(n_2061),
.Y(n_3153)
);

BUFx2_ASAP7_75t_L g3154 ( 
.A(n_2962),
.Y(n_3154)
);

BUFx6f_ASAP7_75t_L g3155 ( 
.A(n_2998),
.Y(n_3155)
);

AND2x6_ASAP7_75t_L g3156 ( 
.A(n_2873),
.B(n_2382),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_2933),
.B(n_2464),
.Y(n_3157)
);

BUFx6f_ASAP7_75t_L g3158 ( 
.A(n_3006),
.Y(n_3158)
);

AND2x4_ASAP7_75t_L g3159 ( 
.A(n_3058),
.B(n_2472),
.Y(n_3159)
);

AND2x4_ASAP7_75t_L g3160 ( 
.A(n_3053),
.B(n_2485),
.Y(n_3160)
);

BUFx12f_ASAP7_75t_L g3161 ( 
.A(n_2974),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_3010),
.Y(n_3162)
);

AND2x4_ASAP7_75t_L g3163 ( 
.A(n_3066),
.B(n_2540),
.Y(n_3163)
);

INVx4_ASAP7_75t_L g3164 ( 
.A(n_2983),
.Y(n_3164)
);

AND2x4_ASAP7_75t_L g3165 ( 
.A(n_2932),
.B(n_2597),
.Y(n_3165)
);

NAND2xp5_ASAP7_75t_L g3166 ( 
.A(n_2890),
.B(n_2126),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_3023),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_3082),
.Y(n_3168)
);

BUFx6f_ASAP7_75t_L g3169 ( 
.A(n_2934),
.Y(n_3169)
);

NOR2xp33_ASAP7_75t_SL g3170 ( 
.A(n_2880),
.B(n_2007),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2891),
.B(n_2892),
.Y(n_3171)
);

INVx2_ASAP7_75t_SL g3172 ( 
.A(n_2986),
.Y(n_3172)
);

BUFx3_ASAP7_75t_L g3173 ( 
.A(n_2893),
.Y(n_3173)
);

BUFx12f_ASAP7_75t_L g3174 ( 
.A(n_3001),
.Y(n_3174)
);

BUFx6f_ASAP7_75t_L g3175 ( 
.A(n_2935),
.Y(n_3175)
);

BUFx12f_ASAP7_75t_L g3176 ( 
.A(n_3005),
.Y(n_3176)
);

INVx5_ASAP7_75t_L g3177 ( 
.A(n_3067),
.Y(n_3177)
);

BUFx6f_ASAP7_75t_L g3178 ( 
.A(n_2936),
.Y(n_3178)
);

BUFx6f_ASAP7_75t_L g3179 ( 
.A(n_2939),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2894),
.Y(n_3180)
);

NAND2xp5_ASAP7_75t_L g3181 ( 
.A(n_2895),
.B(n_2190),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2897),
.Y(n_3182)
);

AND2x4_ASAP7_75t_L g3183 ( 
.A(n_2941),
.B(n_2643),
.Y(n_3183)
);

INVx5_ASAP7_75t_L g3184 ( 
.A(n_2978),
.Y(n_3184)
);

NOR2xp33_ASAP7_75t_L g3185 ( 
.A(n_2992),
.B(n_2258),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2900),
.Y(n_3186)
);

BUFx6f_ASAP7_75t_L g3187 ( 
.A(n_2944),
.Y(n_3187)
);

NOR2xp33_ASAP7_75t_L g3188 ( 
.A(n_3012),
.B(n_2323),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_3033),
.Y(n_3189)
);

INVx3_ASAP7_75t_L g3190 ( 
.A(n_2945),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2902),
.Y(n_3191)
);

BUFx6f_ASAP7_75t_L g3192 ( 
.A(n_2946),
.Y(n_3192)
);

INVx2_ASAP7_75t_SL g3193 ( 
.A(n_3030),
.Y(n_3193)
);

HB1xp67_ASAP7_75t_L g3194 ( 
.A(n_3069),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2904),
.Y(n_3195)
);

BUFx2_ASAP7_75t_L g3196 ( 
.A(n_2898),
.Y(n_3196)
);

INVx5_ASAP7_75t_L g3197 ( 
.A(n_3016),
.Y(n_3197)
);

AND2x2_ASAP7_75t_L g3198 ( 
.A(n_3089),
.B(n_1945),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2906),
.Y(n_3199)
);

BUFx6f_ASAP7_75t_L g3200 ( 
.A(n_2948),
.Y(n_3200)
);

INVx5_ASAP7_75t_L g3201 ( 
.A(n_3025),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2908),
.Y(n_3202)
);

AND2x4_ASAP7_75t_L g3203 ( 
.A(n_2920),
.B(n_2751),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_2925),
.B(n_2850),
.Y(n_3204)
);

INVx5_ASAP7_75t_L g3205 ( 
.A(n_2879),
.Y(n_3205)
);

BUFx6f_ASAP7_75t_L g3206 ( 
.A(n_2949),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2909),
.B(n_2521),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2960),
.B(n_1945),
.Y(n_3208)
);

NOR2xp33_ASAP7_75t_L g3209 ( 
.A(n_2911),
.B(n_2576),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2912),
.B(n_2631),
.Y(n_3210)
);

AND2x4_ASAP7_75t_L g3211 ( 
.A(n_2950),
.B(n_1930),
.Y(n_3211)
);

BUFx6f_ASAP7_75t_L g3212 ( 
.A(n_2951),
.Y(n_3212)
);

BUFx12f_ASAP7_75t_L g3213 ( 
.A(n_2961),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2913),
.B(n_1990),
.Y(n_3214)
);

NOR2xp33_ASAP7_75t_L g3215 ( 
.A(n_2914),
.B(n_2361),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2952),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_2953),
.B(n_1935),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2916),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2917),
.Y(n_3219)
);

AND2x4_ASAP7_75t_L g3220 ( 
.A(n_2954),
.B(n_1939),
.Y(n_3220)
);

INVx3_ASAP7_75t_L g3221 ( 
.A(n_2956),
.Y(n_3221)
);

AND2x4_ASAP7_75t_L g3222 ( 
.A(n_2958),
.B(n_2081),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2963),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2922),
.Y(n_3224)
);

AND2x6_ASAP7_75t_L g3225 ( 
.A(n_2964),
.B(n_2332),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_2966),
.B(n_1957),
.Y(n_3226)
);

AND2x4_ASAP7_75t_L g3227 ( 
.A(n_2965),
.B(n_2086),
.Y(n_3227)
);

INVx4_ASAP7_75t_L g3228 ( 
.A(n_3090),
.Y(n_3228)
);

CKINVDCx5p33_ASAP7_75t_R g3229 ( 
.A(n_2972),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2923),
.B(n_2430),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_2924),
.B(n_2452),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_2926),
.B(n_2455),
.Y(n_3232)
);

BUFx12f_ASAP7_75t_L g3233 ( 
.A(n_2981),
.Y(n_3233)
);

BUFx8_ASAP7_75t_SL g3234 ( 
.A(n_3007),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_2967),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2927),
.Y(n_3236)
);

INVx5_ASAP7_75t_L g3237 ( 
.A(n_2896),
.Y(n_3237)
);

AND2x4_ASAP7_75t_L g3238 ( 
.A(n_2968),
.B(n_2636),
.Y(n_3238)
);

BUFx6f_ASAP7_75t_L g3239 ( 
.A(n_2969),
.Y(n_3239)
);

INVx3_ASAP7_75t_L g3240 ( 
.A(n_2970),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_2929),
.B(n_2644),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2971),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2975),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2976),
.B(n_2708),
.Y(n_3244)
);

BUFx2_ASAP7_75t_L g3245 ( 
.A(n_3026),
.Y(n_3245)
);

NAND2xp33_ASAP7_75t_L g3246 ( 
.A(n_2977),
.B(n_2332),
.Y(n_3246)
);

INVx6_ASAP7_75t_L g3247 ( 
.A(n_2942),
.Y(n_3247)
);

BUFx12f_ASAP7_75t_L g3248 ( 
.A(n_3037),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_3087),
.B(n_2698),
.Y(n_3249)
);

BUFx6f_ASAP7_75t_L g3250 ( 
.A(n_2979),
.Y(n_3250)
);

BUFx6f_ASAP7_75t_L g3251 ( 
.A(n_2980),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2982),
.B(n_2860),
.Y(n_3252)
);

BUFx6f_ASAP7_75t_L g3253 ( 
.A(n_2984),
.Y(n_3253)
);

AND2x2_ASAP7_75t_L g3254 ( 
.A(n_2987),
.B(n_1957),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_L g3255 ( 
.A(n_2988),
.B(n_2867),
.Y(n_3255)
);

INVx5_ASAP7_75t_L g3256 ( 
.A(n_3073),
.Y(n_3256)
);

BUFx8_ASAP7_75t_SL g3257 ( 
.A(n_3075),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_2989),
.B(n_1885),
.Y(n_3258)
);

INVx3_ASAP7_75t_L g3259 ( 
.A(n_2990),
.Y(n_3259)
);

INVx4_ASAP7_75t_L g3260 ( 
.A(n_2991),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2993),
.Y(n_3261)
);

AND2x2_ASAP7_75t_L g3262 ( 
.A(n_2994),
.B(n_1976),
.Y(n_3262)
);

AND2x2_ASAP7_75t_L g3263 ( 
.A(n_2995),
.B(n_1976),
.Y(n_3263)
);

BUFx12f_ASAP7_75t_L g3264 ( 
.A(n_3011),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2999),
.B(n_2332),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3002),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3003),
.B(n_2352),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3004),
.B(n_2352),
.Y(n_3268)
);

BUFx8_ASAP7_75t_SL g3269 ( 
.A(n_3085),
.Y(n_3269)
);

BUFx8_ASAP7_75t_SL g3270 ( 
.A(n_3008),
.Y(n_3270)
);

INVx3_ASAP7_75t_L g3271 ( 
.A(n_3009),
.Y(n_3271)
);

NOR2xp33_ASAP7_75t_L g3272 ( 
.A(n_3013),
.B(n_1886),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3014),
.Y(n_3273)
);

CKINVDCx6p67_ASAP7_75t_R g3274 ( 
.A(n_3015),
.Y(n_3274)
);

BUFx3_ASAP7_75t_L g3275 ( 
.A(n_3019),
.Y(n_3275)
);

BUFx3_ASAP7_75t_L g3276 ( 
.A(n_3020),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_3083),
.B(n_1887),
.Y(n_3277)
);

AND2x6_ASAP7_75t_L g3278 ( 
.A(n_3021),
.B(n_2352),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_3024),
.B(n_2409),
.Y(n_3279)
);

BUFx8_ASAP7_75t_L g3280 ( 
.A(n_3027),
.Y(n_3280)
);

NOR2xp33_ASAP7_75t_L g3281 ( 
.A(n_3080),
.B(n_1888),
.Y(n_3281)
);

INVx3_ASAP7_75t_L g3282 ( 
.A(n_3028),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_3079),
.B(n_1889),
.Y(n_3283)
);

AND2x4_ASAP7_75t_L g3284 ( 
.A(n_3031),
.B(n_1911),
.Y(n_3284)
);

BUFx6f_ASAP7_75t_L g3285 ( 
.A(n_3032),
.Y(n_3285)
);

BUFx6f_ASAP7_75t_L g3286 ( 
.A(n_3034),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3035),
.B(n_2409),
.Y(n_3287)
);

BUFx8_ASAP7_75t_L g3288 ( 
.A(n_3038),
.Y(n_3288)
);

BUFx12f_ASAP7_75t_L g3289 ( 
.A(n_2870),
.Y(n_3289)
);

NOR2xp33_ASAP7_75t_SL g3290 ( 
.A(n_3029),
.B(n_2031),
.Y(n_3290)
);

INVx2_ASAP7_75t_SL g3291 ( 
.A(n_3042),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3044),
.B(n_2409),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3045),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3046),
.B(n_2416),
.Y(n_3294)
);

INVx5_ASAP7_75t_L g3295 ( 
.A(n_3047),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3048),
.B(n_2017),
.Y(n_3296)
);

BUFx12f_ASAP7_75t_L g3297 ( 
.A(n_3050),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_3051),
.B(n_1890),
.Y(n_3298)
);

INVx4_ASAP7_75t_L g3299 ( 
.A(n_3052),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3054),
.B(n_2416),
.Y(n_3300)
);

BUFx12f_ASAP7_75t_L g3301 ( 
.A(n_3055),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3056),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_L g3303 ( 
.A(n_3059),
.B(n_2416),
.Y(n_3303)
);

BUFx8_ASAP7_75t_SL g3304 ( 
.A(n_3060),
.Y(n_3304)
);

NOR2xp33_ASAP7_75t_L g3305 ( 
.A(n_3078),
.B(n_1891),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3061),
.B(n_2457),
.Y(n_3306)
);

INVx5_ASAP7_75t_L g3307 ( 
.A(n_3063),
.Y(n_3307)
);

XOR2x2_ASAP7_75t_L g3308 ( 
.A(n_3064),
.B(n_1922),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3065),
.B(n_2457),
.Y(n_3309)
);

INVx4_ASAP7_75t_L g3310 ( 
.A(n_3071),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3072),
.B(n_2457),
.Y(n_3311)
);

AND2x2_ASAP7_75t_L g3312 ( 
.A(n_3074),
.B(n_2017),
.Y(n_3312)
);

NOR2xp33_ASAP7_75t_L g3313 ( 
.A(n_3076),
.B(n_1892),
.Y(n_3313)
);

BUFx8_ASAP7_75t_L g3314 ( 
.A(n_2905),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_2919),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_2875),
.B(n_1894),
.Y(n_3316)
);

INVx5_ASAP7_75t_L g3317 ( 
.A(n_3040),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2875),
.B(n_2602),
.Y(n_3318)
);

NOR2xp33_ASAP7_75t_L g3319 ( 
.A(n_2875),
.B(n_1895),
.Y(n_3319)
);

AND2x4_ASAP7_75t_L g3320 ( 
.A(n_2955),
.B(n_1958),
.Y(n_3320)
);

INVx5_ASAP7_75t_L g3321 ( 
.A(n_3040),
.Y(n_3321)
);

CKINVDCx5p33_ASAP7_75t_R g3322 ( 
.A(n_2966),
.Y(n_3322)
);

NOR2xp33_ASAP7_75t_L g3323 ( 
.A(n_2875),
.B(n_1898),
.Y(n_3323)
);

HB1xp67_ASAP7_75t_L g3324 ( 
.A(n_2903),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_2881),
.B(n_2059),
.Y(n_3325)
);

INVx5_ASAP7_75t_L g3326 ( 
.A(n_3040),
.Y(n_3326)
);

BUFx6f_ASAP7_75t_L g3327 ( 
.A(n_2919),
.Y(n_3327)
);

INVx5_ASAP7_75t_L g3328 ( 
.A(n_3040),
.Y(n_3328)
);

INVx3_ASAP7_75t_L g3329 ( 
.A(n_2931),
.Y(n_3329)
);

INVx1_ASAP7_75t_L g3330 ( 
.A(n_2884),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_2881),
.B(n_2059),
.Y(n_3331)
);

INVx2_ASAP7_75t_L g3332 ( 
.A(n_2919),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2875),
.B(n_2602),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_2919),
.Y(n_3334)
);

BUFx2_ASAP7_75t_L g3335 ( 
.A(n_2903),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_2875),
.B(n_2602),
.Y(n_3336)
);

AND2x4_ASAP7_75t_L g3337 ( 
.A(n_2955),
.B(n_1967),
.Y(n_3337)
);

INVx2_ASAP7_75t_L g3338 ( 
.A(n_2919),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2884),
.Y(n_3339)
);

BUFx12f_ASAP7_75t_L g3340 ( 
.A(n_2886),
.Y(n_3340)
);

CKINVDCx6p67_ASAP7_75t_R g3341 ( 
.A(n_2881),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2875),
.B(n_2648),
.Y(n_3342)
);

BUFx6f_ASAP7_75t_L g3343 ( 
.A(n_2919),
.Y(n_3343)
);

INVx2_ASAP7_75t_L g3344 ( 
.A(n_2919),
.Y(n_3344)
);

AND2x4_ASAP7_75t_L g3345 ( 
.A(n_2955),
.B(n_1972),
.Y(n_3345)
);

BUFx6f_ASAP7_75t_L g3346 ( 
.A(n_2919),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_2884),
.Y(n_3347)
);

INVx5_ASAP7_75t_L g3348 ( 
.A(n_3040),
.Y(n_3348)
);

INVx3_ASAP7_75t_L g3349 ( 
.A(n_2931),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_2881),
.B(n_2164),
.Y(n_3350)
);

AND2x4_ASAP7_75t_L g3351 ( 
.A(n_2955),
.B(n_2022),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_2875),
.B(n_1899),
.Y(n_3352)
);

INVx2_ASAP7_75t_L g3353 ( 
.A(n_2919),
.Y(n_3353)
);

INVx5_ASAP7_75t_L g3354 ( 
.A(n_3040),
.Y(n_3354)
);

INVx4_ASAP7_75t_L g3355 ( 
.A(n_3036),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_2881),
.B(n_2164),
.Y(n_3356)
);

INVx2_ASAP7_75t_SL g3357 ( 
.A(n_3036),
.Y(n_3357)
);

CKINVDCx20_ASAP7_75t_R g3358 ( 
.A(n_2997),
.Y(n_3358)
);

HB1xp67_ASAP7_75t_L g3359 ( 
.A(n_2903),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2919),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2875),
.B(n_2648),
.Y(n_3361)
);

CKINVDCx5p33_ASAP7_75t_R g3362 ( 
.A(n_2966),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_2875),
.B(n_2648),
.Y(n_3363)
);

CKINVDCx5p33_ASAP7_75t_R g3364 ( 
.A(n_2966),
.Y(n_3364)
);

BUFx3_ASAP7_75t_L g3365 ( 
.A(n_2931),
.Y(n_3365)
);

BUFx12f_ASAP7_75t_L g3366 ( 
.A(n_2886),
.Y(n_3366)
);

BUFx12f_ASAP7_75t_L g3367 ( 
.A(n_2886),
.Y(n_3367)
);

AND2x2_ASAP7_75t_L g3368 ( 
.A(n_2881),
.B(n_2220),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2875),
.B(n_1900),
.Y(n_3369)
);

CKINVDCx5p33_ASAP7_75t_R g3370 ( 
.A(n_2966),
.Y(n_3370)
);

AND2x4_ASAP7_75t_L g3371 ( 
.A(n_2955),
.B(n_2023),
.Y(n_3371)
);

INVxp33_ASAP7_75t_SL g3372 ( 
.A(n_2886),
.Y(n_3372)
);

AND2x4_ASAP7_75t_L g3373 ( 
.A(n_2955),
.B(n_2033),
.Y(n_3373)
);

HB1xp67_ASAP7_75t_L g3374 ( 
.A(n_2903),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_2955),
.B(n_2038),
.Y(n_3375)
);

BUFx12f_ASAP7_75t_L g3376 ( 
.A(n_2886),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_2955),
.B(n_2069),
.Y(n_3377)
);

BUFx6f_ASAP7_75t_L g3378 ( 
.A(n_2919),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2884),
.Y(n_3379)
);

INVx3_ASAP7_75t_L g3380 ( 
.A(n_2931),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2884),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_2875),
.B(n_2666),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2884),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_2881),
.B(n_2220),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2875),
.B(n_2666),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_2875),
.B(n_2666),
.Y(n_3386)
);

BUFx6f_ASAP7_75t_L g3387 ( 
.A(n_2919),
.Y(n_3387)
);

BUFx12f_ASAP7_75t_L g3388 ( 
.A(n_2886),
.Y(n_3388)
);

INVxp67_ASAP7_75t_L g3389 ( 
.A(n_3067),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_2875),
.B(n_2694),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_2884),
.Y(n_3391)
);

BUFx3_ASAP7_75t_L g3392 ( 
.A(n_2931),
.Y(n_3392)
);

AND2x4_ASAP7_75t_L g3393 ( 
.A(n_2955),
.B(n_2099),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_2881),
.B(n_2257),
.Y(n_3394)
);

BUFx8_ASAP7_75t_SL g3395 ( 
.A(n_2997),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_2884),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_2884),
.Y(n_3397)
);

BUFx6f_ASAP7_75t_L g3398 ( 
.A(n_2919),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_L g3399 ( 
.A(n_2875),
.B(n_1901),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_2881),
.B(n_2257),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_2875),
.B(n_2694),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2875),
.B(n_2694),
.Y(n_3402)
);

HB1xp67_ASAP7_75t_L g3403 ( 
.A(n_2903),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2919),
.Y(n_3404)
);

BUFx2_ASAP7_75t_L g3405 ( 
.A(n_2903),
.Y(n_3405)
);

BUFx2_ASAP7_75t_L g3406 ( 
.A(n_2903),
.Y(n_3406)
);

BUFx6f_ASAP7_75t_L g3407 ( 
.A(n_2919),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_2919),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2875),
.B(n_2711),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_2881),
.B(n_2327),
.Y(n_3410)
);

INVx4_ASAP7_75t_L g3411 ( 
.A(n_3036),
.Y(n_3411)
);

AND2x2_ASAP7_75t_SL g3412 ( 
.A(n_2881),
.B(n_2151),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2884),
.Y(n_3413)
);

INVx4_ASAP7_75t_L g3414 ( 
.A(n_3036),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_2919),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_L g3416 ( 
.A(n_2875),
.B(n_2711),
.Y(n_3416)
);

INVx5_ASAP7_75t_L g3417 ( 
.A(n_3040),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_SL g3418 ( 
.A(n_2881),
.B(n_2711),
.Y(n_3418)
);

AND2x4_ASAP7_75t_L g3419 ( 
.A(n_2955),
.B(n_2174),
.Y(n_3419)
);

INVx2_ASAP7_75t_SL g3420 ( 
.A(n_3036),
.Y(n_3420)
);

AND2x4_ASAP7_75t_L g3421 ( 
.A(n_2955),
.B(n_2265),
.Y(n_3421)
);

AND2x4_ASAP7_75t_L g3422 ( 
.A(n_2955),
.B(n_2277),
.Y(n_3422)
);

BUFx3_ASAP7_75t_L g3423 ( 
.A(n_2931),
.Y(n_3423)
);

AND2x4_ASAP7_75t_L g3424 ( 
.A(n_2955),
.B(n_2292),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_2875),
.B(n_2732),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_2881),
.B(n_2327),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_2881),
.B(n_2732),
.Y(n_3427)
);

HB1xp67_ASAP7_75t_L g3428 ( 
.A(n_2903),
.Y(n_3428)
);

AND2x2_ASAP7_75t_L g3429 ( 
.A(n_2881),
.B(n_2330),
.Y(n_3429)
);

HB1xp67_ASAP7_75t_L g3430 ( 
.A(n_2903),
.Y(n_3430)
);

AND2x4_ASAP7_75t_L g3431 ( 
.A(n_2955),
.B(n_2344),
.Y(n_3431)
);

AND2x4_ASAP7_75t_L g3432 ( 
.A(n_2955),
.B(n_2354),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_2875),
.B(n_2732),
.Y(n_3433)
);

AND2x4_ASAP7_75t_L g3434 ( 
.A(n_2955),
.B(n_2386),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3180),
.B(n_2829),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3131),
.Y(n_3436)
);

AND2x4_ASAP7_75t_L g3437 ( 
.A(n_3130),
.B(n_2034),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3140),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3133),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3145),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3242),
.Y(n_3441)
);

INVx3_ASAP7_75t_L g3442 ( 
.A(n_3113),
.Y(n_3442)
);

BUFx6f_ASAP7_75t_L g3443 ( 
.A(n_3193),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_3146),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3191),
.B(n_2829),
.Y(n_3445)
);

BUFx3_ASAP7_75t_L g3446 ( 
.A(n_3137),
.Y(n_3446)
);

BUFx6f_ASAP7_75t_L g3447 ( 
.A(n_3138),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3208),
.B(n_2330),
.Y(n_3448)
);

AND2x4_ASAP7_75t_L g3449 ( 
.A(n_3205),
.B(n_2064),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_3199),
.B(n_2829),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3293),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3169),
.Y(n_3452)
);

AND2x4_ASAP7_75t_L g3453 ( 
.A(n_3103),
.B(n_2087),
.Y(n_3453)
);

BUFx12f_ASAP7_75t_L g3454 ( 
.A(n_3229),
.Y(n_3454)
);

INVx3_ASAP7_75t_L g3455 ( 
.A(n_3119),
.Y(n_3455)
);

AND2x4_ASAP7_75t_L g3456 ( 
.A(n_3317),
.B(n_2095),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3175),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3365),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3178),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3179),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3218),
.B(n_2835),
.Y(n_3461)
);

HB1xp67_ASAP7_75t_L g3462 ( 
.A(n_3194),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3187),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3192),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3155),
.Y(n_3465)
);

NOR2xp33_ASAP7_75t_L g3466 ( 
.A(n_3144),
.B(n_2504),
.Y(n_3466)
);

AND2x4_ASAP7_75t_L g3467 ( 
.A(n_3321),
.B(n_2104),
.Y(n_3467)
);

INVx3_ASAP7_75t_L g3468 ( 
.A(n_3329),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3219),
.B(n_2835),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3158),
.Y(n_3470)
);

BUFx6f_ASAP7_75t_L g3471 ( 
.A(n_3392),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3200),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3206),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3212),
.Y(n_3474)
);

BUFx6f_ASAP7_75t_L g3475 ( 
.A(n_3423),
.Y(n_3475)
);

AND2x2_ASAP7_75t_L g3476 ( 
.A(n_3136),
.B(n_3198),
.Y(n_3476)
);

HB1xp67_ASAP7_75t_L g3477 ( 
.A(n_3107),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3223),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3235),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3162),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3239),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3250),
.Y(n_3482)
);

AND2x4_ASAP7_75t_L g3483 ( 
.A(n_3326),
.B(n_2119),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3251),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3167),
.Y(n_3485)
);

BUFx6f_ASAP7_75t_L g3486 ( 
.A(n_3105),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3253),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3285),
.Y(n_3488)
);

AND2x2_ASAP7_75t_L g3489 ( 
.A(n_3106),
.B(n_2393),
.Y(n_3489)
);

INVx5_ASAP7_75t_L g3490 ( 
.A(n_3269),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_L g3491 ( 
.A(n_3224),
.B(n_2835),
.Y(n_3491)
);

INVx2_ASAP7_75t_L g3492 ( 
.A(n_3168),
.Y(n_3492)
);

XNOR2xp5_ASAP7_75t_L g3493 ( 
.A(n_3358),
.B(n_2121),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3286),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3261),
.Y(n_3495)
);

INVxp33_ASAP7_75t_SL g3496 ( 
.A(n_3120),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_3266),
.Y(n_3497)
);

BUFx6f_ASAP7_75t_L g3498 ( 
.A(n_3124),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3273),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_3177),
.B(n_2393),
.Y(n_3500)
);

AND2x2_ASAP7_75t_L g3501 ( 
.A(n_3389),
.B(n_2427),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3182),
.Y(n_3502)
);

NAND2xp5_ASAP7_75t_L g3503 ( 
.A(n_3316),
.B(n_2837),
.Y(n_3503)
);

BUFx6f_ASAP7_75t_L g3504 ( 
.A(n_3129),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3302),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3186),
.Y(n_3506)
);

AND2x2_ASAP7_75t_L g3507 ( 
.A(n_3123),
.B(n_2427),
.Y(n_3507)
);

BUFx6f_ASAP7_75t_L g3508 ( 
.A(n_3315),
.Y(n_3508)
);

HB1xp67_ASAP7_75t_L g3509 ( 
.A(n_3108),
.Y(n_3509)
);

OR2x6_ASAP7_75t_L g3510 ( 
.A(n_3233),
.B(n_2680),
.Y(n_3510)
);

INVx2_ASAP7_75t_L g3511 ( 
.A(n_3195),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3099),
.Y(n_3512)
);

HB1xp67_ASAP7_75t_L g3513 ( 
.A(n_3154),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3109),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3330),
.Y(n_3515)
);

BUFx2_ASAP7_75t_L g3516 ( 
.A(n_3335),
.Y(n_3516)
);

AND2x4_ASAP7_75t_L g3517 ( 
.A(n_3328),
.B(n_2140),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3339),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3347),
.Y(n_3519)
);

CKINVDCx20_ASAP7_75t_R g3520 ( 
.A(n_3134),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3379),
.Y(n_3521)
);

INVx3_ASAP7_75t_L g3522 ( 
.A(n_3349),
.Y(n_3522)
);

INVx2_ASAP7_75t_L g3523 ( 
.A(n_3202),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3236),
.Y(n_3524)
);

NAND2xp33_ASAP7_75t_SL g3525 ( 
.A(n_3357),
.B(n_2158),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3319),
.B(n_2837),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3381),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3383),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3391),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3396),
.Y(n_3530)
);

BUFx6f_ASAP7_75t_L g3531 ( 
.A(n_3327),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3397),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_3380),
.Y(n_3533)
);

AND2x2_ASAP7_75t_L g3534 ( 
.A(n_3405),
.B(n_2577),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_3413),
.Y(n_3535)
);

BUFx6f_ASAP7_75t_L g3536 ( 
.A(n_3343),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3151),
.Y(n_3537)
);

HB1xp67_ASAP7_75t_L g3538 ( 
.A(n_3406),
.Y(n_3538)
);

BUFx6f_ASAP7_75t_L g3539 ( 
.A(n_3346),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3093),
.Y(n_3540)
);

AND2x6_ASAP7_75t_L g3541 ( 
.A(n_3226),
.B(n_1929),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3097),
.Y(n_3542)
);

XOR2xp5_ASAP7_75t_L g3543 ( 
.A(n_3322),
.B(n_2169),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3171),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3117),
.Y(n_3545)
);

INVx3_ASAP7_75t_L g3546 ( 
.A(n_3297),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3275),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3274),
.B(n_2577),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3276),
.Y(n_3549)
);

NOR2x1_ASAP7_75t_L g3550 ( 
.A(n_3164),
.B(n_2321),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3125),
.Y(n_3551)
);

AND2x6_ASAP7_75t_L g3552 ( 
.A(n_3254),
.B(n_1931),
.Y(n_3552)
);

INVx3_ASAP7_75t_L g3553 ( 
.A(n_3301),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3142),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3323),
.B(n_3352),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3332),
.Y(n_3556)
);

AND2x4_ASAP7_75t_SL g3557 ( 
.A(n_3341),
.B(n_2641),
.Y(n_3557)
);

INVx3_ASAP7_75t_L g3558 ( 
.A(n_3190),
.Y(n_3558)
);

AND2x4_ASAP7_75t_L g3559 ( 
.A(n_3348),
.B(n_2185),
.Y(n_3559)
);

OAI22xp5_ASAP7_75t_SL g3560 ( 
.A1(n_3264),
.A2(n_2223),
.B1(n_2235),
.B2(n_2186),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3216),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3334),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3221),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3338),
.Y(n_3564)
);

BUFx6f_ASAP7_75t_L g3565 ( 
.A(n_3378),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_L g3566 ( 
.A(n_3369),
.B(n_2837),
.Y(n_3566)
);

INVx1_ASAP7_75t_L g3567 ( 
.A(n_3240),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3243),
.Y(n_3568)
);

BUFx8_ASAP7_75t_L g3569 ( 
.A(n_3248),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3399),
.B(n_2331),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3259),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3173),
.B(n_2333),
.Y(n_3572)
);

INVx2_ASAP7_75t_SL g3573 ( 
.A(n_3354),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3271),
.Y(n_3574)
);

INVxp67_ASAP7_75t_L g3575 ( 
.A(n_3153),
.Y(n_3575)
);

BUFx2_ASAP7_75t_L g3576 ( 
.A(n_3314),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3209),
.B(n_3116),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3282),
.Y(n_3578)
);

BUFx6f_ASAP7_75t_L g3579 ( 
.A(n_3387),
.Y(n_3579)
);

AND2x4_ASAP7_75t_L g3580 ( 
.A(n_3417),
.B(n_2239),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3318),
.Y(n_3581)
);

INVx3_ASAP7_75t_L g3582 ( 
.A(n_3260),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3344),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3333),
.Y(n_3584)
);

BUFx6f_ASAP7_75t_L g3585 ( 
.A(n_3398),
.Y(n_3585)
);

AND2x4_ASAP7_75t_L g3586 ( 
.A(n_3262),
.B(n_2273),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3336),
.Y(n_3587)
);

BUFx6f_ASAP7_75t_L g3588 ( 
.A(n_3407),
.Y(n_3588)
);

INVx2_ASAP7_75t_L g3589 ( 
.A(n_3353),
.Y(n_3589)
);

BUFx2_ASAP7_75t_L g3590 ( 
.A(n_3126),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3342),
.Y(n_3591)
);

INVx1_ASAP7_75t_SL g3592 ( 
.A(n_3245),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_3420),
.B(n_1904),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3361),
.Y(n_3594)
);

BUFx3_ASAP7_75t_L g3595 ( 
.A(n_3096),
.Y(n_3595)
);

AND2x6_ASAP7_75t_L g3596 ( 
.A(n_3263),
.B(n_1999),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3296),
.B(n_2336),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3360),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3363),
.Y(n_3599)
);

INVx3_ASAP7_75t_L g3600 ( 
.A(n_3299),
.Y(n_3600)
);

INVx2_ASAP7_75t_L g3601 ( 
.A(n_3404),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3382),
.Y(n_3602)
);

AND2x4_ASAP7_75t_L g3603 ( 
.A(n_3312),
.B(n_2293),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3385),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3091),
.B(n_2339),
.Y(n_3605)
);

AND2x2_ASAP7_75t_L g3606 ( 
.A(n_3172),
.B(n_2641),
.Y(n_3606)
);

XOR2xp5_ASAP7_75t_L g3607 ( 
.A(n_3362),
.B(n_2318),
.Y(n_3607)
);

OA21x2_ASAP7_75t_L g3608 ( 
.A1(n_3127),
.A2(n_2350),
.B(n_2349),
.Y(n_3608)
);

HB1xp67_ASAP7_75t_L g3609 ( 
.A(n_3143),
.Y(n_3609)
);

INVx3_ASAP7_75t_L g3610 ( 
.A(n_3310),
.Y(n_3610)
);

OAI22xp5_ASAP7_75t_L g3611 ( 
.A1(n_3185),
.A2(n_2262),
.B1(n_2635),
.B2(n_1936),
.Y(n_3611)
);

AND2x6_ASAP7_75t_L g3612 ( 
.A(n_3325),
.B(n_2025),
.Y(n_3612)
);

BUFx6f_ASAP7_75t_L g3613 ( 
.A(n_3115),
.Y(n_3613)
);

BUFx6f_ASAP7_75t_L g3614 ( 
.A(n_3340),
.Y(n_3614)
);

BUFx4f_ASAP7_75t_L g3615 ( 
.A(n_3366),
.Y(n_3615)
);

INVx3_ASAP7_75t_L g3616 ( 
.A(n_3284),
.Y(n_3616)
);

INVx2_ASAP7_75t_L g3617 ( 
.A(n_3408),
.Y(n_3617)
);

AND2x2_ASAP7_75t_L g3618 ( 
.A(n_3188),
.B(n_2655),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3415),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3386),
.Y(n_3620)
);

NOR2xp33_ASAP7_75t_L g3621 ( 
.A(n_3147),
.B(n_1905),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3390),
.Y(n_3622)
);

AND2x4_ASAP7_75t_L g3623 ( 
.A(n_3331),
.B(n_2328),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3401),
.Y(n_3624)
);

INVx1_ASAP7_75t_L g3625 ( 
.A(n_3402),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3291),
.Y(n_3626)
);

AND2x4_ASAP7_75t_L g3627 ( 
.A(n_3350),
.B(n_2341),
.Y(n_3627)
);

INVx2_ASAP7_75t_L g3628 ( 
.A(n_3141),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3152),
.B(n_2351),
.Y(n_3629)
);

INVx1_ASAP7_75t_SL g3630 ( 
.A(n_3234),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3409),
.Y(n_3631)
);

BUFx6f_ASAP7_75t_L g3632 ( 
.A(n_3367),
.Y(n_3632)
);

BUFx6f_ASAP7_75t_L g3633 ( 
.A(n_3376),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3416),
.Y(n_3634)
);

INVx3_ASAP7_75t_L g3635 ( 
.A(n_3295),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3425),
.Y(n_3636)
);

INVx2_ASAP7_75t_L g3637 ( 
.A(n_3265),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3433),
.Y(n_3638)
);

NOR2x1_ASAP7_75t_L g3639 ( 
.A(n_3100),
.B(n_2353),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3166),
.B(n_2363),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3267),
.Y(n_3641)
);

BUFx2_ASAP7_75t_L g3642 ( 
.A(n_3148),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3268),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3279),
.Y(n_3644)
);

INVx3_ASAP7_75t_L g3645 ( 
.A(n_3307),
.Y(n_3645)
);

HB1xp67_ASAP7_75t_L g3646 ( 
.A(n_3189),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3287),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3292),
.Y(n_3648)
);

AND2x4_ASAP7_75t_L g3649 ( 
.A(n_3356),
.B(n_2366),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3294),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3300),
.Y(n_3651)
);

BUFx6f_ASAP7_75t_L g3652 ( 
.A(n_3388),
.Y(n_3652)
);

BUFx8_ASAP7_75t_L g3653 ( 
.A(n_3196),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3303),
.Y(n_3654)
);

AND2x4_ASAP7_75t_L g3655 ( 
.A(n_3368),
.B(n_2418),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3384),
.B(n_2655),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3306),
.Y(n_3657)
);

BUFx6f_ASAP7_75t_L g3658 ( 
.A(n_3149),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3309),
.Y(n_3659)
);

INVx2_ASAP7_75t_L g3660 ( 
.A(n_3311),
.Y(n_3660)
);

BUFx2_ASAP7_75t_L g3661 ( 
.A(n_3161),
.Y(n_3661)
);

OA21x2_ASAP7_75t_L g3662 ( 
.A1(n_3139),
.A2(n_2374),
.B(n_2367),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3111),
.Y(n_3663)
);

CKINVDCx5p33_ASAP7_75t_R g3664 ( 
.A(n_3257),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3181),
.B(n_2377),
.Y(n_3665)
);

INVx2_ASAP7_75t_L g3666 ( 
.A(n_3118),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3207),
.B(n_2383),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3210),
.B(n_2388),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3110),
.B(n_2389),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3230),
.Y(n_3670)
);

OR2x6_ASAP7_75t_L g3671 ( 
.A(n_3174),
.B(n_2754),
.Y(n_3671)
);

AND2x4_ASAP7_75t_L g3672 ( 
.A(n_3394),
.B(n_2437),
.Y(n_3672)
);

AND2x2_ASAP7_75t_L g3673 ( 
.A(n_3400),
.B(n_3410),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3122),
.B(n_1907),
.Y(n_3674)
);

BUFx6f_ASAP7_75t_L g3675 ( 
.A(n_3176),
.Y(n_3675)
);

OA21x2_ASAP7_75t_L g3676 ( 
.A1(n_3231),
.A2(n_2406),
.B(n_2404),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_SL g3677 ( 
.A(n_3132),
.B(n_1908),
.Y(n_3677)
);

HB1xp67_ASAP7_75t_L g3678 ( 
.A(n_3324),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3232),
.Y(n_3679)
);

XNOR2xp5_ASAP7_75t_L g3680 ( 
.A(n_3308),
.B(n_2494),
.Y(n_3680)
);

AOI22x1_ASAP7_75t_SL g3681 ( 
.A1(n_3364),
.A2(n_2500),
.B1(n_2514),
.B2(n_2497),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3426),
.B(n_3429),
.Y(n_3682)
);

NAND2xp33_ASAP7_75t_L g3683 ( 
.A(n_3359),
.B(n_1909),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_3241),
.Y(n_3684)
);

AND2x4_ASAP7_75t_L g3685 ( 
.A(n_3160),
.B(n_2532),
.Y(n_3685)
);

BUFx3_ASAP7_75t_L g3686 ( 
.A(n_3372),
.Y(n_3686)
);

INVx3_ASAP7_75t_L g3687 ( 
.A(n_3247),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3121),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3114),
.B(n_2408),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_L g3690 ( 
.A(n_3214),
.B(n_2428),
.Y(n_3690)
);

INVx3_ASAP7_75t_L g3691 ( 
.A(n_3270),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3092),
.Y(n_3692)
);

INVx2_ASAP7_75t_L g3693 ( 
.A(n_3157),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3215),
.B(n_2431),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3098),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3095),
.B(n_1913),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3104),
.Y(n_3697)
);

BUFx6f_ASAP7_75t_L g3698 ( 
.A(n_3256),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3244),
.Y(n_3699)
);

BUFx3_ASAP7_75t_L g3700 ( 
.A(n_3370),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3102),
.B(n_2432),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3252),
.Y(n_3702)
);

BUFx2_ASAP7_75t_L g3703 ( 
.A(n_3395),
.Y(n_3703)
);

BUFx6f_ASAP7_75t_L g3704 ( 
.A(n_3156),
.Y(n_3704)
);

AND2x4_ASAP7_75t_L g3705 ( 
.A(n_3163),
.B(n_3165),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3255),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_3355),
.Y(n_3707)
);

BUFx8_ASAP7_75t_L g3708 ( 
.A(n_3156),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3211),
.Y(n_3709)
);

NOR2xp33_ASAP7_75t_SL g3710 ( 
.A(n_3170),
.B(n_2537),
.Y(n_3710)
);

INVx1_ASAP7_75t_L g3711 ( 
.A(n_3217),
.Y(n_3711)
);

BUFx6f_ASAP7_75t_L g3712 ( 
.A(n_3304),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3220),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3222),
.Y(n_3714)
);

INVx4_ASAP7_75t_L g3715 ( 
.A(n_3411),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3227),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3238),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3258),
.Y(n_3718)
);

CKINVDCx8_ASAP7_75t_R g3719 ( 
.A(n_3184),
.Y(n_3719)
);

BUFx6f_ASAP7_75t_L g3720 ( 
.A(n_3412),
.Y(n_3720)
);

BUFx6f_ASAP7_75t_L g3721 ( 
.A(n_3203),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3128),
.B(n_2683),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3272),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3237),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3277),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3135),
.B(n_2683),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3281),
.Y(n_3727)
);

BUFx6f_ASAP7_75t_L g3728 ( 
.A(n_3204),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3283),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3298),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3305),
.Y(n_3731)
);

BUFx2_ASAP7_75t_L g3732 ( 
.A(n_3374),
.Y(n_3732)
);

BUFx6f_ASAP7_75t_L g3733 ( 
.A(n_3213),
.Y(n_3733)
);

BUFx6f_ASAP7_75t_L g3734 ( 
.A(n_3320),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3313),
.Y(n_3735)
);

INVx3_ASAP7_75t_L g3736 ( 
.A(n_3225),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3290),
.A2(n_2088),
.B1(n_2112),
.B2(n_2037),
.Y(n_3737)
);

INVx3_ASAP7_75t_L g3738 ( 
.A(n_3225),
.Y(n_3738)
);

INVx1_ASAP7_75t_L g3739 ( 
.A(n_3249),
.Y(n_3739)
);

AND2x4_ASAP7_75t_L g3740 ( 
.A(n_3183),
.B(n_2551),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3337),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3345),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3351),
.Y(n_3743)
);

BUFx6f_ASAP7_75t_L g3744 ( 
.A(n_3371),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3373),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3375),
.Y(n_3746)
);

AND2x4_ASAP7_75t_L g3747 ( 
.A(n_3150),
.B(n_2589),
.Y(n_3747)
);

OA21x2_ASAP7_75t_L g3748 ( 
.A1(n_3418),
.A2(n_2439),
.B(n_2435),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3377),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3393),
.Y(n_3750)
);

INVx2_ASAP7_75t_L g3751 ( 
.A(n_3419),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3421),
.Y(n_3752)
);

INVx5_ASAP7_75t_L g3753 ( 
.A(n_3197),
.Y(n_3753)
);

INVx5_ASAP7_75t_L g3754 ( 
.A(n_3201),
.Y(n_3754)
);

BUFx6f_ASAP7_75t_L g3755 ( 
.A(n_3422),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3424),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3431),
.Y(n_3757)
);

AND2x2_ASAP7_75t_L g3758 ( 
.A(n_3159),
.B(n_3403),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3432),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_SL g3760 ( 
.A(n_3414),
.B(n_1914),
.Y(n_3760)
);

NAND3xp33_ASAP7_75t_L g3761 ( 
.A(n_3228),
.B(n_1916),
.C(n_1915),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3428),
.B(n_2703),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3434),
.Y(n_3763)
);

AND2x4_ASAP7_75t_L g3764 ( 
.A(n_3094),
.B(n_2630),
.Y(n_3764)
);

INVx2_ASAP7_75t_L g3765 ( 
.A(n_3101),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3246),
.Y(n_3766)
);

INVx3_ASAP7_75t_L g3767 ( 
.A(n_3278),
.Y(n_3767)
);

OAI22xp33_ASAP7_75t_L g3768 ( 
.A1(n_3555),
.A2(n_3289),
.B1(n_2665),
.B2(n_2679),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_SL g3769 ( 
.A(n_3707),
.B(n_3430),
.Y(n_3769)
);

AND3x2_ASAP7_75t_L g3770 ( 
.A(n_3576),
.B(n_2831),
.C(n_3280),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3512),
.Y(n_3771)
);

AND2x4_ASAP7_75t_L g3772 ( 
.A(n_3443),
.B(n_3427),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3577),
.B(n_3278),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3485),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_SL g3775 ( 
.A(n_3575),
.B(n_3112),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3492),
.Y(n_3776)
);

INVx2_ASAP7_75t_L g3777 ( 
.A(n_3502),
.Y(n_3777)
);

BUFx2_ASAP7_75t_L g3778 ( 
.A(n_3516),
.Y(n_3778)
);

NAND2xp33_ASAP7_75t_L g3779 ( 
.A(n_3718),
.B(n_1918),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_3621),
.B(n_1919),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3506),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3511),
.Y(n_3782)
);

CKINVDCx5p33_ASAP7_75t_R g3783 ( 
.A(n_3664),
.Y(n_3783)
);

INVx3_ASAP7_75t_L g3784 ( 
.A(n_3446),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3514),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3523),
.Y(n_3786)
);

INVx5_ASAP7_75t_L g3787 ( 
.A(n_3613),
.Y(n_3787)
);

OA22x2_ASAP7_75t_L g3788 ( 
.A1(n_3680),
.A2(n_3288),
.B1(n_2166),
.B2(n_2171),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3524),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3441),
.Y(n_3790)
);

BUFx6f_ASAP7_75t_L g3791 ( 
.A(n_3614),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3451),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3515),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_3540),
.Y(n_3794)
);

BUFx6f_ASAP7_75t_L g3795 ( 
.A(n_3632),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3723),
.B(n_3725),
.Y(n_3796)
);

INVx1_ASAP7_75t_SL g3797 ( 
.A(n_3592),
.Y(n_3797)
);

BUFx3_ASAP7_75t_L g3798 ( 
.A(n_3454),
.Y(n_3798)
);

INVx3_ASAP7_75t_L g3799 ( 
.A(n_3447),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3552),
.A2(n_2700),
.B1(n_2717),
.B2(n_2654),
.Y(n_3800)
);

INVx2_ASAP7_75t_L g3801 ( 
.A(n_3542),
.Y(n_3801)
);

OR2x2_ASAP7_75t_L g3802 ( 
.A(n_3462),
.B(n_2128),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3518),
.Y(n_3803)
);

INVx2_ASAP7_75t_L g3804 ( 
.A(n_3545),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3519),
.Y(n_3805)
);

NOR2xp33_ASAP7_75t_L g3806 ( 
.A(n_3696),
.B(n_2172),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3521),
.Y(n_3807)
);

INVx2_ASAP7_75t_L g3808 ( 
.A(n_3551),
.Y(n_3808)
);

INVx3_ASAP7_75t_L g3809 ( 
.A(n_3458),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3556),
.Y(n_3810)
);

NAND2xp33_ASAP7_75t_L g3811 ( 
.A(n_3727),
.B(n_1923),
.Y(n_3811)
);

AOI22xp33_ASAP7_75t_L g3812 ( 
.A1(n_3552),
.A2(n_2730),
.B1(n_2757),
.B2(n_2727),
.Y(n_3812)
);

INVxp67_ASAP7_75t_SL g3813 ( 
.A(n_3513),
.Y(n_3813)
);

NAND2xp33_ASAP7_75t_SL g3814 ( 
.A(n_3715),
.B(n_2779),
.Y(n_3814)
);

NAND2xp5_ASAP7_75t_SL g3815 ( 
.A(n_3729),
.B(n_1924),
.Y(n_3815)
);

INVxp33_ASAP7_75t_SL g3816 ( 
.A(n_3686),
.Y(n_3816)
);

NAND2xp33_ASAP7_75t_SL g3817 ( 
.A(n_3618),
.B(n_2782),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3527),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_SL g3819 ( 
.A(n_3730),
.B(n_1926),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_SL g3820 ( 
.A(n_3731),
.B(n_1946),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3562),
.Y(n_3821)
);

NAND2xp5_ASAP7_75t_SL g3822 ( 
.A(n_3735),
.B(n_1947),
.Y(n_3822)
);

INVx4_ASAP7_75t_L g3823 ( 
.A(n_3633),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3564),
.Y(n_3824)
);

INVx2_ASAP7_75t_L g3825 ( 
.A(n_3583),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3589),
.Y(n_3826)
);

OAI22xp5_ASAP7_75t_L g3827 ( 
.A1(n_3739),
.A2(n_1949),
.B1(n_1952),
.B2(n_1948),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_3692),
.B(n_3695),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3697),
.B(n_1953),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3537),
.B(n_1954),
.Y(n_3830)
);

INVx2_ASAP7_75t_SL g3831 ( 
.A(n_3758),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3528),
.Y(n_3832)
);

INVx3_ASAP7_75t_L g3833 ( 
.A(n_3471),
.Y(n_3833)
);

INVxp67_ASAP7_75t_L g3834 ( 
.A(n_3538),
.Y(n_3834)
);

NAND3xp33_ASAP7_75t_L g3835 ( 
.A(n_3466),
.B(n_1968),
.C(n_1960),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3598),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3529),
.Y(n_3837)
);

AOI22xp33_ASAP7_75t_L g3838 ( 
.A1(n_3596),
.A2(n_3544),
.B1(n_3644),
.B2(n_3637),
.Y(n_3838)
);

HB1xp67_ASAP7_75t_SL g3839 ( 
.A(n_3569),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3601),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3530),
.Y(n_3841)
);

INVx3_ASAP7_75t_L g3842 ( 
.A(n_3475),
.Y(n_3842)
);

INVxp33_ASAP7_75t_L g3843 ( 
.A(n_3493),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3617),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3532),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3535),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3476),
.B(n_2787),
.Y(n_3847)
);

INVx3_ASAP7_75t_L g3848 ( 
.A(n_3486),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3663),
.B(n_1969),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3495),
.Y(n_3850)
);

INVx2_ASAP7_75t_L g3851 ( 
.A(n_3619),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3436),
.Y(n_3852)
);

BUFx3_ASAP7_75t_L g3853 ( 
.A(n_3595),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3497),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3439),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3499),
.Y(n_3856)
);

INVx3_ASAP7_75t_L g3857 ( 
.A(n_3498),
.Y(n_3857)
);

INVx2_ASAP7_75t_SL g3858 ( 
.A(n_3732),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3440),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3670),
.B(n_1974),
.Y(n_3860)
);

INVx8_ASAP7_75t_L g3861 ( 
.A(n_3658),
.Y(n_3861)
);

NAND3xp33_ASAP7_75t_L g3862 ( 
.A(n_3679),
.B(n_1977),
.C(n_1975),
.Y(n_3862)
);

BUFx6f_ASAP7_75t_L g3863 ( 
.A(n_3652),
.Y(n_3863)
);

INVx2_ASAP7_75t_L g3864 ( 
.A(n_3505),
.Y(n_3864)
);

INVx2_ASAP7_75t_L g3865 ( 
.A(n_3561),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3563),
.Y(n_3866)
);

INVx2_ASAP7_75t_SL g3867 ( 
.A(n_3705),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3567),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3684),
.B(n_1980),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3606),
.B(n_1981),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3568),
.Y(n_3871)
);

BUFx2_ASAP7_75t_L g3872 ( 
.A(n_3437),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_3571),
.Y(n_3873)
);

AND3x2_ASAP7_75t_L g3874 ( 
.A(n_3703),
.B(n_2400),
.C(n_2387),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3574),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3578),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3554),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_3699),
.B(n_1982),
.Y(n_3878)
);

INVx1_ASAP7_75t_L g3879 ( 
.A(n_3657),
.Y(n_3879)
);

AND2x2_ASAP7_75t_L g3880 ( 
.A(n_3507),
.B(n_2801),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3660),
.Y(n_3881)
);

AND2x4_ASAP7_75t_L g3882 ( 
.A(n_3590),
.B(n_2803),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3435),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3445),
.Y(n_3884)
);

INVx1_ASAP7_75t_L g3885 ( 
.A(n_3450),
.Y(n_3885)
);

AND2x2_ASAP7_75t_L g3886 ( 
.A(n_3534),
.B(n_2805),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_SL g3887 ( 
.A(n_3706),
.B(n_1985),
.Y(n_3887)
);

INVx2_ASAP7_75t_SL g3888 ( 
.A(n_3720),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_SL g3889 ( 
.A(n_3702),
.B(n_1986),
.Y(n_3889)
);

AOI21x1_ASAP7_75t_L g3890 ( 
.A1(n_3461),
.A2(n_2448),
.B(n_2446),
.Y(n_3890)
);

BUFx6f_ASAP7_75t_SL g3891 ( 
.A(n_3675),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3693),
.Y(n_3892)
);

CKINVDCx6p67_ASAP7_75t_R g3893 ( 
.A(n_3520),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3469),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3581),
.B(n_1989),
.Y(n_3895)
);

AND2x2_ASAP7_75t_L g3896 ( 
.A(n_3673),
.B(n_2826),
.Y(n_3896)
);

CKINVDCx20_ASAP7_75t_R g3897 ( 
.A(n_3700),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3608),
.Y(n_3898)
);

NOR2xp33_ASAP7_75t_L g3899 ( 
.A(n_3496),
.B(n_2177),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3584),
.B(n_1992),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3491),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3662),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3572),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_L g3904 ( 
.A(n_3587),
.B(n_1993),
.Y(n_3904)
);

BUFx6f_ASAP7_75t_L g3905 ( 
.A(n_3698),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3591),
.B(n_1994),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3641),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3701),
.B(n_1995),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3643),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_3594),
.B(n_1997),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3647),
.Y(n_3911)
);

INVx3_ASAP7_75t_L g3912 ( 
.A(n_3504),
.Y(n_3912)
);

INVx3_ASAP7_75t_L g3913 ( 
.A(n_3508),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3648),
.Y(n_3914)
);

AOI22xp33_ASAP7_75t_L g3915 ( 
.A1(n_3596),
.A2(n_2839),
.B1(n_2833),
.B2(n_2238),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3650),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3651),
.Y(n_3917)
);

INVx2_ASAP7_75t_SL g3918 ( 
.A(n_3682),
.Y(n_3918)
);

BUFx6f_ASAP7_75t_L g3919 ( 
.A(n_3615),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3547),
.Y(n_3920)
);

OR2x2_ASAP7_75t_L g3921 ( 
.A(n_3586),
.B(n_2180),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3654),
.Y(n_3922)
);

NAND2xp33_ASAP7_75t_L g3923 ( 
.A(n_3639),
.B(n_1998),
.Y(n_3923)
);

INVx3_ASAP7_75t_L g3924 ( 
.A(n_3531),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3659),
.Y(n_3925)
);

INVxp67_ASAP7_75t_SL g3926 ( 
.A(n_3721),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3549),
.Y(n_3927)
);

INVx2_ASAP7_75t_L g3928 ( 
.A(n_3558),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_SL g3929 ( 
.A(n_3582),
.B(n_2002),
.Y(n_3929)
);

OR2x6_ASAP7_75t_L g3930 ( 
.A(n_3642),
.B(n_3661),
.Y(n_3930)
);

INVx2_ASAP7_75t_L g3931 ( 
.A(n_3676),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3599),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_SL g3933 ( 
.A(n_3600),
.B(n_2003),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3626),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3602),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3766),
.Y(n_3936)
);

INVx2_ASAP7_75t_SL g3937 ( 
.A(n_3449),
.Y(n_3937)
);

NAND3xp33_ASAP7_75t_L g3938 ( 
.A(n_3570),
.B(n_2006),
.C(n_2005),
.Y(n_3938)
);

NOR2x1p5_ASAP7_75t_L g3939 ( 
.A(n_3691),
.B(n_3546),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_L g3940 ( 
.A(n_3604),
.B(n_2011),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3620),
.Y(n_3941)
);

HB1xp67_ASAP7_75t_L g3942 ( 
.A(n_3609),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3622),
.Y(n_3943)
);

BUFx3_ASAP7_75t_L g3944 ( 
.A(n_3653),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3624),
.Y(n_3945)
);

NAND2xp5_ASAP7_75t_L g3946 ( 
.A(n_3625),
.B(n_3631),
.Y(n_3946)
);

CKINVDCx5p33_ASAP7_75t_R g3947 ( 
.A(n_3630),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3634),
.Y(n_3948)
);

INVx2_ASAP7_75t_SL g3949 ( 
.A(n_3646),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3610),
.B(n_3762),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3636),
.Y(n_3951)
);

OR2x2_ASAP7_75t_L g3952 ( 
.A(n_3603),
.B(n_2268),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3638),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_SL g3954 ( 
.A(n_3689),
.B(n_2013),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3629),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3438),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3444),
.Y(n_3957)
);

NOR2xp33_ASAP7_75t_L g3958 ( 
.A(n_3656),
.B(n_2291),
.Y(n_3958)
);

NOR2xp33_ASAP7_75t_L g3959 ( 
.A(n_3448),
.B(n_2299),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3640),
.B(n_2014),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3665),
.B(n_2015),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_L g3962 ( 
.A(n_3667),
.B(n_2016),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3605),
.B(n_2019),
.Y(n_3963)
);

CKINVDCx5p33_ASAP7_75t_R g3964 ( 
.A(n_3719),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_3668),
.B(n_2024),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3669),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3465),
.Y(n_3967)
);

BUFx3_ASAP7_75t_L g3968 ( 
.A(n_3753),
.Y(n_3968)
);

BUFx6f_ASAP7_75t_L g3969 ( 
.A(n_3728),
.Y(n_3969)
);

BUFx6f_ASAP7_75t_L g3970 ( 
.A(n_3536),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3489),
.B(n_2027),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3470),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3748),
.Y(n_3973)
);

INVx2_ASAP7_75t_L g3974 ( 
.A(n_3480),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3597),
.Y(n_3975)
);

HB1xp67_ASAP7_75t_SL g3976 ( 
.A(n_3708),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3765),
.Y(n_3977)
);

INVx2_ASAP7_75t_L g3978 ( 
.A(n_3452),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_SL g3979 ( 
.A(n_3503),
.B(n_2028),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3457),
.Y(n_3980)
);

INVx2_ASAP7_75t_L g3981 ( 
.A(n_3459),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_L g3982 ( 
.A(n_3548),
.B(n_2311),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_3526),
.B(n_2036),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3460),
.Y(n_3984)
);

INVx1_ASAP7_75t_SL g3985 ( 
.A(n_3678),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3463),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3566),
.B(n_2041),
.Y(n_3987)
);

INVx2_ASAP7_75t_L g3988 ( 
.A(n_3464),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3690),
.B(n_2043),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3472),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3550),
.B(n_2044),
.Y(n_3991)
);

INVx2_ASAP7_75t_SL g3992 ( 
.A(n_3734),
.Y(n_3992)
);

CKINVDCx5p33_ASAP7_75t_R g3993 ( 
.A(n_3754),
.Y(n_3993)
);

BUFx6f_ASAP7_75t_L g3994 ( 
.A(n_3539),
.Y(n_3994)
);

INVxp33_ASAP7_75t_L g3995 ( 
.A(n_3543),
.Y(n_3995)
);

INVx3_ASAP7_75t_L g3996 ( 
.A(n_3565),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3473),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3474),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3478),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3479),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3481),
.Y(n_4001)
);

INVx2_ASAP7_75t_SL g4002 ( 
.A(n_3744),
.Y(n_4002)
);

INVx2_ASAP7_75t_L g4003 ( 
.A(n_3482),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3694),
.B(n_2045),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3484),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3501),
.B(n_2046),
.Y(n_4006)
);

OR2x6_ASAP7_75t_L g4007 ( 
.A(n_3712),
.B(n_2422),
.Y(n_4007)
);

NOR2x1p5_ASAP7_75t_L g4008 ( 
.A(n_3553),
.B(n_2047),
.Y(n_4008)
);

INVx2_ASAP7_75t_SL g4009 ( 
.A(n_3755),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3487),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3488),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3616),
.B(n_2048),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3494),
.Y(n_4013)
);

OR2x2_ASAP7_75t_L g4014 ( 
.A(n_3623),
.B(n_2355),
.Y(n_4014)
);

BUFx6f_ASAP7_75t_L g4015 ( 
.A(n_3579),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3442),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3455),
.Y(n_4017)
);

BUFx2_ASAP7_75t_L g4018 ( 
.A(n_3740),
.Y(n_4018)
);

BUFx2_ASAP7_75t_L g4019 ( 
.A(n_3685),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3468),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3522),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3533),
.B(n_2049),
.Y(n_4022)
);

AOI21x1_ASAP7_75t_L g4023 ( 
.A1(n_3674),
.A2(n_2458),
.B(n_2450),
.Y(n_4023)
);

CKINVDCx6p67_ASAP7_75t_R g4024 ( 
.A(n_3490),
.Y(n_4024)
);

INVx1_ASAP7_75t_L g4025 ( 
.A(n_3741),
.Y(n_4025)
);

BUFx2_ASAP7_75t_L g4026 ( 
.A(n_3747),
.Y(n_4026)
);

NAND3xp33_ASAP7_75t_L g4027 ( 
.A(n_3611),
.B(n_2052),
.C(n_2050),
.Y(n_4027)
);

INVx8_ASAP7_75t_L g4028 ( 
.A(n_3671),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3585),
.Y(n_4029)
);

NAND2xp33_ASAP7_75t_L g4030 ( 
.A(n_3677),
.B(n_2056),
.Y(n_4030)
);

INVx2_ASAP7_75t_L g4031 ( 
.A(n_3588),
.Y(n_4031)
);

OAI22xp33_ASAP7_75t_SL g4032 ( 
.A1(n_3710),
.A2(n_2395),
.B1(n_2415),
.B2(n_2371),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3746),
.Y(n_4033)
);

AND2x4_ASAP7_75t_L g4034 ( 
.A(n_3733),
.B(n_2509),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3749),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3666),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3752),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3756),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3761),
.B(n_2058),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3757),
.Y(n_4040)
);

INVx5_ASAP7_75t_L g4041 ( 
.A(n_3704),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3688),
.Y(n_4042)
);

BUFx2_ASAP7_75t_L g4043 ( 
.A(n_3453),
.Y(n_4043)
);

AOI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_3683),
.A2(n_2538),
.B1(n_2584),
.B2(n_2518),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_SL g4045 ( 
.A(n_3737),
.B(n_2060),
.Y(n_4045)
);

BUFx2_ASAP7_75t_L g4046 ( 
.A(n_3456),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3742),
.B(n_2062),
.Y(n_4047)
);

INVx1_ASAP7_75t_L g4048 ( 
.A(n_3759),
.Y(n_4048)
);

INVx2_ASAP7_75t_L g4049 ( 
.A(n_3724),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3743),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_SL g4051 ( 
.A(n_3525),
.B(n_2063),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3628),
.Y(n_4052)
);

INVx1_ASAP7_75t_L g4053 ( 
.A(n_3745),
.Y(n_4053)
);

AO21x2_ASAP7_75t_L g4054 ( 
.A1(n_3593),
.A2(n_2465),
.B(n_2460),
.Y(n_4054)
);

NAND2xp33_ASAP7_75t_L g4055 ( 
.A(n_3760),
.B(n_2065),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3750),
.Y(n_4056)
);

INVx2_ASAP7_75t_L g4057 ( 
.A(n_3751),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3763),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3711),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_3713),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3736),
.Y(n_4061)
);

BUFx3_ASAP7_75t_L g4062 ( 
.A(n_3573),
.Y(n_4062)
);

INVx1_ASAP7_75t_L g4063 ( 
.A(n_3716),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3738),
.Y(n_4064)
);

INVx2_ASAP7_75t_L g4065 ( 
.A(n_3767),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3709),
.Y(n_4066)
);

BUFx3_ASAP7_75t_L g4067 ( 
.A(n_3687),
.Y(n_4067)
);

INVx2_ASAP7_75t_SL g4068 ( 
.A(n_3500),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_SL g4069 ( 
.A(n_3722),
.B(n_2067),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3714),
.B(n_2073),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3717),
.B(n_3541),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_L g4072 ( 
.A(n_3541),
.B(n_2075),
.Y(n_4072)
);

NOR2xp33_ASAP7_75t_L g4073 ( 
.A(n_3806),
.B(n_3627),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3771),
.Y(n_4074)
);

BUFx3_ASAP7_75t_L g4075 ( 
.A(n_3897),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3785),
.Y(n_4076)
);

INVxp67_ASAP7_75t_SL g4077 ( 
.A(n_3778),
.Y(n_4077)
);

AND2x2_ASAP7_75t_L g4078 ( 
.A(n_3797),
.B(n_3649),
.Y(n_4078)
);

XOR2xp5_ASAP7_75t_L g4079 ( 
.A(n_3783),
.B(n_3607),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3793),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3803),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3805),
.Y(n_4082)
);

NOR2xp33_ASAP7_75t_L g4083 ( 
.A(n_3899),
.B(n_3655),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3807),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_3847),
.B(n_3896),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3774),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3818),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_3832),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3837),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3858),
.B(n_3672),
.Y(n_4090)
);

BUFx8_ASAP7_75t_L g4091 ( 
.A(n_3891),
.Y(n_4091)
);

INVx1_ASAP7_75t_L g4092 ( 
.A(n_3841),
.Y(n_4092)
);

AND2x4_ASAP7_75t_L g4093 ( 
.A(n_3853),
.B(n_3557),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3845),
.Y(n_4094)
);

INVxp33_ASAP7_75t_L g4095 ( 
.A(n_3802),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3846),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3850),
.Y(n_4097)
);

XOR2xp5_ASAP7_75t_L g4098 ( 
.A(n_3947),
.B(n_3560),
.Y(n_4098)
);

XOR2xp5_ASAP7_75t_L g4099 ( 
.A(n_3964),
.B(n_3681),
.Y(n_4099)
);

INVx2_ASAP7_75t_L g4100 ( 
.A(n_3776),
.Y(n_4100)
);

AND2x2_ASAP7_75t_L g4101 ( 
.A(n_3958),
.B(n_3726),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_3854),
.Y(n_4102)
);

OR2x2_ASAP7_75t_L g4103 ( 
.A(n_3985),
.B(n_3764),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3856),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3852),
.Y(n_4105)
);

NOR2xp33_ASAP7_75t_L g4106 ( 
.A(n_3816),
.B(n_3467),
.Y(n_4106)
);

XOR2xp5_ASAP7_75t_L g4107 ( 
.A(n_3843),
.B(n_3483),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3855),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_3859),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_3880),
.B(n_3886),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3864),
.Y(n_4111)
);

INVx1_ASAP7_75t_SL g4112 ( 
.A(n_3949),
.Y(n_4112)
);

CKINVDCx20_ASAP7_75t_R g4113 ( 
.A(n_3893),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_3959),
.B(n_3517),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3955),
.B(n_3612),
.Y(n_4115)
);

XNOR2x2_ASAP7_75t_L g4116 ( 
.A(n_4044),
.B(n_2601),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3828),
.B(n_3559),
.Y(n_4117)
);

INVx3_ASAP7_75t_L g4118 ( 
.A(n_3861),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_3982),
.B(n_3580),
.Y(n_4119)
);

INVx2_ASAP7_75t_L g4120 ( 
.A(n_3777),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3936),
.Y(n_4121)
);

NOR2xp33_ASAP7_75t_L g4122 ( 
.A(n_3834),
.B(n_3612),
.Y(n_4122)
);

NOR2xp67_ASAP7_75t_L g4123 ( 
.A(n_3787),
.B(n_3477),
.Y(n_4123)
);

INVx1_ASAP7_75t_L g4124 ( 
.A(n_3879),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3881),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3941),
.Y(n_4126)
);

BUFx3_ASAP7_75t_L g4127 ( 
.A(n_3861),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3781),
.Y(n_4128)
);

NOR2xp33_ASAP7_75t_L g4129 ( 
.A(n_3813),
.B(n_3509),
.Y(n_4129)
);

INVx1_ASAP7_75t_L g4130 ( 
.A(n_3948),
.Y(n_4130)
);

INVx2_ASAP7_75t_L g4131 ( 
.A(n_3782),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3775),
.B(n_3510),
.Y(n_4132)
);

INVxp67_ASAP7_75t_L g4133 ( 
.A(n_3942),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3951),
.Y(n_4134)
);

INVx1_ASAP7_75t_L g4135 ( 
.A(n_4025),
.Y(n_4135)
);

AND2x6_ASAP7_75t_L g4136 ( 
.A(n_3919),
.B(n_3635),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4033),
.Y(n_4137)
);

INVx2_ASAP7_75t_SL g4138 ( 
.A(n_3969),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_3787),
.B(n_3645),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4035),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_3831),
.B(n_2703),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4037),
.Y(n_4142)
);

INVx2_ASAP7_75t_L g4143 ( 
.A(n_3786),
.Y(n_4143)
);

NOR2xp33_ASAP7_75t_L g4144 ( 
.A(n_3780),
.B(n_2603),
.Y(n_4144)
);

AOI21xp5_ASAP7_75t_L g4145 ( 
.A1(n_3796),
.A2(n_2471),
.B(n_2466),
.Y(n_4145)
);

INVx1_ASAP7_75t_SL g4146 ( 
.A(n_3872),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_4038),
.Y(n_4147)
);

AND2x6_ASAP7_75t_L g4148 ( 
.A(n_3919),
.B(n_2474),
.Y(n_4148)
);

NOR2xp33_ASAP7_75t_L g4149 ( 
.A(n_3966),
.B(n_2696),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4040),
.Y(n_4150)
);

INVx2_ASAP7_75t_L g4151 ( 
.A(n_3789),
.Y(n_4151)
);

AND2x4_ASAP7_75t_SL g4152 ( 
.A(n_3823),
.B(n_2766),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4048),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4056),
.Y(n_4154)
);

INVx1_ASAP7_75t_L g4155 ( 
.A(n_4057),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_4050),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_4053),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_SL g4158 ( 
.A(n_3798),
.B(n_2740),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4058),
.Y(n_4159)
);

NOR2xp33_ASAP7_75t_L g4160 ( 
.A(n_3975),
.B(n_2753),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3790),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_3792),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3907),
.Y(n_4163)
);

NOR2xp33_ASAP7_75t_L g4164 ( 
.A(n_3918),
.B(n_2778),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_3909),
.Y(n_4165)
);

INVx1_ASAP7_75t_L g4166 ( 
.A(n_3911),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3914),
.Y(n_4167)
);

NOR2xp33_ASAP7_75t_L g4168 ( 
.A(n_3768),
.B(n_2076),
.Y(n_4168)
);

NOR2xp67_ASAP7_75t_L g4169 ( 
.A(n_4041),
.B(n_2077),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_L g4170 ( 
.A(n_3950),
.B(n_2079),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_3916),
.Y(n_4171)
);

XNOR2xp5_ASAP7_75t_L g4172 ( 
.A(n_3995),
.B(n_2082),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3917),
.Y(n_4173)
);

NAND2xp5_ASAP7_75t_L g4174 ( 
.A(n_3946),
.B(n_2475),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3922),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_3925),
.Y(n_4176)
);

OAI21xp5_ASAP7_75t_L g4177 ( 
.A1(n_3773),
.A2(n_2478),
.B(n_2477),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3932),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3935),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_3888),
.B(n_3800),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_3812),
.B(n_2766),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_3943),
.Y(n_4182)
);

BUFx6f_ASAP7_75t_SL g4183 ( 
.A(n_3944),
.Y(n_4183)
);

AND2x4_ASAP7_75t_L g4184 ( 
.A(n_3930),
.B(n_2482),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_3945),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3953),
.Y(n_4186)
);

XNOR2x1_ASAP7_75t_L g4187 ( 
.A(n_3882),
.B(n_2083),
.Y(n_4187)
);

HB1xp67_ASAP7_75t_L g4188 ( 
.A(n_3867),
.Y(n_4188)
);

NOR2xp33_ASAP7_75t_L g4189 ( 
.A(n_3971),
.B(n_2084),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3877),
.Y(n_4190)
);

XOR2xp5_ASAP7_75t_L g4191 ( 
.A(n_3993),
.B(n_2085),
.Y(n_4191)
);

AND2x6_ASAP7_75t_SL g4192 ( 
.A(n_4007),
.B(n_2483),
.Y(n_4192)
);

INVx1_ASAP7_75t_L g4193 ( 
.A(n_4059),
.Y(n_4193)
);

OR2x2_ASAP7_75t_L g4194 ( 
.A(n_3921),
.B(n_2487),
.Y(n_4194)
);

OAI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_3830),
.A2(n_2492),
.B(n_2490),
.Y(n_4195)
);

NAND2xp33_ASAP7_75t_R g4196 ( 
.A(n_3930),
.B(n_2089),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4060),
.Y(n_4197)
);

AND2x2_ASAP7_75t_L g4198 ( 
.A(n_3915),
.B(n_2863),
.Y(n_4198)
);

INVx2_ASAP7_75t_L g4199 ( 
.A(n_3977),
.Y(n_4199)
);

NAND2x1p5_ASAP7_75t_L g4200 ( 
.A(n_4041),
.B(n_3969),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_4063),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4066),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_3952),
.B(n_2863),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_3873),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_3875),
.Y(n_4205)
);

XNOR2xp5_ASAP7_75t_L g4206 ( 
.A(n_3839),
.B(n_2091),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3865),
.Y(n_4207)
);

NOR2xp33_ASAP7_75t_L g4208 ( 
.A(n_3870),
.B(n_2092),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4014),
.B(n_2869),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_3866),
.Y(n_4210)
);

INVx1_ASAP7_75t_L g4211 ( 
.A(n_3868),
.Y(n_4211)
);

NOR2xp67_ASAP7_75t_L g4212 ( 
.A(n_3784),
.B(n_2093),
.Y(n_4212)
);

BUFx3_ASAP7_75t_L g4213 ( 
.A(n_3791),
.Y(n_4213)
);

NAND2xp33_ASAP7_75t_SL g4214 ( 
.A(n_4008),
.B(n_2094),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_3871),
.Y(n_4215)
);

INVx2_ASAP7_75t_L g4216 ( 
.A(n_3794),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_3876),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3892),
.Y(n_4218)
);

CKINVDCx20_ASAP7_75t_R g4219 ( 
.A(n_4024),
.Y(n_4219)
);

INVx1_ASAP7_75t_L g4220 ( 
.A(n_3801),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3804),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_3808),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3810),
.Y(n_4223)
);

HB1xp67_ASAP7_75t_L g4224 ( 
.A(n_4018),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_3817),
.B(n_2096),
.Y(n_4225)
);

INVx2_ASAP7_75t_L g4226 ( 
.A(n_3821),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3824),
.Y(n_4227)
);

INVxp33_ASAP7_75t_L g4228 ( 
.A(n_4034),
.Y(n_4228)
);

INVxp33_ASAP7_75t_L g4229 ( 
.A(n_3905),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3825),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3826),
.Y(n_4231)
);

OAI21xp5_ASAP7_75t_L g4232 ( 
.A1(n_3849),
.A2(n_2498),
.B(n_2496),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_L g4233 ( 
.A(n_3903),
.B(n_2507),
.Y(n_4233)
);

XOR2xp5_ASAP7_75t_L g4234 ( 
.A(n_3791),
.B(n_2098),
.Y(n_4234)
);

AND2x4_ASAP7_75t_L g4235 ( 
.A(n_3992),
.B(n_4002),
.Y(n_4235)
);

XOR2xp5_ASAP7_75t_L g4236 ( 
.A(n_3795),
.B(n_2102),
.Y(n_4236)
);

BUFx3_ASAP7_75t_L g4237 ( 
.A(n_3795),
.Y(n_4237)
);

AND2x4_ASAP7_75t_L g4238 ( 
.A(n_4009),
.B(n_2515),
.Y(n_4238)
);

NOR2xp33_ASAP7_75t_SL g4239 ( 
.A(n_3863),
.B(n_2105),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_3772),
.B(n_2522),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3836),
.Y(n_4241)
);

BUFx8_ASAP7_75t_L g4242 ( 
.A(n_3863),
.Y(n_4242)
);

XNOR2xp5_ASAP7_75t_L g4243 ( 
.A(n_3976),
.B(n_2108),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_3840),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_3989),
.B(n_2523),
.Y(n_4245)
);

INVx1_ASAP7_75t_L g4246 ( 
.A(n_3844),
.Y(n_4246)
);

BUFx6f_ASAP7_75t_L g4247 ( 
.A(n_3970),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_3851),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_3934),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4004),
.B(n_2535),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_3920),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_3927),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3986),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_3990),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3999),
.Y(n_4255)
);

NOR2xp33_ASAP7_75t_L g4256 ( 
.A(n_3769),
.B(n_2109),
.Y(n_4256)
);

NOR2xp33_ASAP7_75t_SL g4257 ( 
.A(n_4028),
.B(n_2110),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_3898),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_3931),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4001),
.Y(n_4260)
);

INVx1_ASAP7_75t_L g4261 ( 
.A(n_4011),
.Y(n_4261)
);

NAND2x1p5_ASAP7_75t_L g4262 ( 
.A(n_3905),
.B(n_3799),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_3978),
.Y(n_4263)
);

INVxp67_ASAP7_75t_SL g4264 ( 
.A(n_3926),
.Y(n_4264)
);

INVx1_ASAP7_75t_L g4265 ( 
.A(n_3980),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_3981),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_4043),
.B(n_2542),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_3984),
.Y(n_4268)
);

XNOR2x2_ASAP7_75t_L g4269 ( 
.A(n_3788),
.B(n_2546),
.Y(n_4269)
);

AND2x4_ASAP7_75t_L g4270 ( 
.A(n_3939),
.B(n_2550),
.Y(n_4270)
);

XNOR2x2_ASAP7_75t_L g4271 ( 
.A(n_3827),
.B(n_2553),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_3988),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_3997),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_3998),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4000),
.Y(n_4275)
);

NAND2xp33_ASAP7_75t_R g4276 ( 
.A(n_4046),
.B(n_2111),
.Y(n_4276)
);

INVx1_ASAP7_75t_L g4277 ( 
.A(n_4003),
.Y(n_4277)
);

OR2x6_ASAP7_75t_L g4278 ( 
.A(n_4028),
.B(n_2440),
.Y(n_4278)
);

INVxp33_ASAP7_75t_L g4279 ( 
.A(n_4019),
.Y(n_4279)
);

XOR2xp5_ASAP7_75t_L g4280 ( 
.A(n_3968),
.B(n_2113),
.Y(n_4280)
);

BUFx8_ASAP7_75t_L g4281 ( 
.A(n_4026),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4005),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_4010),
.Y(n_4283)
);

INVx1_ASAP7_75t_L g4284 ( 
.A(n_4013),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_3928),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4068),
.B(n_2557),
.Y(n_4286)
);

XOR2xp5_ASAP7_75t_L g4287 ( 
.A(n_4027),
.B(n_2115),
.Y(n_4287)
);

NAND2xp33_ASAP7_75t_R g4288 ( 
.A(n_3809),
.B(n_3833),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3960),
.B(n_2563),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_3956),
.Y(n_4290)
);

INVxp33_ASAP7_75t_L g4291 ( 
.A(n_3970),
.Y(n_4291)
);

NOR2xp33_ASAP7_75t_L g4292 ( 
.A(n_4006),
.B(n_2116),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_3838),
.B(n_2570),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3957),
.Y(n_4294)
);

INVxp67_ASAP7_75t_L g4295 ( 
.A(n_4071),
.Y(n_4295)
);

INVxp67_ASAP7_75t_SL g4296 ( 
.A(n_3842),
.Y(n_4296)
);

NOR2xp33_ASAP7_75t_L g4297 ( 
.A(n_3878),
.B(n_2117),
.Y(n_4297)
);

OAI21xp5_ASAP7_75t_L g4298 ( 
.A1(n_3829),
.A2(n_2586),
.B(n_2583),
.Y(n_4298)
);

INVxp33_ASAP7_75t_SL g4299 ( 
.A(n_4062),
.Y(n_4299)
);

BUFx6f_ASAP7_75t_SL g4300 ( 
.A(n_4007),
.Y(n_4300)
);

AOI21xp5_ASAP7_75t_L g4301 ( 
.A1(n_3987),
.A2(n_2596),
.B(n_2590),
.Y(n_4301)
);

BUFx3_ASAP7_75t_L g4302 ( 
.A(n_3994),
.Y(n_4302)
);

AND2x4_ASAP7_75t_L g4303 ( 
.A(n_3937),
.B(n_2598),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_3967),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_3973),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_3961),
.B(n_2599),
.Y(n_4306)
);

AND2x2_ASAP7_75t_L g4307 ( 
.A(n_3962),
.B(n_2607),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_3972),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_3974),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_3902),
.Y(n_4310)
);

INVx1_ASAP7_75t_L g4311 ( 
.A(n_4052),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4049),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4036),
.Y(n_4313)
);

INVx2_ASAP7_75t_L g4314 ( 
.A(n_4042),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_4016),
.Y(n_4315)
);

AND2x2_ASAP7_75t_SL g4316 ( 
.A(n_3779),
.B(n_2469),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4017),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4020),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4021),
.Y(n_4319)
);

INVx1_ASAP7_75t_L g4320 ( 
.A(n_4061),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4064),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4065),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3890),
.Y(n_4323)
);

INVx1_ASAP7_75t_L g4324 ( 
.A(n_3883),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_3884),
.Y(n_4325)
);

NAND2xp33_ASAP7_75t_R g4326 ( 
.A(n_3770),
.B(n_2118),
.Y(n_4326)
);

OR2x6_ASAP7_75t_L g4327 ( 
.A(n_3994),
.B(n_2501),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_3885),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3894),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_3901),
.Y(n_4330)
);

INVx1_ASAP7_75t_L g4331 ( 
.A(n_3895),
.Y(n_4331)
);

INVx1_ASAP7_75t_L g4332 ( 
.A(n_3900),
.Y(n_4332)
);

NOR2xp33_ASAP7_75t_L g4333 ( 
.A(n_3887),
.B(n_2120),
.Y(n_4333)
);

NOR2xp33_ASAP7_75t_L g4334 ( 
.A(n_3954),
.B(n_2123),
.Y(n_4334)
);

NOR2xp33_ASAP7_75t_L g4335 ( 
.A(n_3815),
.B(n_2124),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_3904),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_L g4337 ( 
.A(n_3965),
.B(n_2608),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3906),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_3910),
.Y(n_4339)
);

INVx2_ASAP7_75t_L g4340 ( 
.A(n_4023),
.Y(n_4340)
);

CKINVDCx16_ASAP7_75t_R g4341 ( 
.A(n_3814),
.Y(n_4341)
);

INVxp67_ASAP7_75t_SL g4342 ( 
.A(n_4067),
.Y(n_4342)
);

NAND2x1p5_ASAP7_75t_L g4343 ( 
.A(n_4015),
.B(n_2614),
.Y(n_4343)
);

HB1xp67_ASAP7_75t_L g4344 ( 
.A(n_4015),
.Y(n_4344)
);

XOR2xp5_ASAP7_75t_L g4345 ( 
.A(n_3835),
.B(n_2125),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3940),
.Y(n_4346)
);

AND2x2_ASAP7_75t_L g4347 ( 
.A(n_3860),
.B(n_2616),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4054),
.Y(n_4348)
);

OAI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_3869),
.A2(n_2623),
.B(n_2622),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4047),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4070),
.Y(n_4351)
);

CKINVDCx5p33_ASAP7_75t_R g4352 ( 
.A(n_3848),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4012),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3889),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3862),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3991),
.Y(n_4356)
);

CKINVDCx20_ASAP7_75t_R g4357 ( 
.A(n_3857),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3963),
.Y(n_4358)
);

INVx2_ASAP7_75t_SL g4359 ( 
.A(n_3912),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_3938),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_3811),
.B(n_2628),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4029),
.Y(n_4362)
);

XOR2xp5_ASAP7_75t_L g4363 ( 
.A(n_4032),
.B(n_4051),
.Y(n_4363)
);

AND2x2_ASAP7_75t_L g4364 ( 
.A(n_4072),
.B(n_2629),
.Y(n_4364)
);

NAND2xp33_ASAP7_75t_R g4365 ( 
.A(n_3874),
.B(n_2127),
.Y(n_4365)
);

NOR2xp33_ASAP7_75t_L g4366 ( 
.A(n_3819),
.B(n_2129),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4022),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_3908),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_3923),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_4031),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_3913),
.Y(n_4371)
);

XOR2x2_ASAP7_75t_L g4372 ( 
.A(n_4045),
.B(n_4069),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_3820),
.Y(n_4373)
);

INVx8_ASAP7_75t_L g4374 ( 
.A(n_4183),
.Y(n_4374)
);

INVxp67_ASAP7_75t_L g4375 ( 
.A(n_4077),
.Y(n_4375)
);

NOR2xp67_ASAP7_75t_L g4376 ( 
.A(n_4118),
.B(n_3924),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4105),
.Y(n_4377)
);

NAND2xp33_ASAP7_75t_L g4378 ( 
.A(n_4331),
.B(n_4039),
.Y(n_4378)
);

NAND2xp5_ASAP7_75t_L g4379 ( 
.A(n_4144),
.B(n_3822),
.Y(n_4379)
);

INVx1_ASAP7_75t_L g4380 ( 
.A(n_4163),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_SL g4381 ( 
.A(n_4112),
.B(n_3929),
.Y(n_4381)
);

NOR2xp67_ASAP7_75t_L g4382 ( 
.A(n_4127),
.B(n_3996),
.Y(n_4382)
);

INVx2_ASAP7_75t_SL g4383 ( 
.A(n_4075),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_4073),
.B(n_4149),
.Y(n_4384)
);

NOR2xp33_ASAP7_75t_L g4385 ( 
.A(n_4083),
.B(n_3933),
.Y(n_4385)
);

NOR2xp33_ASAP7_75t_L g4386 ( 
.A(n_4332),
.B(n_4336),
.Y(n_4386)
);

A2O1A1Ixp33_ASAP7_75t_L g4387 ( 
.A1(n_4195),
.A2(n_4055),
.B(n_4030),
.C(n_3983),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4160),
.B(n_3979),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_4338),
.B(n_2131),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_4339),
.B(n_2134),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4108),
.Y(n_4391)
);

NAND2xp5_ASAP7_75t_L g4392 ( 
.A(n_4346),
.B(n_2136),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4165),
.Y(n_4393)
);

OR2x2_ASAP7_75t_L g4394 ( 
.A(n_4103),
.B(n_2137),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_4101),
.B(n_2139),
.Y(n_4395)
);

NAND2xp5_ASAP7_75t_L g4396 ( 
.A(n_4292),
.B(n_2147),
.Y(n_4396)
);

AOI22xp33_ASAP7_75t_L g4397 ( 
.A1(n_4181),
.A2(n_2149),
.B1(n_2155),
.B2(n_2148),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4166),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_4316),
.B(n_4307),
.Y(n_4399)
);

OR2x6_ASAP7_75t_L g4400 ( 
.A(n_4200),
.B(n_2508),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4109),
.Y(n_4401)
);

BUFx6f_ASAP7_75t_L g4402 ( 
.A(n_4247),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_4167),
.Y(n_4403)
);

INVx2_ASAP7_75t_SL g4404 ( 
.A(n_4242),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4171),
.B(n_2156),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_SL g4406 ( 
.A(n_4299),
.B(n_2157),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_SL g4407 ( 
.A(n_4129),
.B(n_2159),
.Y(n_4407)
);

NAND2x1p5_ASAP7_75t_L g4408 ( 
.A(n_4213),
.B(n_2633),
.Y(n_4408)
);

AND2x6_ASAP7_75t_L g4409 ( 
.A(n_4324),
.B(n_2642),
.Y(n_4409)
);

INVx2_ASAP7_75t_L g4410 ( 
.A(n_4111),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_4173),
.B(n_2161),
.Y(n_4411)
);

BUFx2_ASAP7_75t_L g4412 ( 
.A(n_4281),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4175),
.B(n_2162),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_L g4414 ( 
.A1(n_4085),
.A2(n_2165),
.B1(n_2167),
.B2(n_2163),
.Y(n_4414)
);

NOR2xp67_ASAP7_75t_L g4415 ( 
.A(n_4106),
.B(n_2170),
.Y(n_4415)
);

AND2x4_ASAP7_75t_L g4416 ( 
.A(n_4093),
.B(n_2647),
.Y(n_4416)
);

NAND2xp33_ASAP7_75t_L g4417 ( 
.A(n_4353),
.B(n_2173),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_4133),
.B(n_2179),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_L g4419 ( 
.A(n_4176),
.B(n_4178),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_4179),
.B(n_2181),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_L g4421 ( 
.A(n_4182),
.B(n_2182),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4185),
.B(n_2183),
.Y(n_4422)
);

BUFx6f_ASAP7_75t_L g4423 ( 
.A(n_4247),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_4245),
.A2(n_2662),
.B(n_2659),
.Y(n_4424)
);

OR2x2_ASAP7_75t_L g4425 ( 
.A(n_4146),
.B(n_2187),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_SL g4426 ( 
.A(n_4122),
.B(n_2188),
.Y(n_4426)
);

AOI22xp5_ASAP7_75t_L g4427 ( 
.A1(n_4168),
.A2(n_2192),
.B1(n_2194),
.B2(n_2191),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4186),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4350),
.B(n_2196),
.Y(n_4429)
);

INVx2_ASAP7_75t_L g4430 ( 
.A(n_4126),
.Y(n_4430)
);

NAND2x1p5_ASAP7_75t_L g4431 ( 
.A(n_4237),
.B(n_2668),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4110),
.B(n_2197),
.Y(n_4432)
);

INVx1_ASAP7_75t_L g4433 ( 
.A(n_4074),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4351),
.B(n_2199),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_4347),
.B(n_2200),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_4232),
.B(n_2201),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4076),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_4298),
.B(n_2204),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_4349),
.B(n_2205),
.Y(n_4439)
);

NOR3xp33_ASAP7_75t_L g4440 ( 
.A(n_4335),
.B(n_2676),
.C(n_2675),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4325),
.B(n_2207),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_L g4442 ( 
.A(n_4328),
.B(n_2210),
.Y(n_4442)
);

BUFx6f_ASAP7_75t_L g4443 ( 
.A(n_4302),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4329),
.B(n_2211),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4080),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_4130),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_4081),
.Y(n_4447)
);

AOI21xp5_ASAP7_75t_L g4448 ( 
.A1(n_4250),
.A2(n_2687),
.B(n_2681),
.Y(n_4448)
);

A2O1A1Ixp33_ASAP7_75t_L g4449 ( 
.A1(n_4355),
.A2(n_2702),
.B(n_2704),
.C(n_2699),
.Y(n_4449)
);

AND2x2_ASAP7_75t_L g4450 ( 
.A(n_4114),
.B(n_2213),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_4134),
.Y(n_4451)
);

INVx2_ASAP7_75t_SL g4452 ( 
.A(n_4139),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_SL g4453 ( 
.A(n_4257),
.B(n_2216),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4330),
.B(n_2218),
.Y(n_4454)
);

BUFx3_ASAP7_75t_L g4455 ( 
.A(n_4091),
.Y(n_4455)
);

NOR2xp33_ASAP7_75t_R g4456 ( 
.A(n_4113),
.B(n_2221),
.Y(n_4456)
);

AOI22xp5_ASAP7_75t_L g4457 ( 
.A1(n_4090),
.A2(n_2225),
.B1(n_2228),
.B2(n_2224),
.Y(n_4457)
);

HB1xp67_ASAP7_75t_L g4458 ( 
.A(n_4224),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4082),
.Y(n_4459)
);

NAND2xp5_ASAP7_75t_L g4460 ( 
.A(n_4174),
.B(n_4084),
.Y(n_4460)
);

INVx2_ASAP7_75t_L g4461 ( 
.A(n_4207),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4225),
.A2(n_2232),
.B1(n_2233),
.B2(n_2230),
.Y(n_4462)
);

INVxp67_ASAP7_75t_L g4463 ( 
.A(n_4078),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_SL g4464 ( 
.A(n_4119),
.B(n_2236),
.Y(n_4464)
);

INVx2_ASAP7_75t_L g4465 ( 
.A(n_4210),
.Y(n_4465)
);

INVx2_ASAP7_75t_SL g4466 ( 
.A(n_4352),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_SL g4467 ( 
.A(n_4341),
.B(n_2237),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_SL g4468 ( 
.A(n_4138),
.B(n_2241),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_SL g4469 ( 
.A(n_4235),
.B(n_2242),
.Y(n_4469)
);

NAND2xp5_ASAP7_75t_L g4470 ( 
.A(n_4087),
.B(n_2245),
.Y(n_4470)
);

AOI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4117),
.A2(n_2247),
.B1(n_2248),
.B2(n_2246),
.Y(n_4471)
);

INVx1_ASAP7_75t_L g4472 ( 
.A(n_4088),
.Y(n_4472)
);

NAND2xp5_ASAP7_75t_SL g4473 ( 
.A(n_4239),
.B(n_2251),
.Y(n_4473)
);

INVx2_ASAP7_75t_L g4474 ( 
.A(n_4211),
.Y(n_4474)
);

INVx1_ASAP7_75t_L g4475 ( 
.A(n_4089),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4092),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4203),
.B(n_2253),
.Y(n_4477)
);

NAND2xp5_ASAP7_75t_L g4478 ( 
.A(n_4094),
.B(n_2260),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4096),
.B(n_2263),
.Y(n_4479)
);

INVx2_ASAP7_75t_SL g4480 ( 
.A(n_4136),
.Y(n_4480)
);

INVxp33_ASAP7_75t_L g4481 ( 
.A(n_4095),
.Y(n_4481)
);

NOR2xp33_ASAP7_75t_SL g4482 ( 
.A(n_4219),
.B(n_2264),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4097),
.B(n_2266),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_SL g4484 ( 
.A(n_4132),
.B(n_2267),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_4102),
.B(n_2270),
.Y(n_4485)
);

NOR2xp33_ASAP7_75t_L g4486 ( 
.A(n_4228),
.B(n_2271),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4215),
.Y(n_4487)
);

O2A1O1Ixp5_ASAP7_75t_L g4488 ( 
.A1(n_4289),
.A2(n_2714),
.B(n_2716),
.C(n_2710),
.Y(n_4488)
);

INVx2_ASAP7_75t_SL g4489 ( 
.A(n_4136),
.Y(n_4489)
);

NOR2xp33_ASAP7_75t_L g4490 ( 
.A(n_4279),
.B(n_2272),
.Y(n_4490)
);

NOR2xp33_ASAP7_75t_L g4491 ( 
.A(n_4115),
.B(n_2275),
.Y(n_4491)
);

BUFx6f_ASAP7_75t_L g4492 ( 
.A(n_4262),
.Y(n_4492)
);

INVx1_ASAP7_75t_L g4493 ( 
.A(n_4104),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_SL g4494 ( 
.A(n_4256),
.B(n_2276),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_4293),
.B(n_2278),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_SL g4496 ( 
.A(n_4164),
.B(n_2279),
.Y(n_4496)
);

NOR2xp33_ASAP7_75t_SL g4497 ( 
.A(n_4300),
.B(n_2281),
.Y(n_4497)
);

OAI22xp33_ASAP7_75t_L g4498 ( 
.A1(n_4361),
.A2(n_2285),
.B1(n_2286),
.B2(n_2282),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4135),
.B(n_2287),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_4137),
.B(n_2289),
.Y(n_4500)
);

O2A1O1Ixp33_ASAP7_75t_L g4501 ( 
.A1(n_4306),
.A2(n_2726),
.B(n_2729),
.C(n_2723),
.Y(n_4501)
);

NAND2xp5_ASAP7_75t_SL g4502 ( 
.A(n_4184),
.B(n_2290),
.Y(n_4502)
);

AND2x2_ASAP7_75t_L g4503 ( 
.A(n_4209),
.B(n_2295),
.Y(n_4503)
);

INVx1_ASAP7_75t_SL g4504 ( 
.A(n_4357),
.Y(n_4504)
);

NAND2xp33_ASAP7_75t_L g4505 ( 
.A(n_4373),
.B(n_2296),
.Y(n_4505)
);

NOR2xp67_ASAP7_75t_L g4506 ( 
.A(n_4295),
.B(n_2300),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4240),
.B(n_2301),
.Y(n_4507)
);

BUFx8_ASAP7_75t_L g4508 ( 
.A(n_4148),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_4140),
.B(n_2302),
.Y(n_4509)
);

INVx2_ASAP7_75t_SL g4510 ( 
.A(n_4136),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_SL g4511 ( 
.A(n_4177),
.B(n_2306),
.Y(n_4511)
);

AOI22xp33_ASAP7_75t_L g4512 ( 
.A1(n_4198),
.A2(n_2309),
.B1(n_2310),
.B2(n_2307),
.Y(n_4512)
);

INVx2_ASAP7_75t_L g4513 ( 
.A(n_4217),
.Y(n_4513)
);

INVx2_ASAP7_75t_L g4514 ( 
.A(n_4161),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4142),
.B(n_2312),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4147),
.B(n_2313),
.Y(n_4516)
);

AND2x2_ASAP7_75t_L g4517 ( 
.A(n_4267),
.B(n_2314),
.Y(n_4517)
);

AND2x2_ASAP7_75t_L g4518 ( 
.A(n_4180),
.B(n_2316),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4150),
.B(n_4153),
.Y(n_4519)
);

INVx1_ASAP7_75t_L g4520 ( 
.A(n_4193),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_4197),
.B(n_2317),
.Y(n_4521)
);

AOI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_4337),
.A2(n_2737),
.B(n_2733),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4201),
.B(n_2319),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_4162),
.Y(n_4524)
);

BUFx5_ASAP7_75t_L g4525 ( 
.A(n_4121),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4364),
.B(n_4233),
.Y(n_4526)
);

NAND2xp33_ASAP7_75t_L g4527 ( 
.A(n_4360),
.B(n_2320),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4124),
.B(n_4125),
.Y(n_4528)
);

HB1xp67_ASAP7_75t_L g4529 ( 
.A(n_4188),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_4204),
.Y(n_4530)
);

AOI22xp5_ASAP7_75t_L g4531 ( 
.A1(n_4287),
.A2(n_2324),
.B1(n_2325),
.B2(n_2322),
.Y(n_4531)
);

NAND2xp5_ASAP7_75t_SL g4532 ( 
.A(n_4158),
.B(n_2326),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4156),
.Y(n_4533)
);

NAND2x1_ASAP7_75t_L g4534 ( 
.A(n_4320),
.B(n_2738),
.Y(n_4534)
);

AOI21xp5_ASAP7_75t_L g4535 ( 
.A1(n_4358),
.A2(n_2744),
.B(n_2739),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4205),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_4264),
.B(n_4253),
.Y(n_4537)
);

AND2x4_ASAP7_75t_L g4538 ( 
.A(n_4342),
.B(n_2748),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_SL g4539 ( 
.A(n_4270),
.B(n_2329),
.Y(n_4539)
);

AND2x6_ASAP7_75t_SL g4540 ( 
.A(n_4278),
.B(n_4327),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_SL g4541 ( 
.A(n_4297),
.B(n_2334),
.Y(n_4541)
);

NAND2xp5_ASAP7_75t_L g4542 ( 
.A(n_4254),
.B(n_4255),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4260),
.B(n_4261),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4368),
.A2(n_2338),
.B1(n_2342),
.B2(n_2335),
.Y(n_4544)
);

AND2x6_ASAP7_75t_SL g4545 ( 
.A(n_4278),
.B(n_2755),
.Y(n_4545)
);

OAI22xp33_ASAP7_75t_L g4546 ( 
.A1(n_4196),
.A2(n_2345),
.B1(n_2346),
.B2(n_2343),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_SL g4547 ( 
.A(n_4123),
.B(n_2347),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4157),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_L g4549 ( 
.A(n_4251),
.B(n_2348),
.Y(n_4549)
);

NOR2xp33_ASAP7_75t_L g4550 ( 
.A(n_4271),
.B(n_2356),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_SL g4551 ( 
.A(n_4333),
.B(n_2357),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4252),
.B(n_2358),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_4159),
.B(n_4202),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_4116),
.A2(n_2360),
.B1(n_2362),
.B2(n_2359),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4141),
.B(n_2364),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4154),
.Y(n_4556)
);

NOR3xp33_ASAP7_75t_L g4557 ( 
.A(n_4366),
.B(n_2767),
.C(n_2764),
.Y(n_4557)
);

NAND2xp5_ASAP7_75t_L g4558 ( 
.A(n_4190),
.B(n_2365),
.Y(n_4558)
);

OR2x6_ASAP7_75t_L g4559 ( 
.A(n_4327),
.B(n_2511),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4155),
.B(n_2368),
.Y(n_4560)
);

OR2x2_ASAP7_75t_L g4561 ( 
.A(n_4194),
.B(n_2369),
.Y(n_4561)
);

INVx2_ASAP7_75t_L g4562 ( 
.A(n_4086),
.Y(n_4562)
);

AOI22xp33_ASAP7_75t_SL g4563 ( 
.A1(n_4187),
.A2(n_4269),
.B1(n_4189),
.B2(n_4208),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_SL g4564 ( 
.A(n_4291),
.B(n_2370),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4354),
.B(n_2372),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4100),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4286),
.B(n_2373),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4303),
.B(n_2375),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_4263),
.B(n_2376),
.Y(n_4569)
);

INVx2_ASAP7_75t_SL g4570 ( 
.A(n_4344),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4265),
.Y(n_4571)
);

AOI22xp33_ASAP7_75t_L g4572 ( 
.A1(n_4363),
.A2(n_2379),
.B1(n_2380),
.B2(n_2378),
.Y(n_4572)
);

OR2x2_ASAP7_75t_L g4573 ( 
.A(n_4107),
.B(n_2381),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4266),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4120),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4268),
.Y(n_4576)
);

BUFx6f_ASAP7_75t_L g4577 ( 
.A(n_4359),
.Y(n_4577)
);

INVx1_ASAP7_75t_L g4578 ( 
.A(n_4272),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4273),
.B(n_2385),
.Y(n_4579)
);

NOR2xp33_ASAP7_75t_L g4580 ( 
.A(n_4356),
.B(n_2390),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4274),
.Y(n_4581)
);

AOI22xp5_ASAP7_75t_L g4582 ( 
.A1(n_4334),
.A2(n_4276),
.B1(n_4372),
.B2(n_4288),
.Y(n_4582)
);

NAND2xp5_ASAP7_75t_L g4583 ( 
.A(n_4275),
.B(n_2391),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_L g4584 ( 
.A(n_4277),
.B(n_2392),
.Y(n_4584)
);

INVxp67_ASAP7_75t_SL g4585 ( 
.A(n_4296),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_SL g4586 ( 
.A(n_4169),
.B(n_2394),
.Y(n_4586)
);

NAND2xp5_ASAP7_75t_L g4587 ( 
.A(n_4282),
.B(n_2396),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4283),
.B(n_2397),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4238),
.B(n_4343),
.Y(n_4589)
);

BUFx3_ASAP7_75t_L g4590 ( 
.A(n_4371),
.Y(n_4590)
);

NOR2xp33_ASAP7_75t_L g4591 ( 
.A(n_4369),
.B(n_2398),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_SL g4592 ( 
.A(n_4229),
.B(n_2399),
.Y(n_4592)
);

NOR2xp33_ASAP7_75t_L g4593 ( 
.A(n_4367),
.B(n_2401),
.Y(n_4593)
);

BUFx8_ASAP7_75t_L g4594 ( 
.A(n_4148),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4284),
.Y(n_4595)
);

OAI22xp5_ASAP7_75t_L g4596 ( 
.A1(n_4315),
.A2(n_2405),
.B1(n_2407),
.B2(n_2403),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4128),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_4199),
.B(n_2410),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_4218),
.B(n_2411),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4249),
.B(n_2413),
.Y(n_4600)
);

INVx1_ASAP7_75t_L g4601 ( 
.A(n_4220),
.Y(n_4601)
);

NAND2xp5_ASAP7_75t_L g4602 ( 
.A(n_4221),
.B(n_2414),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_4131),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_L g4604 ( 
.A(n_4222),
.B(n_2419),
.Y(n_4604)
);

INVx2_ASAP7_75t_L g4605 ( 
.A(n_4143),
.Y(n_4605)
);

NOR2xp67_ASAP7_75t_L g4606 ( 
.A(n_4285),
.B(n_2420),
.Y(n_4606)
);

AOI22xp5_ASAP7_75t_L g4607 ( 
.A1(n_4345),
.A2(n_2423),
.B1(n_2425),
.B2(n_2421),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4223),
.B(n_2426),
.Y(n_4608)
);

BUFx8_ASAP7_75t_L g4609 ( 
.A(n_4148),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4151),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4227),
.B(n_2429),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4230),
.B(n_4231),
.Y(n_4612)
);

AND2x2_ASAP7_75t_L g4613 ( 
.A(n_4172),
.B(n_2433),
.Y(n_4613)
);

NAND2xp5_ASAP7_75t_SL g4614 ( 
.A(n_4212),
.B(n_2434),
.Y(n_4614)
);

INVx1_ASAP7_75t_L g4615 ( 
.A(n_4241),
.Y(n_4615)
);

NOR2xp33_ASAP7_75t_L g4616 ( 
.A(n_4319),
.B(n_2436),
.Y(n_4616)
);

INVx2_ASAP7_75t_SL g4617 ( 
.A(n_4152),
.Y(n_4617)
);

NAND2xp5_ASAP7_75t_SL g4618 ( 
.A(n_4170),
.B(n_2438),
.Y(n_4618)
);

NOR2xp67_ASAP7_75t_L g4619 ( 
.A(n_4321),
.B(n_2441),
.Y(n_4619)
);

NOR2xp33_ASAP7_75t_L g4620 ( 
.A(n_4322),
.B(n_2442),
.Y(n_4620)
);

INVx2_ASAP7_75t_SL g4621 ( 
.A(n_4079),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4244),
.B(n_2443),
.Y(n_4622)
);

NOR2xp33_ASAP7_75t_SL g4623 ( 
.A(n_4098),
.B(n_2444),
.Y(n_4623)
);

NOR2xp67_ASAP7_75t_L g4624 ( 
.A(n_4362),
.B(n_2445),
.Y(n_4624)
);

NAND2xp5_ASAP7_75t_L g4625 ( 
.A(n_4246),
.B(n_2447),
.Y(n_4625)
);

INVxp67_ASAP7_75t_L g4626 ( 
.A(n_4234),
.Y(n_4626)
);

AOI22xp5_ASAP7_75t_L g4627 ( 
.A1(n_4214),
.A2(n_2451),
.B1(n_2453),
.B2(n_2449),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4216),
.Y(n_4628)
);

INVx5_ASAP7_75t_L g4629 ( 
.A(n_4192),
.Y(n_4629)
);

INVx3_ASAP7_75t_L g4630 ( 
.A(n_4370),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_4317),
.B(n_2454),
.Y(n_4631)
);

INVx1_ASAP7_75t_L g4632 ( 
.A(n_4226),
.Y(n_4632)
);

INVxp33_ASAP7_75t_L g4633 ( 
.A(n_4236),
.Y(n_4633)
);

AOI22xp5_ASAP7_75t_L g4634 ( 
.A1(n_4191),
.A2(n_2459),
.B1(n_2461),
.B2(n_2456),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_SL g4635 ( 
.A(n_4318),
.B(n_2462),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4248),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4314),
.B(n_2463),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_4258),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_4243),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4311),
.B(n_2467),
.Y(n_4640)
);

NAND2xp33_ASAP7_75t_L g4641 ( 
.A(n_4340),
.B(n_2470),
.Y(n_4641)
);

INVx3_ASAP7_75t_L g4642 ( 
.A(n_4312),
.Y(n_4642)
);

INVx2_ASAP7_75t_L g4643 ( 
.A(n_4259),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4313),
.B(n_2473),
.Y(n_4644)
);

BUFx6f_ASAP7_75t_L g4645 ( 
.A(n_4290),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4301),
.B(n_2479),
.Y(n_4646)
);

INVx2_ASAP7_75t_L g4647 ( 
.A(n_4305),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4294),
.B(n_2480),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4304),
.B(n_2484),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4308),
.Y(n_4650)
);

AND2x4_ASAP7_75t_L g4651 ( 
.A(n_4309),
.B(n_2768),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_SL g4652 ( 
.A(n_4145),
.B(n_4206),
.Y(n_4652)
);

AOI22xp5_ASAP7_75t_L g4653 ( 
.A1(n_4365),
.A2(n_2488),
.B1(n_2489),
.B2(n_2486),
.Y(n_4653)
);

INVxp67_ASAP7_75t_L g4654 ( 
.A(n_4280),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_SL g4655 ( 
.A(n_4348),
.B(n_4323),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_L g4656 ( 
.A(n_4310),
.B(n_2491),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4099),
.Y(n_4657)
);

INVx2_ASAP7_75t_L g4658 ( 
.A(n_4326),
.Y(n_4658)
);

INVx1_ASAP7_75t_L g4659 ( 
.A(n_4163),
.Y(n_4659)
);

INVx1_ASAP7_75t_L g4660 ( 
.A(n_4163),
.Y(n_4660)
);

NOR2xp33_ASAP7_75t_SL g4661 ( 
.A(n_4127),
.B(n_2495),
.Y(n_4661)
);

NOR2xp33_ASAP7_75t_L g4662 ( 
.A(n_4073),
.B(n_2499),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4144),
.B(n_2502),
.Y(n_4663)
);

NAND2xp33_ASAP7_75t_L g4664 ( 
.A(n_4331),
.B(n_2503),
.Y(n_4664)
);

INVx2_ASAP7_75t_SL g4665 ( 
.A(n_4127),
.Y(n_4665)
);

INVx4_ASAP7_75t_L g4666 ( 
.A(n_4127),
.Y(n_4666)
);

AOI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_4460),
.A2(n_4387),
.B(n_4641),
.Y(n_4667)
);

INVx1_ASAP7_75t_L g4668 ( 
.A(n_4528),
.Y(n_4668)
);

NAND2xp5_ASAP7_75t_L g4669 ( 
.A(n_4384),
.B(n_2505),
.Y(n_4669)
);

AO21x1_ASAP7_75t_L g4670 ( 
.A1(n_4511),
.A2(n_2783),
.B(n_2773),
.Y(n_4670)
);

AOI21xp5_ASAP7_75t_L g4671 ( 
.A1(n_4378),
.A2(n_2792),
.B(n_2791),
.Y(n_4671)
);

NOR2xp33_ASAP7_75t_L g4672 ( 
.A(n_4385),
.B(n_2506),
.Y(n_4672)
);

AO21x1_ASAP7_75t_L g4673 ( 
.A1(n_4379),
.A2(n_2796),
.B(n_2793),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4386),
.B(n_2510),
.Y(n_4674)
);

AOI21xp5_ASAP7_75t_L g4675 ( 
.A1(n_4419),
.A2(n_4542),
.B(n_4519),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4662),
.B(n_2512),
.Y(n_4676)
);

A2O1A1Ixp33_ASAP7_75t_L g4677 ( 
.A1(n_4396),
.A2(n_2814),
.B(n_2817),
.C(n_2800),
.Y(n_4677)
);

OAI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_4663),
.A2(n_4591),
.B(n_4438),
.Y(n_4678)
);

AOI21xp5_ASAP7_75t_L g4679 ( 
.A1(n_4543),
.A2(n_2819),
.B(n_2818),
.Y(n_4679)
);

AOI21xp5_ASAP7_75t_L g4680 ( 
.A1(n_4537),
.A2(n_2827),
.B(n_2824),
.Y(n_4680)
);

AND2x2_ASAP7_75t_L g4681 ( 
.A(n_4517),
.B(n_2513),
.Y(n_4681)
);

NOR2xp33_ASAP7_75t_R g4682 ( 
.A(n_4639),
.B(n_4482),
.Y(n_4682)
);

NOR2xp33_ASAP7_75t_L g4683 ( 
.A(n_4573),
.B(n_2516),
.Y(n_4683)
);

AOI21xp5_ASAP7_75t_L g4684 ( 
.A1(n_4664),
.A2(n_2842),
.B(n_2838),
.Y(n_4684)
);

NOR3xp33_ASAP7_75t_L g4685 ( 
.A(n_4550),
.B(n_2848),
.C(n_2847),
.Y(n_4685)
);

AOI21xp5_ASAP7_75t_L g4686 ( 
.A1(n_4417),
.A2(n_4553),
.B(n_4526),
.Y(n_4686)
);

AOI21xp5_ASAP7_75t_L g4687 ( 
.A1(n_4388),
.A2(n_2857),
.B(n_2854),
.Y(n_4687)
);

AOI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4585),
.A2(n_2865),
.B(n_2582),
.Y(n_4688)
);

NOR2xp33_ASAP7_75t_L g4689 ( 
.A(n_4375),
.B(n_2517),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4518),
.B(n_2519),
.Y(n_4690)
);

NOR3xp33_ASAP7_75t_L g4691 ( 
.A(n_4541),
.B(n_2600),
.C(n_2562),
.Y(n_4691)
);

OR2x6_ASAP7_75t_L g4692 ( 
.A(n_4374),
.B(n_2618),
.Y(n_4692)
);

OAI21xp33_ASAP7_75t_L g4693 ( 
.A1(n_4436),
.A2(n_2524),
.B(n_2520),
.Y(n_4693)
);

NAND2xp5_ASAP7_75t_SL g4694 ( 
.A(n_4582),
.B(n_2525),
.Y(n_4694)
);

AND2x4_ASAP7_75t_L g4695 ( 
.A(n_4666),
.B(n_2660),
.Y(n_4695)
);

AOI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4551),
.A2(n_4655),
.B(n_4407),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_SL g4697 ( 
.A(n_4399),
.B(n_2526),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_L g4698 ( 
.A(n_4463),
.B(n_4450),
.Y(n_4698)
);

OAI21xp5_ASAP7_75t_L g4699 ( 
.A1(n_4439),
.A2(n_2743),
.B(n_2695),
.Y(n_4699)
);

AOI21xp5_ASAP7_75t_L g4700 ( 
.A1(n_4527),
.A2(n_2752),
.B(n_2749),
.Y(n_4700)
);

OAI21x1_ASAP7_75t_L g4701 ( 
.A1(n_4534),
.A2(n_2795),
.B(n_2789),
.Y(n_4701)
);

NAND2xp5_ASAP7_75t_L g4702 ( 
.A(n_4432),
.B(n_2527),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4533),
.Y(n_4703)
);

INVx2_ASAP7_75t_L g4704 ( 
.A(n_4377),
.Y(n_4704)
);

BUFx3_ASAP7_75t_L g4705 ( 
.A(n_4443),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_SL g4706 ( 
.A(n_4525),
.B(n_2528),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4507),
.B(n_2529),
.Y(n_4707)
);

OAI21xp5_ASAP7_75t_L g4708 ( 
.A1(n_4488),
.A2(n_2830),
.B(n_2815),
.Y(n_4708)
);

BUFx6f_ASAP7_75t_L g4709 ( 
.A(n_4443),
.Y(n_4709)
);

NOR2xp33_ASAP7_75t_L g4710 ( 
.A(n_4613),
.B(n_2531),
.Y(n_4710)
);

AOI21xp5_ASAP7_75t_L g4711 ( 
.A1(n_4618),
.A2(n_2536),
.B(n_2533),
.Y(n_4711)
);

NOR2x2_ASAP7_75t_L g4712 ( 
.A(n_4559),
.B(n_2539),
.Y(n_4712)
);

A2O1A1Ixp33_ASAP7_75t_L g4713 ( 
.A1(n_4501),
.A2(n_2543),
.B(n_2544),
.C(n_2541),
.Y(n_4713)
);

AND2x2_ASAP7_75t_L g4714 ( 
.A(n_4477),
.B(n_2545),
.Y(n_4714)
);

INVx1_ASAP7_75t_L g4715 ( 
.A(n_4380),
.Y(n_4715)
);

AO21x1_ASAP7_75t_L g4716 ( 
.A1(n_4440),
.A2(n_4),
.B(n_5),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4391),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4503),
.B(n_4409),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4409),
.B(n_2547),
.Y(n_4719)
);

OAI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_4580),
.A2(n_2549),
.B(n_2548),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_SL g4721 ( 
.A(n_4525),
.B(n_2552),
.Y(n_4721)
);

AOI21xp5_ASAP7_75t_L g4722 ( 
.A1(n_4494),
.A2(n_2555),
.B(n_2554),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4409),
.B(n_2558),
.Y(n_4723)
);

AND2x2_ASAP7_75t_L g4724 ( 
.A(n_4589),
.B(n_2559),
.Y(n_4724)
);

OAI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4593),
.A2(n_2561),
.B(n_2560),
.Y(n_4725)
);

AOI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_4426),
.A2(n_2567),
.B(n_2566),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4458),
.B(n_2568),
.Y(n_4727)
);

NOR2xp67_ASAP7_75t_L g4728 ( 
.A(n_4621),
.B(n_1829),
.Y(n_4728)
);

INVx3_ASAP7_75t_L g4729 ( 
.A(n_4402),
.Y(n_4729)
);

AOI21xp5_ASAP7_75t_L g4730 ( 
.A1(n_4393),
.A2(n_2571),
.B(n_2569),
.Y(n_4730)
);

AND2x6_ASAP7_75t_L g4731 ( 
.A(n_4658),
.B(n_1830),
.Y(n_4731)
);

NOR2xp67_ASAP7_75t_L g4732 ( 
.A(n_4665),
.B(n_4466),
.Y(n_4732)
);

INVx3_ASAP7_75t_L g4733 ( 
.A(n_4402),
.Y(n_4733)
);

AO21x1_ASAP7_75t_L g4734 ( 
.A1(n_4557),
.A2(n_5),
.B(n_6),
.Y(n_4734)
);

INVxp67_ASAP7_75t_L g4735 ( 
.A(n_4529),
.Y(n_4735)
);

AOI21xp5_ASAP7_75t_L g4736 ( 
.A1(n_4398),
.A2(n_2573),
.B(n_2572),
.Y(n_4736)
);

NAND2xp5_ASAP7_75t_L g4737 ( 
.A(n_4495),
.B(n_2574),
.Y(n_4737)
);

NOR2x1p5_ASAP7_75t_SL g4738 ( 
.A(n_4525),
.B(n_1831),
.Y(n_4738)
);

AOI22xp5_ASAP7_75t_L g4739 ( 
.A1(n_4563),
.A2(n_2578),
.B1(n_2579),
.B2(n_2575),
.Y(n_4739)
);

O2A1O1Ixp33_ASAP7_75t_L g4740 ( 
.A1(n_4546),
.A2(n_2581),
.B(n_2585),
.C(n_2580),
.Y(n_4740)
);

AOI21xp5_ASAP7_75t_L g4741 ( 
.A1(n_4403),
.A2(n_2588),
.B(n_2587),
.Y(n_4741)
);

AOI21xp5_ASAP7_75t_L g4742 ( 
.A1(n_4428),
.A2(n_2593),
.B(n_2591),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_L g4743 ( 
.A(n_4555),
.B(n_2595),
.Y(n_4743)
);

NOR2xp67_ASAP7_75t_L g4744 ( 
.A(n_4617),
.B(n_4480),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_SL g4745 ( 
.A(n_4525),
.B(n_2604),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4561),
.B(n_2605),
.Y(n_4746)
);

NAND2xp5_ASAP7_75t_L g4747 ( 
.A(n_4435),
.B(n_4433),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_4437),
.A2(n_2610),
.B(n_2606),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4445),
.Y(n_4749)
);

AOI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_4447),
.A2(n_2612),
.B(n_2611),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4459),
.B(n_4472),
.Y(n_4751)
);

AND2x2_ASAP7_75t_SL g4752 ( 
.A(n_4412),
.B(n_7),
.Y(n_4752)
);

BUFx4f_ASAP7_75t_L g4753 ( 
.A(n_4374),
.Y(n_4753)
);

O2A1O1Ixp33_ASAP7_75t_L g4754 ( 
.A1(n_4449),
.A2(n_2615),
.B(n_2619),
.C(n_2613),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4475),
.B(n_2620),
.Y(n_4755)
);

AOI22xp33_ASAP7_75t_L g4756 ( 
.A1(n_4572),
.A2(n_2625),
.B1(n_2626),
.B2(n_2624),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_4401),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4476),
.B(n_2627),
.Y(n_4758)
);

BUFx6f_ASAP7_75t_L g4759 ( 
.A(n_4423),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_SL g4760 ( 
.A(n_4415),
.B(n_4661),
.Y(n_4760)
);

AOI21xp5_ASAP7_75t_L g4761 ( 
.A1(n_4493),
.A2(n_2634),
.B(n_2632),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4520),
.B(n_2637),
.Y(n_4762)
);

NAND2xp5_ASAP7_75t_L g4763 ( 
.A(n_4530),
.B(n_2638),
.Y(n_4763)
);

INVx2_ASAP7_75t_L g4764 ( 
.A(n_4410),
.Y(n_4764)
);

AND2x4_ASAP7_75t_L g4765 ( 
.A(n_4452),
.B(n_2639),
.Y(n_4765)
);

OAI22xp5_ASAP7_75t_L g4766 ( 
.A1(n_4397),
.A2(n_2645),
.B1(n_2646),
.B2(n_2640),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4568),
.B(n_2649),
.Y(n_4767)
);

INVx4_ASAP7_75t_L g4768 ( 
.A(n_4423),
.Y(n_4768)
);

AOI21xp5_ASAP7_75t_L g4769 ( 
.A1(n_4536),
.A2(n_2651),
.B(n_2650),
.Y(n_4769)
);

NAND2xp5_ASAP7_75t_L g4770 ( 
.A(n_4659),
.B(n_2652),
.Y(n_4770)
);

AOI21xp5_ASAP7_75t_L g4771 ( 
.A1(n_4660),
.A2(n_2656),
.B(n_2653),
.Y(n_4771)
);

BUFx6f_ASAP7_75t_L g4772 ( 
.A(n_4492),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4395),
.B(n_2657),
.Y(n_4773)
);

CKINVDCx5p33_ASAP7_75t_R g4774 ( 
.A(n_4455),
.Y(n_4774)
);

AOI21xp5_ASAP7_75t_L g4775 ( 
.A1(n_4505),
.A2(n_2661),
.B(n_2658),
.Y(n_4775)
);

NAND2xp5_ASAP7_75t_L g4776 ( 
.A(n_4567),
.B(n_2663),
.Y(n_4776)
);

NOR2x1_ASAP7_75t_L g4777 ( 
.A(n_4382),
.B(n_2664),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4570),
.B(n_4548),
.Y(n_4778)
);

BUFx6f_ASAP7_75t_L g4779 ( 
.A(n_4492),
.Y(n_4779)
);

AOI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4496),
.A2(n_2669),
.B(n_2667),
.Y(n_4780)
);

INVx4_ASAP7_75t_L g4781 ( 
.A(n_4400),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4394),
.B(n_2670),
.Y(n_4782)
);

INVx4_ASAP7_75t_L g4783 ( 
.A(n_4400),
.Y(n_4783)
);

BUFx4f_ASAP7_75t_L g4784 ( 
.A(n_4404),
.Y(n_4784)
);

CKINVDCx5p33_ASAP7_75t_R g4785 ( 
.A(n_4456),
.Y(n_4785)
);

O2A1O1Ixp33_ASAP7_75t_L g4786 ( 
.A1(n_4498),
.A2(n_2672),
.B(n_2674),
.C(n_2671),
.Y(n_4786)
);

AOI22xp33_ASAP7_75t_L g4787 ( 
.A1(n_4512),
.A2(n_2682),
.B1(n_2684),
.B2(n_2678),
.Y(n_4787)
);

O2A1O1Ixp33_ASAP7_75t_L g4788 ( 
.A1(n_4389),
.A2(n_2686),
.B(n_2690),
.C(n_2685),
.Y(n_4788)
);

OAI21xp5_ASAP7_75t_L g4789 ( 
.A1(n_4390),
.A2(n_2693),
.B(n_2692),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4486),
.B(n_2697),
.Y(n_4790)
);

INVx3_ASAP7_75t_L g4791 ( 
.A(n_4577),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4430),
.Y(n_4792)
);

AOI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_4656),
.A2(n_2706),
.B(n_2701),
.Y(n_4793)
);

INVxp67_ASAP7_75t_L g4794 ( 
.A(n_4425),
.Y(n_4794)
);

A2O1A1Ixp33_ASAP7_75t_L g4795 ( 
.A1(n_4535),
.A2(n_2712),
.B(n_2713),
.C(n_2709),
.Y(n_4795)
);

BUFx6f_ASAP7_75t_L g4796 ( 
.A(n_4577),
.Y(n_4796)
);

AND2x4_ASAP7_75t_L g4797 ( 
.A(n_4489),
.B(n_2715),
.Y(n_4797)
);

OAI21xp33_ASAP7_75t_L g4798 ( 
.A1(n_4427),
.A2(n_2719),
.B(n_2718),
.Y(n_4798)
);

INVx1_ASAP7_75t_SL g4799 ( 
.A(n_4504),
.Y(n_4799)
);

NAND2xp5_ASAP7_75t_SL g4800 ( 
.A(n_4547),
.B(n_2720),
.Y(n_4800)
);

INVx1_ASAP7_75t_L g4801 ( 
.A(n_4571),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_4446),
.Y(n_4802)
);

NOR2xp33_ASAP7_75t_L g4803 ( 
.A(n_4654),
.B(n_2722),
.Y(n_4803)
);

A2O1A1Ixp33_ASAP7_75t_L g4804 ( 
.A1(n_4424),
.A2(n_2725),
.B(n_2728),
.C(n_2724),
.Y(n_4804)
);

OAI21xp5_ASAP7_75t_L g4805 ( 
.A1(n_4392),
.A2(n_2734),
.B(n_2731),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4623),
.B(n_2735),
.Y(n_4806)
);

AOI22xp33_ASAP7_75t_L g4807 ( 
.A1(n_4554),
.A2(n_2742),
.B1(n_2745),
.B2(n_2741),
.Y(n_4807)
);

AOI21xp5_ASAP7_75t_L g4808 ( 
.A1(n_4429),
.A2(n_4434),
.B(n_4565),
.Y(n_4808)
);

OAI21xp5_ASAP7_75t_L g4809 ( 
.A1(n_4616),
.A2(n_2750),
.B(n_2747),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4574),
.Y(n_4810)
);

NAND2xp5_ASAP7_75t_L g4811 ( 
.A(n_4451),
.B(n_2756),
.Y(n_4811)
);

CKINVDCx5p33_ASAP7_75t_R g4812 ( 
.A(n_4508),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_L g4813 ( 
.A(n_4461),
.B(n_2759),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_L g4814 ( 
.A(n_4465),
.B(n_2760),
.Y(n_4814)
);

BUFx12f_ASAP7_75t_L g4815 ( 
.A(n_4594),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4576),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4474),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4487),
.B(n_2761),
.Y(n_4818)
);

INVx4_ASAP7_75t_L g4819 ( 
.A(n_4540),
.Y(n_4819)
);

OAI21xp5_ASAP7_75t_L g4820 ( 
.A1(n_4620),
.A2(n_2763),
.B(n_2762),
.Y(n_4820)
);

INVx3_ASAP7_75t_L g4821 ( 
.A(n_4590),
.Y(n_4821)
);

NAND2xp5_ASAP7_75t_L g4822 ( 
.A(n_4513),
.B(n_4514),
.Y(n_4822)
);

AO22x1_ASAP7_75t_L g4823 ( 
.A1(n_4609),
.A2(n_2770),
.B1(n_2771),
.B2(n_2765),
.Y(n_4823)
);

AOI21xp33_ASAP7_75t_L g4824 ( 
.A1(n_4491),
.A2(n_2775),
.B(n_2772),
.Y(n_4824)
);

AND2x4_ASAP7_75t_L g4825 ( 
.A(n_4510),
.B(n_2777),
.Y(n_4825)
);

NAND2xp33_ASAP7_75t_L g4826 ( 
.A(n_4441),
.B(n_2780),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4614),
.A2(n_2784),
.B(n_2781),
.Y(n_4827)
);

NAND2xp5_ASAP7_75t_L g4828 ( 
.A(n_4524),
.B(n_2785),
.Y(n_4828)
);

AOI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_4612),
.A2(n_2790),
.B(n_2786),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4538),
.B(n_2794),
.Y(n_4830)
);

AOI21xp5_ASAP7_75t_L g4831 ( 
.A1(n_4631),
.A2(n_4635),
.B(n_4646),
.Y(n_4831)
);

BUFx3_ASAP7_75t_L g4832 ( 
.A(n_4383),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4490),
.B(n_2797),
.Y(n_4833)
);

OAI321xp33_ASAP7_75t_L g4834 ( 
.A1(n_4531),
.A2(n_2807),
.A3(n_2804),
.B1(n_2808),
.B2(n_2806),
.C(n_2799),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4556),
.Y(n_4835)
);

INVx4_ASAP7_75t_L g4836 ( 
.A(n_4559),
.Y(n_4836)
);

NOR2xp33_ASAP7_75t_R g4837 ( 
.A(n_4497),
.B(n_4545),
.Y(n_4837)
);

AOI22xp33_ASAP7_75t_L g4838 ( 
.A1(n_4652),
.A2(n_4633),
.B1(n_4651),
.B2(n_4626),
.Y(n_4838)
);

AOI21xp5_ASAP7_75t_L g4839 ( 
.A1(n_4464),
.A2(n_2810),
.B(n_2809),
.Y(n_4839)
);

AOI21xp5_ASAP7_75t_L g4840 ( 
.A1(n_4442),
.A2(n_2812),
.B(n_2811),
.Y(n_4840)
);

OR2x2_ASAP7_75t_L g4841 ( 
.A(n_4578),
.B(n_2813),
.Y(n_4841)
);

O2A1O1Ixp33_ASAP7_75t_L g4842 ( 
.A1(n_4453),
.A2(n_2822),
.B(n_2823),
.C(n_2821),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4408),
.B(n_2825),
.Y(n_4843)
);

NOR2xp33_ASAP7_75t_L g4844 ( 
.A(n_4532),
.B(n_2832),
.Y(n_4844)
);

AND2x4_ASAP7_75t_L g4845 ( 
.A(n_4376),
.B(n_2834),
.Y(n_4845)
);

AOI21xp5_ASAP7_75t_L g4846 ( 
.A1(n_4444),
.A2(n_2840),
.B(n_2836),
.Y(n_4846)
);

AOI21x1_ASAP7_75t_L g4847 ( 
.A1(n_4606),
.A2(n_1833),
.B(n_1832),
.Y(n_4847)
);

INVx2_ASAP7_75t_L g4848 ( 
.A(n_4581),
.Y(n_4848)
);

AND2x2_ASAP7_75t_L g4849 ( 
.A(n_4431),
.B(n_2844),
.Y(n_4849)
);

AOI21xp5_ASAP7_75t_L g4850 ( 
.A1(n_4454),
.A2(n_2846),
.B(n_2845),
.Y(n_4850)
);

INVx3_ASAP7_75t_L g4851 ( 
.A(n_4645),
.Y(n_4851)
);

AOI21xp5_ASAP7_75t_L g4852 ( 
.A1(n_4381),
.A2(n_2851),
.B(n_2849),
.Y(n_4852)
);

AOI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4405),
.A2(n_2859),
.B(n_2852),
.Y(n_4853)
);

INVx6_ASAP7_75t_L g4854 ( 
.A(n_4629),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_4653),
.B(n_2862),
.Y(n_4855)
);

INVx3_ASAP7_75t_L g4856 ( 
.A(n_4645),
.Y(n_4856)
);

NAND2xp5_ASAP7_75t_SL g4857 ( 
.A(n_4506),
.B(n_2866),
.Y(n_4857)
);

INVxp67_ASAP7_75t_L g4858 ( 
.A(n_4416),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4411),
.A2(n_4420),
.B(n_4413),
.Y(n_4859)
);

NOR2xp33_ASAP7_75t_L g4860 ( 
.A(n_4539),
.B(n_2868),
.Y(n_4860)
);

BUFx10_ASAP7_75t_L g4861 ( 
.A(n_4595),
.Y(n_4861)
);

AOI21xp5_ASAP7_75t_L g4862 ( 
.A1(n_4421),
.A2(n_1835),
.B(n_1834),
.Y(n_4862)
);

O2A1O1Ixp33_ASAP7_75t_L g4863 ( 
.A1(n_4473),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_4863)
);

NAND2xp5_ASAP7_75t_L g4864 ( 
.A(n_4642),
.B(n_9),
.Y(n_4864)
);

AOI21x1_ASAP7_75t_L g4865 ( 
.A1(n_4619),
.A2(n_1838),
.B(n_1836),
.Y(n_4865)
);

NOR2xp33_ASAP7_75t_L g4866 ( 
.A(n_4634),
.B(n_10),
.Y(n_4866)
);

OAI22xp5_ASAP7_75t_L g4867 ( 
.A1(n_4462),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_SL g4868 ( 
.A(n_4624),
.B(n_11),
.Y(n_4868)
);

AND2x4_ASAP7_75t_L g4869 ( 
.A(n_4630),
.B(n_1841),
.Y(n_4869)
);

INVx1_ASAP7_75t_SL g4870 ( 
.A(n_4481),
.Y(n_4870)
);

AOI21xp5_ASAP7_75t_L g4871 ( 
.A1(n_4422),
.A2(n_1848),
.B(n_1842),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4601),
.B(n_12),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4615),
.B(n_13),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4650),
.B(n_13),
.Y(n_4874)
);

O2A1O1Ixp5_ASAP7_75t_L g4875 ( 
.A1(n_4586),
.A2(n_16),
.B(n_14),
.C(n_15),
.Y(n_4875)
);

AOI21xp5_ASAP7_75t_L g4876 ( 
.A1(n_4470),
.A2(n_1859),
.B(n_1854),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_SL g4877 ( 
.A(n_4629),
.B(n_14),
.Y(n_4877)
);

AOI21xp5_ASAP7_75t_L g4878 ( 
.A1(n_4478),
.A2(n_1862),
.B(n_1861),
.Y(n_4878)
);

INVx4_ASAP7_75t_L g4879 ( 
.A(n_4629),
.Y(n_4879)
);

AOI22xp5_ASAP7_75t_L g4880 ( 
.A1(n_4607),
.A2(n_4502),
.B1(n_4467),
.B2(n_4418),
.Y(n_4880)
);

INVx2_ASAP7_75t_L g4881 ( 
.A(n_4562),
.Y(n_4881)
);

AOI21xp5_ASAP7_75t_L g4882 ( 
.A1(n_4479),
.A2(n_1864),
.B(n_1863),
.Y(n_4882)
);

A2O1A1Ixp33_ASAP7_75t_L g4883 ( 
.A1(n_4448),
.A2(n_17),
.B(n_15),
.C(n_16),
.Y(n_4883)
);

INVxp67_ASAP7_75t_L g4884 ( 
.A(n_4406),
.Y(n_4884)
);

NOR2xp67_ASAP7_75t_L g4885 ( 
.A(n_4657),
.B(n_1865),
.Y(n_4885)
);

NOR2xp33_ASAP7_75t_L g4886 ( 
.A(n_4484),
.B(n_4457),
.Y(n_4886)
);

NAND2x1p5_ASAP7_75t_L g4887 ( 
.A(n_4564),
.B(n_1866),
.Y(n_4887)
);

OR2x2_ASAP7_75t_SL g4888 ( 
.A(n_4483),
.B(n_17),
.Y(n_4888)
);

AOI21x1_ASAP7_75t_L g4889 ( 
.A1(n_4522),
.A2(n_1871),
.B(n_1868),
.Y(n_4889)
);

BUFx2_ASAP7_75t_L g4890 ( 
.A(n_4598),
.Y(n_4890)
);

OAI22xp5_ASAP7_75t_L g4891 ( 
.A1(n_4414),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_4891)
);

NAND2xp5_ASAP7_75t_L g4892 ( 
.A(n_4632),
.B(n_4636),
.Y(n_4892)
);

INVx2_ASAP7_75t_SL g4893 ( 
.A(n_4592),
.Y(n_4893)
);

BUFx6f_ASAP7_75t_L g4894 ( 
.A(n_4566),
.Y(n_4894)
);

OR2x2_ASAP7_75t_L g4895 ( 
.A(n_4485),
.B(n_18),
.Y(n_4895)
);

INVx2_ASAP7_75t_SL g4896 ( 
.A(n_4575),
.Y(n_4896)
);

O2A1O1Ixp5_ASAP7_75t_L g4897 ( 
.A1(n_4468),
.A2(n_22),
.B(n_19),
.C(n_21),
.Y(n_4897)
);

BUFx6f_ASAP7_75t_L g4898 ( 
.A(n_4597),
.Y(n_4898)
);

AOI21x1_ASAP7_75t_L g4899 ( 
.A1(n_4560),
.A2(n_1874),
.B(n_1873),
.Y(n_4899)
);

NOR2xp33_ASAP7_75t_L g4900 ( 
.A(n_4627),
.B(n_21),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4647),
.B(n_24),
.Y(n_4901)
);

CKINVDCx20_ASAP7_75t_R g4902 ( 
.A(n_4469),
.Y(n_4902)
);

AOI21xp5_ASAP7_75t_L g4903 ( 
.A1(n_4499),
.A2(n_1882),
.B(n_1877),
.Y(n_4903)
);

NAND2xp5_ASAP7_75t_L g4904 ( 
.A(n_4603),
.B(n_24),
.Y(n_4904)
);

INVx2_ASAP7_75t_L g4905 ( 
.A(n_4605),
.Y(n_4905)
);

HB1xp67_ASAP7_75t_L g4906 ( 
.A(n_4610),
.Y(n_4906)
);

INVx4_ASAP7_75t_L g4907 ( 
.A(n_4628),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4638),
.Y(n_4908)
);

AOI21xp5_ASAP7_75t_L g4909 ( 
.A1(n_4500),
.A2(n_25),
.B(n_27),
.Y(n_4909)
);

OAI21xp5_ASAP7_75t_L g4910 ( 
.A1(n_4509),
.A2(n_29),
.B(n_30),
.Y(n_4910)
);

INVx1_ASAP7_75t_L g4911 ( 
.A(n_4643),
.Y(n_4911)
);

NAND2x1_ASAP7_75t_L g4912 ( 
.A(n_4599),
.B(n_29),
.Y(n_4912)
);

NOR2xp33_ASAP7_75t_L g4913 ( 
.A(n_4544),
.B(n_30),
.Y(n_4913)
);

A2O1A1Ixp33_ASAP7_75t_L g4914 ( 
.A1(n_4549),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4637),
.Y(n_4915)
);

NOR2xp33_ASAP7_75t_L g4916 ( 
.A(n_4515),
.B(n_31),
.Y(n_4916)
);

AOI21xp5_ASAP7_75t_L g4917 ( 
.A1(n_4516),
.A2(n_32),
.B(n_33),
.Y(n_4917)
);

NAND2x1_ASAP7_75t_L g4918 ( 
.A(n_4600),
.B(n_4602),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4521),
.B(n_34),
.Y(n_4919)
);

AOI22xp5_ASAP7_75t_L g4920 ( 
.A1(n_4596),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_SL g4921 ( 
.A(n_4523),
.B(n_35),
.Y(n_4921)
);

INVx3_ASAP7_75t_L g4922 ( 
.A(n_4604),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_L g4923 ( 
.A(n_4471),
.B(n_37),
.Y(n_4923)
);

OAI21xp33_ASAP7_75t_L g4924 ( 
.A1(n_4552),
.A2(n_37),
.B(n_38),
.Y(n_4924)
);

AOI21x1_ASAP7_75t_L g4925 ( 
.A1(n_4649),
.A2(n_38),
.B(n_39),
.Y(n_4925)
);

AOI22xp33_ASAP7_75t_L g4926 ( 
.A1(n_4608),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_4926)
);

OR2x6_ASAP7_75t_L g4927 ( 
.A(n_4558),
.B(n_40),
.Y(n_4927)
);

BUFx2_ASAP7_75t_L g4928 ( 
.A(n_4569),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_SL g4929 ( 
.A(n_4579),
.B(n_4583),
.Y(n_4929)
);

OAI21xp5_ASAP7_75t_L g4930 ( 
.A1(n_4584),
.A2(n_41),
.B(n_43),
.Y(n_4930)
);

OAI22xp5_ASAP7_75t_L g4931 ( 
.A1(n_4672),
.A2(n_4588),
.B1(n_4587),
.B2(n_4611),
.Y(n_4931)
);

A2O1A1Ixp33_ASAP7_75t_L g4932 ( 
.A1(n_4678),
.A2(n_4625),
.B(n_4640),
.C(n_4622),
.Y(n_4932)
);

AND2x4_ASAP7_75t_L g4933 ( 
.A(n_4705),
.B(n_4644),
.Y(n_4933)
);

AOI21xp5_ASAP7_75t_L g4934 ( 
.A1(n_4667),
.A2(n_4648),
.B(n_43),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_SL g4935 ( 
.A(n_4686),
.B(n_44),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4668),
.B(n_44),
.Y(n_4936)
);

O2A1O1Ixp5_ASAP7_75t_L g4937 ( 
.A1(n_4910),
.A2(n_4930),
.B(n_4918),
.C(n_4900),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4675),
.A2(n_45),
.B(n_46),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4747),
.B(n_45),
.Y(n_4939)
);

NAND3xp33_ASAP7_75t_L g4940 ( 
.A(n_4913),
.B(n_47),
.C(n_48),
.Y(n_4940)
);

O2A1O1Ixp33_ASAP7_75t_SL g4941 ( 
.A1(n_4914),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_4941)
);

BUFx3_ASAP7_75t_L g4942 ( 
.A(n_4709),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_L g4943 ( 
.A(n_4799),
.B(n_49),
.Y(n_4943)
);

AOI21xp5_ASAP7_75t_L g4944 ( 
.A1(n_4859),
.A2(n_50),
.B(n_51),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_L g4945 ( 
.A(n_4928),
.B(n_50),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_SL g4946 ( 
.A(n_4718),
.B(n_52),
.Y(n_4946)
);

HB1xp67_ASAP7_75t_L g4947 ( 
.A(n_4735),
.Y(n_4947)
);

OAI22xp5_ASAP7_75t_L g4948 ( 
.A1(n_4676),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_4948)
);

OAI22xp5_ASAP7_75t_L g4949 ( 
.A1(n_4866),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_4949)
);

BUFx4f_ASAP7_75t_L g4950 ( 
.A(n_4815),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4890),
.B(n_55),
.Y(n_4951)
);

BUFx10_ASAP7_75t_L g4952 ( 
.A(n_4785),
.Y(n_4952)
);

OAI22xp5_ASAP7_75t_L g4953 ( 
.A1(n_4916),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_4953)
);

AOI21xp5_ASAP7_75t_L g4954 ( 
.A1(n_4808),
.A2(n_56),
.B(n_57),
.Y(n_4954)
);

AOI21xp5_ASAP7_75t_L g4955 ( 
.A1(n_4706),
.A2(n_58),
.B(n_59),
.Y(n_4955)
);

O2A1O1Ixp33_ASAP7_75t_SL g4956 ( 
.A1(n_4883),
.A2(n_4867),
.B(n_4745),
.C(n_4721),
.Y(n_4956)
);

NOR2xp33_ASAP7_75t_SL g4957 ( 
.A(n_4753),
.B(n_60),
.Y(n_4957)
);

INVx2_ASAP7_75t_L g4958 ( 
.A(n_4704),
.Y(n_4958)
);

AOI22xp33_ASAP7_75t_L g4959 ( 
.A1(n_4685),
.A2(n_62),
.B1(n_60),
.B2(n_61),
.Y(n_4959)
);

AOI21xp5_ASAP7_75t_L g4960 ( 
.A1(n_4929),
.A2(n_61),
.B(n_63),
.Y(n_4960)
);

A2O1A1Ixp33_ASAP7_75t_L g4961 ( 
.A1(n_4693),
.A2(n_65),
.B(n_63),
.C(n_64),
.Y(n_4961)
);

OA22x2_ASAP7_75t_L g4962 ( 
.A1(n_4880),
.A2(n_68),
.B1(n_65),
.B2(n_67),
.Y(n_4962)
);

NOR2xp33_ASAP7_75t_L g4963 ( 
.A(n_4710),
.B(n_69),
.Y(n_4963)
);

AOI21x1_ASAP7_75t_L g4964 ( 
.A1(n_4673),
.A2(n_4899),
.B(n_4696),
.Y(n_4964)
);

A2O1A1Ixp33_ASAP7_75t_L g4965 ( 
.A1(n_4886),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_4965)
);

NAND2xp5_ASAP7_75t_L g4966 ( 
.A(n_4915),
.B(n_70),
.Y(n_4966)
);

NAND2xp5_ASAP7_75t_L g4967 ( 
.A(n_4794),
.B(n_71),
.Y(n_4967)
);

INVx2_ASAP7_75t_L g4968 ( 
.A(n_4717),
.Y(n_4968)
);

BUFx6f_ASAP7_75t_L g4969 ( 
.A(n_4709),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4751),
.Y(n_4970)
);

INVx3_ASAP7_75t_L g4971 ( 
.A(n_4759),
.Y(n_4971)
);

AOI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_4831),
.A2(n_72),
.B(n_73),
.Y(n_4972)
);

OAI22xp5_ASAP7_75t_L g4973 ( 
.A1(n_4923),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_4973)
);

NOR2xp33_ASAP7_75t_L g4974 ( 
.A(n_4803),
.B(n_74),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_SL g4975 ( 
.A(n_4922),
.B(n_75),
.Y(n_4975)
);

NAND2xp5_ASAP7_75t_L g4976 ( 
.A(n_4698),
.B(n_76),
.Y(n_4976)
);

OAI22xp5_ASAP7_75t_L g4977 ( 
.A1(n_4919),
.A2(n_78),
.B1(n_76),
.B2(n_77),
.Y(n_4977)
);

NOR2xp33_ASAP7_75t_SL g4978 ( 
.A(n_4784),
.B(n_77),
.Y(n_4978)
);

HB1xp67_ASAP7_75t_L g4979 ( 
.A(n_4778),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4862),
.A2(n_80),
.B(n_81),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_SL g4981 ( 
.A(n_4861),
.B(n_81),
.Y(n_4981)
);

O2A1O1Ixp5_ASAP7_75t_L g4982 ( 
.A1(n_4670),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4724),
.B(n_83),
.Y(n_4983)
);

NAND2xp5_ASAP7_75t_SL g4984 ( 
.A(n_4851),
.B(n_84),
.Y(n_4984)
);

AOI22xp5_ASAP7_75t_L g4985 ( 
.A1(n_4683),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_4985)
);

INVx1_ASAP7_75t_L g4986 ( 
.A(n_4848),
.Y(n_4986)
);

A2O1A1Ixp33_ASAP7_75t_L g4987 ( 
.A1(n_4924),
.A2(n_87),
.B(n_85),
.C(n_86),
.Y(n_4987)
);

OAI22xp5_ASAP7_75t_L g4988 ( 
.A1(n_4927),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4715),
.B(n_88),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_SL g4990 ( 
.A(n_4856),
.B(n_90),
.Y(n_4990)
);

AOI22xp33_ASAP7_75t_L g4991 ( 
.A1(n_4838),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_4991)
);

AOI21xp5_ASAP7_75t_L g4992 ( 
.A1(n_4871),
.A2(n_4878),
.B(n_4876),
.Y(n_4992)
);

AOI21xp5_ASAP7_75t_L g4993 ( 
.A1(n_4882),
.A2(n_92),
.B(n_93),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4903),
.A2(n_94),
.B(n_95),
.Y(n_4994)
);

AOI21xp5_ASAP7_75t_L g4995 ( 
.A1(n_4826),
.A2(n_94),
.B(n_95),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4703),
.Y(n_4996)
);

BUFx3_ASAP7_75t_L g4997 ( 
.A(n_4796),
.Y(n_4997)
);

AOI21xp5_ASAP7_75t_L g4998 ( 
.A1(n_4864),
.A2(n_96),
.B(n_97),
.Y(n_4998)
);

AOI33xp33_ASAP7_75t_L g4999 ( 
.A1(n_4756),
.A2(n_98),
.A3(n_101),
.B1(n_96),
.B2(n_97),
.B3(n_100),
.Y(n_4999)
);

BUFx3_ASAP7_75t_L g5000 ( 
.A(n_4796),
.Y(n_5000)
);

INVxp67_ASAP7_75t_L g5001 ( 
.A(n_4870),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4749),
.Y(n_5002)
);

INVx1_ASAP7_75t_SL g5003 ( 
.A(n_4682),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4701),
.A2(n_100),
.B(n_101),
.Y(n_5004)
);

INVxp67_ASAP7_75t_L g5005 ( 
.A(n_4759),
.Y(n_5005)
);

NAND2xp5_ASAP7_75t_SL g5006 ( 
.A(n_4732),
.B(n_102),
.Y(n_5006)
);

AOI21xp5_ASAP7_75t_L g5007 ( 
.A1(n_4872),
.A2(n_102),
.B(n_103),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_SL g5008 ( 
.A(n_4834),
.B(n_103),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4801),
.B(n_104),
.Y(n_5009)
);

OAI22xp5_ASAP7_75t_L g5010 ( 
.A1(n_4927),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4810),
.B(n_4816),
.Y(n_5011)
);

AOI21x1_ASAP7_75t_L g5012 ( 
.A1(n_4671),
.A2(n_105),
.B(n_106),
.Y(n_5012)
);

AOI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_4873),
.A2(n_107),
.B(n_109),
.Y(n_5013)
);

O2A1O1Ixp33_ASAP7_75t_L g5014 ( 
.A1(n_4824),
.A2(n_4720),
.B(n_4725),
.C(n_4809),
.Y(n_5014)
);

AND2x2_ASAP7_75t_L g5015 ( 
.A(n_4690),
.B(n_4681),
.Y(n_5015)
);

INVx2_ASAP7_75t_L g5016 ( 
.A(n_4757),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_L g5017 ( 
.A(n_4674),
.B(n_110),
.Y(n_5017)
);

NAND2xp5_ASAP7_75t_SL g5018 ( 
.A(n_4832),
.B(n_110),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4822),
.B(n_111),
.Y(n_5019)
);

NAND2x1p5_ASAP7_75t_L g5020 ( 
.A(n_4781),
.B(n_111),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4821),
.B(n_112),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4892),
.Y(n_5022)
);

NOR2x1_ASAP7_75t_L g5023 ( 
.A(n_4760),
.B(n_113),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4764),
.B(n_113),
.Y(n_5024)
);

AOI21x1_ASAP7_75t_L g5025 ( 
.A1(n_4889),
.A2(n_114),
.B(n_115),
.Y(n_5025)
);

NOR2xp33_ASAP7_75t_L g5026 ( 
.A(n_4884),
.B(n_114),
.Y(n_5026)
);

AOI21x1_ASAP7_75t_L g5027 ( 
.A1(n_4847),
.A2(n_115),
.B(n_116),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4792),
.B(n_116),
.Y(n_5028)
);

INVx5_ASAP7_75t_L g5029 ( 
.A(n_4731),
.Y(n_5029)
);

INVxp67_ASAP7_75t_SL g5030 ( 
.A(n_4906),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4874),
.A2(n_117),
.B(n_118),
.Y(n_5031)
);

O2A1O1Ixp5_ASAP7_75t_L g5032 ( 
.A1(n_4716),
.A2(n_121),
.B(n_119),
.C(n_120),
.Y(n_5032)
);

O2A1O1Ixp33_ASAP7_75t_L g5033 ( 
.A1(n_4820),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_5033)
);

NOR2xp33_ASAP7_75t_SL g5034 ( 
.A(n_4774),
.B(n_123),
.Y(n_5034)
);

HB1xp67_ASAP7_75t_L g5035 ( 
.A(n_4802),
.Y(n_5035)
);

AOI22xp5_ASAP7_75t_L g5036 ( 
.A1(n_4739),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_5036)
);

OAI22xp5_ASAP7_75t_L g5037 ( 
.A1(n_4920),
.A2(n_4895),
.B1(n_4926),
.B2(n_4833),
.Y(n_5037)
);

OR2x2_ASAP7_75t_SL g5038 ( 
.A(n_4854),
.B(n_4719),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4912),
.A2(n_125),
.B(n_126),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4817),
.B(n_127),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4835),
.B(n_127),
.Y(n_5041)
);

AOI33xp33_ASAP7_75t_L g5042 ( 
.A1(n_4807),
.A2(n_132),
.A3(n_134),
.B1(n_128),
.B2(n_131),
.B3(n_133),
.Y(n_5042)
);

AOI21xp5_ASAP7_75t_L g5043 ( 
.A1(n_4921),
.A2(n_4917),
.B(n_4909),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4908),
.Y(n_5044)
);

O2A1O1Ixp33_ASAP7_75t_L g5045 ( 
.A1(n_4677),
.A2(n_134),
.B(n_128),
.C(n_131),
.Y(n_5045)
);

AOI21xp5_ASAP7_75t_L g5046 ( 
.A1(n_4699),
.A2(n_135),
.B(n_136),
.Y(n_5046)
);

INVx1_ASAP7_75t_L g5047 ( 
.A(n_4911),
.Y(n_5047)
);

NAND2xp5_ASAP7_75t_L g5048 ( 
.A(n_4669),
.B(n_135),
.Y(n_5048)
);

OAI21xp5_ASAP7_75t_L g5049 ( 
.A1(n_4790),
.A2(n_136),
.B(n_137),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4836),
.B(n_137),
.Y(n_5050)
);

A2O1A1Ixp33_ASAP7_75t_L g5051 ( 
.A1(n_4754),
.A2(n_4786),
.B(n_4788),
.C(n_4700),
.Y(n_5051)
);

AND2x2_ASAP7_75t_SL g5052 ( 
.A(n_4752),
.B(n_138),
.Y(n_5052)
);

NOR2xp33_ASAP7_75t_L g5053 ( 
.A(n_4858),
.B(n_138),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_L g5054 ( 
.A1(n_4865),
.A2(n_140),
.B(n_141),
.Y(n_5054)
);

CKINVDCx20_ASAP7_75t_R g5055 ( 
.A(n_4812),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4783),
.B(n_140),
.Y(n_5056)
);

AOI21xp5_ASAP7_75t_L g5057 ( 
.A1(n_4789),
.A2(n_141),
.B(n_143),
.Y(n_5057)
);

NAND2x1p5_ASAP7_75t_L g5058 ( 
.A(n_4768),
.B(n_4879),
.Y(n_5058)
);

NOR2xp33_ASAP7_75t_L g5059 ( 
.A(n_4888),
.B(n_144),
.Y(n_5059)
);

BUFx2_ASAP7_75t_L g5060 ( 
.A(n_4729),
.Y(n_5060)
);

AOI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_4805),
.A2(n_144),
.B(n_145),
.Y(n_5061)
);

OAI22xp5_ASAP7_75t_L g5062 ( 
.A1(n_4713),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_5062)
);

NAND2x1p5_ASAP7_75t_L g5063 ( 
.A(n_4772),
.B(n_146),
.Y(n_5063)
);

AOI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_4680),
.A2(n_147),
.B(n_148),
.Y(n_5064)
);

AOI22xp5_ASAP7_75t_L g5065 ( 
.A1(n_4806),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_5065)
);

INVx2_ASAP7_75t_SL g5066 ( 
.A(n_4854),
.Y(n_5066)
);

OAI22xp5_ASAP7_75t_L g5067 ( 
.A1(n_4723),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_5067)
);

O2A1O1Ixp33_ASAP7_75t_L g5068 ( 
.A1(n_4740),
.A2(n_154),
.B(n_152),
.C(n_153),
.Y(n_5068)
);

AOI33xp33_ASAP7_75t_L g5069 ( 
.A1(n_4787),
.A2(n_154),
.A3(n_156),
.B1(n_152),
.B2(n_153),
.B3(n_155),
.Y(n_5069)
);

OAI21x1_ASAP7_75t_L g5070 ( 
.A1(n_4925),
.A2(n_155),
.B(n_156),
.Y(n_5070)
);

INVx1_ASAP7_75t_SL g5071 ( 
.A(n_4772),
.Y(n_5071)
);

AOI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4863),
.A2(n_157),
.B(n_158),
.Y(n_5072)
);

BUFx6f_ASAP7_75t_L g5073 ( 
.A(n_4779),
.Y(n_5073)
);

AND2x2_ASAP7_75t_L g5074 ( 
.A(n_4714),
.B(n_159),
.Y(n_5074)
);

OR2x2_ASAP7_75t_L g5075 ( 
.A(n_4841),
.B(n_159),
.Y(n_5075)
);

O2A1O1Ixp33_ASAP7_75t_L g5076 ( 
.A1(n_4891),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_5076)
);

NOR2xp33_ASAP7_75t_L g5077 ( 
.A(n_4800),
.B(n_160),
.Y(n_5077)
);

NOR2xp33_ASAP7_75t_L g5078 ( 
.A(n_4694),
.B(n_161),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4907),
.B(n_162),
.Y(n_5079)
);

INVx2_ASAP7_75t_L g5080 ( 
.A(n_4881),
.Y(n_5080)
);

NAND2xp5_ASAP7_75t_SL g5081 ( 
.A(n_4885),
.B(n_163),
.Y(n_5081)
);

AND2x4_ASAP7_75t_L g5082 ( 
.A(n_4791),
.B(n_164),
.Y(n_5082)
);

NOR2xp33_ASAP7_75t_L g5083 ( 
.A(n_4733),
.B(n_164),
.Y(n_5083)
);

AOI21xp5_ASAP7_75t_L g5084 ( 
.A1(n_4734),
.A2(n_165),
.B(n_166),
.Y(n_5084)
);

NAND3xp33_ASAP7_75t_L g5085 ( 
.A(n_4844),
.B(n_4691),
.C(n_4855),
.Y(n_5085)
);

AOI21xp5_ASAP7_75t_L g5086 ( 
.A1(n_4904),
.A2(n_165),
.B(n_167),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_4767),
.B(n_4843),
.Y(n_5087)
);

NOR2xp33_ASAP7_75t_L g5088 ( 
.A(n_4902),
.B(n_167),
.Y(n_5088)
);

OAI22x1_ASAP7_75t_L g5089 ( 
.A1(n_4819),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_5089)
);

OAI22xp5_ASAP7_75t_L g5090 ( 
.A1(n_4689),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_5090)
);

NOR2xp33_ASAP7_75t_SL g5091 ( 
.A(n_4692),
.B(n_4744),
.Y(n_5091)
);

O2A1O1Ixp5_ASAP7_75t_L g5092 ( 
.A1(n_4875),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_4896),
.B(n_171),
.Y(n_5093)
);

A2O1A1Ixp33_ASAP7_75t_L g5094 ( 
.A1(n_4684),
.A2(n_174),
.B(n_172),
.C(n_173),
.Y(n_5094)
);

INVx3_ASAP7_75t_L g5095 ( 
.A(n_4779),
.Y(n_5095)
);

AOI22xp5_ASAP7_75t_L g5096 ( 
.A1(n_4860),
.A2(n_177),
.B1(n_175),
.B2(n_176),
.Y(n_5096)
);

NOR2xp67_ASAP7_75t_L g5097 ( 
.A(n_4893),
.B(n_175),
.Y(n_5097)
);

AOI21xp5_ASAP7_75t_L g5098 ( 
.A1(n_4901),
.A2(n_176),
.B(n_179),
.Y(n_5098)
);

BUFx12f_ASAP7_75t_L g5099 ( 
.A(n_4692),
.Y(n_5099)
);

NOR2xp67_ASAP7_75t_L g5100 ( 
.A(n_4765),
.B(n_179),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4905),
.Y(n_5101)
);

OAI22xp5_ASAP7_75t_L g5102 ( 
.A1(n_4746),
.A2(n_183),
.B1(n_180),
.B2(n_181),
.Y(n_5102)
);

OAI22xp5_ASAP7_75t_L g5103 ( 
.A1(n_4795),
.A2(n_183),
.B1(n_180),
.B2(n_181),
.Y(n_5103)
);

A2O1A1Ixp33_ASAP7_75t_L g5104 ( 
.A1(n_4687),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_5104)
);

NAND2xp5_ASAP7_75t_L g5105 ( 
.A(n_4679),
.B(n_4894),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_4894),
.B(n_186),
.Y(n_5106)
);

NAND2xp5_ASAP7_75t_SL g5107 ( 
.A(n_4728),
.B(n_187),
.Y(n_5107)
);

AOI21xp5_ASAP7_75t_L g5108 ( 
.A1(n_4776),
.A2(n_189),
.B(n_190),
.Y(n_5108)
);

HB1xp67_ASAP7_75t_L g5109 ( 
.A(n_4898),
.Y(n_5109)
);

OR2x2_ASAP7_75t_L g5110 ( 
.A(n_4727),
.B(n_189),
.Y(n_5110)
);

OAI22x1_ASAP7_75t_L g5111 ( 
.A1(n_4877),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_5111)
);

OAI21x1_ASAP7_75t_L g5112 ( 
.A1(n_4708),
.A2(n_191),
.B(n_193),
.Y(n_5112)
);

BUFx3_ASAP7_75t_L g5113 ( 
.A(n_4695),
.Y(n_5113)
);

INVx3_ASAP7_75t_L g5114 ( 
.A(n_4869),
.Y(n_5114)
);

OR2x6_ASAP7_75t_SL g5115 ( 
.A(n_4707),
.B(n_194),
.Y(n_5115)
);

OAI22xp5_ASAP7_75t_L g5116 ( 
.A1(n_4702),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_5116)
);

INVx1_ASAP7_75t_L g5117 ( 
.A(n_4898),
.Y(n_5117)
);

NAND2xp5_ASAP7_75t_L g5118 ( 
.A(n_4849),
.B(n_196),
.Y(n_5118)
);

AND2x2_ASAP7_75t_L g5119 ( 
.A(n_4830),
.B(n_197),
.Y(n_5119)
);

AOI21xp5_ASAP7_75t_L g5120 ( 
.A1(n_4697),
.A2(n_199),
.B(n_200),
.Y(n_5120)
);

OAI21xp33_ASAP7_75t_L g5121 ( 
.A1(n_4798),
.A2(n_199),
.B(n_201),
.Y(n_5121)
);

HB1xp67_ASAP7_75t_L g5122 ( 
.A(n_4797),
.Y(n_5122)
);

NOR3xp33_ASAP7_75t_L g5123 ( 
.A(n_4897),
.B(n_202),
.C(n_203),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_4825),
.B(n_203),
.Y(n_5124)
);

OR2x6_ASAP7_75t_SL g5125 ( 
.A(n_4712),
.B(n_4782),
.Y(n_5125)
);

INVx2_ASAP7_75t_L g5126 ( 
.A(n_4887),
.Y(n_5126)
);

A2O1A1Ixp33_ASAP7_75t_L g5127 ( 
.A1(n_4775),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_5127)
);

BUFx6f_ASAP7_75t_L g5128 ( 
.A(n_4845),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_4737),
.A2(n_204),
.B(n_205),
.Y(n_5129)
);

OR2x6_ASAP7_75t_L g5130 ( 
.A(n_4823),
.B(n_206),
.Y(n_5130)
);

OAI21x1_ASAP7_75t_L g5131 ( 
.A1(n_4688),
.A2(n_207),
.B(n_210),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4755),
.B(n_207),
.Y(n_5132)
);

AOI21xp5_ASAP7_75t_L g5133 ( 
.A1(n_4773),
.A2(n_210),
.B(n_211),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_4731),
.Y(n_5134)
);

AOI21xp5_ASAP7_75t_L g5135 ( 
.A1(n_4829),
.A2(n_211),
.B(n_212),
.Y(n_5135)
);

OAI22xp5_ASAP7_75t_L g5136 ( 
.A1(n_4743),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_5136)
);

AOI21xp5_ASAP7_75t_L g5137 ( 
.A1(n_4857),
.A2(n_213),
.B(n_215),
.Y(n_5137)
);

INVx1_ASAP7_75t_L g5138 ( 
.A(n_4731),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_4811),
.Y(n_5139)
);

NOR2xp33_ASAP7_75t_L g5140 ( 
.A(n_4868),
.B(n_216),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_4758),
.A2(n_217),
.B(n_218),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_SL g5142 ( 
.A(n_4837),
.B(n_217),
.Y(n_5142)
);

NAND2xp33_ASAP7_75t_L g5143 ( 
.A(n_4777),
.B(n_218),
.Y(n_5143)
);

NAND2xp5_ASAP7_75t_SL g5144 ( 
.A(n_4762),
.B(n_219),
.Y(n_5144)
);

AOI21xp5_ASAP7_75t_L g5145 ( 
.A1(n_4763),
.A2(n_219),
.B(n_220),
.Y(n_5145)
);

AOI21xp5_ASAP7_75t_L g5146 ( 
.A1(n_4770),
.A2(n_220),
.B(n_221),
.Y(n_5146)
);

AOI33xp33_ASAP7_75t_L g5147 ( 
.A1(n_4842),
.A2(n_223),
.A3(n_227),
.B1(n_221),
.B2(n_222),
.B3(n_224),
.Y(n_5147)
);

AOI21xp5_ASAP7_75t_L g5148 ( 
.A1(n_4738),
.A2(n_223),
.B(n_229),
.Y(n_5148)
);

AOI21xp5_ASAP7_75t_L g5149 ( 
.A1(n_4793),
.A2(n_4846),
.B(n_4840),
.Y(n_5149)
);

INVx1_ASAP7_75t_L g5150 ( 
.A(n_4813),
.Y(n_5150)
);

INVx1_ASAP7_75t_L g5151 ( 
.A(n_4814),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4850),
.A2(n_230),
.B(n_231),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_4818),
.Y(n_5153)
);

INVx4_ASAP7_75t_L g5154 ( 
.A(n_4730),
.Y(n_5154)
);

INVx1_ASAP7_75t_L g5155 ( 
.A(n_4828),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_SL g5156 ( 
.A(n_4853),
.B(n_230),
.Y(n_5156)
);

BUFx6f_ASAP7_75t_L g5157 ( 
.A(n_4736),
.Y(n_5157)
);

AND2x4_ASAP7_75t_L g5158 ( 
.A(n_4804),
.B(n_4741),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4742),
.B(n_231),
.Y(n_5159)
);

O2A1O1Ixp33_ASAP7_75t_SL g5160 ( 
.A1(n_4748),
.A2(n_4750),
.B(n_4769),
.C(n_4761),
.Y(n_5160)
);

AOI21xp5_ASAP7_75t_L g5161 ( 
.A1(n_4771),
.A2(n_232),
.B(n_233),
.Y(n_5161)
);

INVx4_ASAP7_75t_L g5162 ( 
.A(n_4827),
.Y(n_5162)
);

AOI22xp5_ASAP7_75t_L g5163 ( 
.A1(n_4766),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_5163)
);

AOI22x1_ASAP7_75t_L g5164 ( 
.A1(n_4726),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_5164)
);

OR2x6_ASAP7_75t_L g5165 ( 
.A(n_4852),
.B(n_4839),
.Y(n_5165)
);

AND2x2_ASAP7_75t_SL g5166 ( 
.A(n_4711),
.B(n_235),
.Y(n_5166)
);

A2O1A1Ixp33_ASAP7_75t_L g5167 ( 
.A1(n_4722),
.A2(n_238),
.B(n_236),
.C(n_237),
.Y(n_5167)
);

AOI21xp5_ASAP7_75t_L g5168 ( 
.A1(n_4780),
.A2(n_239),
.B(n_240),
.Y(n_5168)
);

AO31x2_ASAP7_75t_L g5169 ( 
.A1(n_5134),
.A2(n_244),
.A3(n_240),
.B(n_242),
.Y(n_5169)
);

OAI22xp5_ASAP7_75t_L g5170 ( 
.A1(n_4963),
.A2(n_4940),
.B1(n_4985),
.B2(n_5014),
.Y(n_5170)
);

AOI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_4992),
.A2(n_242),
.B(n_244),
.Y(n_5171)
);

AOI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_4935),
.A2(n_245),
.B(n_246),
.Y(n_5172)
);

BUFx4_ASAP7_75t_SL g5173 ( 
.A(n_5055),
.Y(n_5173)
);

INVx1_ASAP7_75t_L g5174 ( 
.A(n_5002),
.Y(n_5174)
);

OAI21x1_ASAP7_75t_L g5175 ( 
.A1(n_4964),
.A2(n_246),
.B(n_247),
.Y(n_5175)
);

CKINVDCx5p33_ASAP7_75t_R g5176 ( 
.A(n_4950),
.Y(n_5176)
);

OAI21x1_ASAP7_75t_SL g5177 ( 
.A1(n_5049),
.A2(n_248),
.B(n_249),
.Y(n_5177)
);

OAI21x1_ASAP7_75t_L g5178 ( 
.A1(n_5025),
.A2(n_5027),
.B(n_5054),
.Y(n_5178)
);

AO31x2_ASAP7_75t_L g5179 ( 
.A1(n_5138),
.A2(n_252),
.A3(n_250),
.B(n_251),
.Y(n_5179)
);

OAI21x1_ASAP7_75t_L g5180 ( 
.A1(n_5004),
.A2(n_250),
.B(n_251),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_4979),
.B(n_252),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_4970),
.B(n_253),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_4937),
.A2(n_253),
.B(n_254),
.Y(n_5183)
);

OAI21x1_ASAP7_75t_SL g5184 ( 
.A1(n_5033),
.A2(n_254),
.B(n_255),
.Y(n_5184)
);

OAI21x1_ASAP7_75t_L g5185 ( 
.A1(n_4934),
.A2(n_255),
.B(n_256),
.Y(n_5185)
);

AOI21xp5_ASAP7_75t_L g5186 ( 
.A1(n_4956),
.A2(n_257),
.B(n_258),
.Y(n_5186)
);

AND2x2_ASAP7_75t_SL g5187 ( 
.A(n_5052),
.B(n_5091),
.Y(n_5187)
);

NAND2xp5_ASAP7_75t_L g5188 ( 
.A(n_4947),
.B(n_257),
.Y(n_5188)
);

OAI21xp33_ASAP7_75t_L g5189 ( 
.A1(n_5096),
.A2(n_259),
.B(n_260),
.Y(n_5189)
);

AND2x2_ASAP7_75t_L g5190 ( 
.A(n_5015),
.B(n_259),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_5011),
.Y(n_5191)
);

INVx1_ASAP7_75t_L g5192 ( 
.A(n_4996),
.Y(n_5192)
);

BUFx2_ASAP7_75t_L g5193 ( 
.A(n_5030),
.Y(n_5193)
);

HB1xp67_ASAP7_75t_L g5194 ( 
.A(n_5022),
.Y(n_5194)
);

AO21x1_ASAP7_75t_L g5195 ( 
.A1(n_4949),
.A2(n_260),
.B(n_261),
.Y(n_5195)
);

INVx2_ASAP7_75t_L g5196 ( 
.A(n_4958),
.Y(n_5196)
);

NOR4xp25_ASAP7_75t_L g5197 ( 
.A(n_4988),
.B(n_263),
.C(n_261),
.D(n_262),
.Y(n_5197)
);

AND2x2_ASAP7_75t_L g5198 ( 
.A(n_5087),
.B(n_262),
.Y(n_5198)
);

OAI21x1_ASAP7_75t_L g5199 ( 
.A1(n_5043),
.A2(n_263),
.B(n_264),
.Y(n_5199)
);

OAI21x1_ASAP7_75t_L g5200 ( 
.A1(n_5112),
.A2(n_264),
.B(n_265),
.Y(n_5200)
);

A2O1A1Ixp33_ASAP7_75t_L g5201 ( 
.A1(n_4974),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_5201)
);

OAI22x1_ASAP7_75t_L g5202 ( 
.A1(n_5059),
.A2(n_269),
.B1(n_266),
.B2(n_268),
.Y(n_5202)
);

OAI21x1_ASAP7_75t_L g5203 ( 
.A1(n_4938),
.A2(n_268),
.B(n_269),
.Y(n_5203)
);

AOI21xp5_ASAP7_75t_L g5204 ( 
.A1(n_4932),
.A2(n_270),
.B(n_271),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_SL g5205 ( 
.A1(n_4987),
.A2(n_270),
.B(n_271),
.Y(n_5205)
);

AND2x2_ASAP7_75t_L g5206 ( 
.A(n_4983),
.B(n_272),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_4968),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_5150),
.B(n_272),
.Y(n_5208)
);

AOI221x1_ASAP7_75t_L g5209 ( 
.A1(n_5089),
.A2(n_275),
.B1(n_273),
.B2(n_274),
.C(n_276),
.Y(n_5209)
);

OAI21x1_ASAP7_75t_L g5210 ( 
.A1(n_4980),
.A2(n_273),
.B(n_274),
.Y(n_5210)
);

OAI21x1_ASAP7_75t_L g5211 ( 
.A1(n_4993),
.A2(n_275),
.B(n_277),
.Y(n_5211)
);

NAND2xp5_ASAP7_75t_L g5212 ( 
.A(n_5151),
.B(n_277),
.Y(n_5212)
);

OAI21x1_ASAP7_75t_L g5213 ( 
.A1(n_4994),
.A2(n_4954),
.B(n_4944),
.Y(n_5213)
);

OA21x2_ASAP7_75t_L g5214 ( 
.A1(n_5070),
.A2(n_5084),
.B(n_5148),
.Y(n_5214)
);

OAI21x1_ASAP7_75t_SL g5215 ( 
.A1(n_5057),
.A2(n_278),
.B(n_279),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_5016),
.Y(n_5216)
);

AOI21xp5_ASAP7_75t_L g5217 ( 
.A1(n_5029),
.A2(n_278),
.B(n_279),
.Y(n_5217)
);

INVxp67_ASAP7_75t_SL g5218 ( 
.A(n_5105),
.Y(n_5218)
);

AOI21xp5_ASAP7_75t_L g5219 ( 
.A1(n_5029),
.A2(n_280),
.B(n_281),
.Y(n_5219)
);

BUFx2_ASAP7_75t_L g5220 ( 
.A(n_5060),
.Y(n_5220)
);

INVx3_ASAP7_75t_L g5221 ( 
.A(n_4969),
.Y(n_5221)
);

AOI21xp5_ASAP7_75t_L g5222 ( 
.A1(n_5029),
.A2(n_280),
.B(n_282),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4972),
.A2(n_282),
.B(n_283),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_5153),
.B(n_283),
.Y(n_5224)
);

BUFx2_ASAP7_75t_L g5225 ( 
.A(n_5038),
.Y(n_5225)
);

NAND2xp5_ASAP7_75t_L g5226 ( 
.A(n_5155),
.B(n_284),
.Y(n_5226)
);

AOI21x1_ASAP7_75t_L g5227 ( 
.A1(n_5012),
.A2(n_285),
.B(n_286),
.Y(n_5227)
);

OAI21x1_ASAP7_75t_L g5228 ( 
.A1(n_5126),
.A2(n_285),
.B(n_286),
.Y(n_5228)
);

AO31x2_ASAP7_75t_L g5229 ( 
.A1(n_5044),
.A2(n_5047),
.A3(n_4986),
.B(n_5080),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_5035),
.Y(n_5230)
);

OR2x6_ASAP7_75t_L g5231 ( 
.A(n_5099),
.B(n_287),
.Y(n_5231)
);

AND2x2_ASAP7_75t_L g5232 ( 
.A(n_5074),
.B(n_287),
.Y(n_5232)
);

AOI21xp5_ASAP7_75t_L g5233 ( 
.A1(n_4931),
.A2(n_5046),
.B(n_5037),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_5101),
.Y(n_5234)
);

AO31x2_ASAP7_75t_L g5235 ( 
.A1(n_5154),
.A2(n_290),
.A3(n_288),
.B(n_289),
.Y(n_5235)
);

BUFx2_ASAP7_75t_L g5236 ( 
.A(n_4997),
.Y(n_5236)
);

OAI21x1_ASAP7_75t_L g5237 ( 
.A1(n_5131),
.A2(n_288),
.B(n_289),
.Y(n_5237)
);

NOR2x1_ASAP7_75t_L g5238 ( 
.A(n_5023),
.B(n_291),
.Y(n_5238)
);

NAND2xp5_ASAP7_75t_L g5239 ( 
.A(n_5001),
.B(n_292),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_L g5240 ( 
.A(n_5139),
.B(n_292),
.Y(n_5240)
);

OAI21xp33_ASAP7_75t_L g5241 ( 
.A1(n_4999),
.A2(n_293),
.B(n_294),
.Y(n_5241)
);

OAI22xp5_ASAP7_75t_L g5242 ( 
.A1(n_5036),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_5242)
);

OAI22xp5_ASAP7_75t_L g5243 ( 
.A1(n_5065),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_5243)
);

OAI21x1_ASAP7_75t_L g5244 ( 
.A1(n_5149),
.A2(n_297),
.B(n_298),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_SL g5245 ( 
.A(n_5157),
.B(n_299),
.Y(n_5245)
);

OAI21x1_ASAP7_75t_L g5246 ( 
.A1(n_5092),
.A2(n_299),
.B(n_300),
.Y(n_5246)
);

OAI21x1_ASAP7_75t_L g5247 ( 
.A1(n_4955),
.A2(n_5039),
.B(n_5072),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_5117),
.Y(n_5248)
);

AO32x2_ASAP7_75t_L g5249 ( 
.A1(n_4953),
.A2(n_303),
.A3(n_300),
.B1(n_302),
.B2(n_305),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_4989),
.Y(n_5250)
);

AOI21xp5_ASAP7_75t_L g5251 ( 
.A1(n_5061),
.A2(n_302),
.B(n_303),
.Y(n_5251)
);

NOR2xp33_ASAP7_75t_L g5252 ( 
.A(n_5034),
.B(n_305),
.Y(n_5252)
);

OAI21x1_ASAP7_75t_L g5253 ( 
.A1(n_4982),
.A2(n_307),
.B(n_308),
.Y(n_5253)
);

AND2x4_ASAP7_75t_L g5254 ( 
.A(n_4942),
.B(n_308),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_4939),
.B(n_309),
.Y(n_5255)
);

NOR2xp67_ASAP7_75t_L g5256 ( 
.A(n_5066),
.B(n_309),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_5032),
.A2(n_310),
.B(n_311),
.Y(n_5257)
);

NOR2x1_ASAP7_75t_L g5258 ( 
.A(n_4936),
.B(n_5009),
.Y(n_5258)
);

O2A1O1Ixp33_ASAP7_75t_SL g5259 ( 
.A1(n_4965),
.A2(n_313),
.B(n_310),
.C(n_312),
.Y(n_5259)
);

NAND2xp5_ASAP7_75t_L g5260 ( 
.A(n_5019),
.B(n_312),
.Y(n_5260)
);

OAI21x1_ASAP7_75t_L g5261 ( 
.A1(n_5164),
.A2(n_313),
.B(n_314),
.Y(n_5261)
);

INVx3_ASAP7_75t_L g5262 ( 
.A(n_4969),
.Y(n_5262)
);

AOI21xp5_ASAP7_75t_L g5263 ( 
.A1(n_5051),
.A2(n_314),
.B(n_315),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_4951),
.B(n_315),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_4945),
.B(n_316),
.Y(n_5265)
);

NAND2x1_ASAP7_75t_L g5266 ( 
.A(n_5162),
.B(n_316),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_4976),
.B(n_317),
.Y(n_5267)
);

AND2x2_ASAP7_75t_L g5268 ( 
.A(n_5119),
.B(n_317),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_SL g5269 ( 
.A(n_5157),
.B(n_318),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_L g5270 ( 
.A(n_4966),
.B(n_318),
.Y(n_5270)
);

AND2x4_ASAP7_75t_L g5271 ( 
.A(n_5000),
.B(n_319),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_5109),
.B(n_320),
.Y(n_5272)
);

OAI21xp5_ASAP7_75t_L g5273 ( 
.A1(n_4995),
.A2(n_320),
.B(n_322),
.Y(n_5273)
);

AOI21xp5_ASAP7_75t_L g5274 ( 
.A1(n_5160),
.A2(n_322),
.B(n_323),
.Y(n_5274)
);

NAND2xp5_ASAP7_75t_L g5275 ( 
.A(n_5024),
.B(n_324),
.Y(n_5275)
);

INVx1_ASAP7_75t_L g5276 ( 
.A(n_5028),
.Y(n_5276)
);

AND2x2_ASAP7_75t_SL g5277 ( 
.A(n_5166),
.B(n_325),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_4941),
.A2(n_326),
.B(n_327),
.Y(n_5278)
);

NAND3xp33_ASAP7_75t_L g5279 ( 
.A(n_5042),
.B(n_326),
.C(n_328),
.Y(n_5279)
);

NAND2xp5_ASAP7_75t_L g5280 ( 
.A(n_5040),
.B(n_5041),
.Y(n_5280)
);

OAI21x1_ASAP7_75t_L g5281 ( 
.A1(n_5086),
.A2(n_328),
.B(n_329),
.Y(n_5281)
);

OAI21x1_ASAP7_75t_L g5282 ( 
.A1(n_5098),
.A2(n_329),
.B(n_330),
.Y(n_5282)
);

AOI21xp5_ASAP7_75t_L g5283 ( 
.A1(n_5121),
.A2(n_5158),
.B(n_5076),
.Y(n_5283)
);

OAI21x1_ASAP7_75t_L g5284 ( 
.A1(n_5168),
.A2(n_331),
.B(n_332),
.Y(n_5284)
);

OAI21x1_ASAP7_75t_L g5285 ( 
.A1(n_5135),
.A2(n_331),
.B(n_332),
.Y(n_5285)
);

OAI21x1_ASAP7_75t_L g5286 ( 
.A1(n_5161),
.A2(n_333),
.B(n_334),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_5124),
.B(n_334),
.Y(n_5287)
);

OR2x2_ASAP7_75t_L g5288 ( 
.A(n_5075),
.B(n_335),
.Y(n_5288)
);

AND2x2_ASAP7_75t_L g5289 ( 
.A(n_5005),
.B(n_335),
.Y(n_5289)
);

AND2x2_ASAP7_75t_L g5290 ( 
.A(n_4971),
.B(n_4933),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_L g5291 ( 
.A(n_5071),
.B(n_336),
.Y(n_5291)
);

INVx1_ASAP7_75t_SL g5292 ( 
.A(n_5003),
.Y(n_5292)
);

AOI211x1_ASAP7_75t_L g5293 ( 
.A1(n_5010),
.A2(n_340),
.B(n_337),
.C(n_339),
.Y(n_5293)
);

OAI21xp5_ASAP7_75t_L g5294 ( 
.A1(n_4961),
.A2(n_337),
.B(n_339),
.Y(n_5294)
);

NAND2x1p5_ASAP7_75t_L g5295 ( 
.A(n_5073),
.B(n_341),
.Y(n_5295)
);

AO32x2_ASAP7_75t_L g5296 ( 
.A1(n_4973),
.A2(n_343),
.A3(n_341),
.B1(n_342),
.B2(n_344),
.Y(n_5296)
);

OAI21xp5_ASAP7_75t_L g5297 ( 
.A1(n_5064),
.A2(n_342),
.B(n_344),
.Y(n_5297)
);

AOI21xp5_ASAP7_75t_L g5298 ( 
.A1(n_5165),
.A2(n_345),
.B(n_346),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_L g5299 ( 
.A(n_5114),
.B(n_347),
.Y(n_5299)
);

AO21x1_ASAP7_75t_L g5300 ( 
.A1(n_4977),
.A2(n_347),
.B(n_348),
.Y(n_5300)
);

OAI21x1_ASAP7_75t_L g5301 ( 
.A1(n_5152),
.A2(n_350),
.B(n_351),
.Y(n_5301)
);

OAI22xp5_ASAP7_75t_L g5302 ( 
.A1(n_4959),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_5302)
);

OAI21x1_ASAP7_75t_L g5303 ( 
.A1(n_4960),
.A2(n_355),
.B(n_356),
.Y(n_5303)
);

INVx1_ASAP7_75t_SL g5304 ( 
.A(n_5113),
.Y(n_5304)
);

AOI21xp5_ASAP7_75t_L g5305 ( 
.A1(n_5165),
.A2(n_5068),
.B(n_5045),
.Y(n_5305)
);

CKINVDCx11_ASAP7_75t_R g5306 ( 
.A(n_4952),
.Y(n_5306)
);

NAND2xp5_ASAP7_75t_L g5307 ( 
.A(n_5122),
.B(n_356),
.Y(n_5307)
);

OAI21x1_ASAP7_75t_L g5308 ( 
.A1(n_4998),
.A2(n_357),
.B(n_358),
.Y(n_5308)
);

INVxp67_ASAP7_75t_SL g5309 ( 
.A(n_5093),
.Y(n_5309)
);

INVx2_ASAP7_75t_L g5310 ( 
.A(n_5106),
.Y(n_5310)
);

OAI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_5104),
.A2(n_357),
.B(n_359),
.Y(n_5311)
);

AOI21xp5_ASAP7_75t_L g5312 ( 
.A1(n_5008),
.A2(n_360),
.B(n_361),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_5079),
.Y(n_5313)
);

CKINVDCx5p33_ASAP7_75t_R g5314 ( 
.A(n_5073),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_4967),
.B(n_361),
.Y(n_5315)
);

AO31x2_ASAP7_75t_L g5316 ( 
.A1(n_5062),
.A2(n_364),
.A3(n_362),
.B(n_363),
.Y(n_5316)
);

INVx2_ASAP7_75t_SL g5317 ( 
.A(n_5095),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_L g5318 ( 
.A(n_5026),
.B(n_362),
.Y(n_5318)
);

AND2x2_ASAP7_75t_L g5319 ( 
.A(n_5118),
.B(n_363),
.Y(n_5319)
);

OAI21x1_ASAP7_75t_SL g5320 ( 
.A1(n_5007),
.A2(n_364),
.B(n_365),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_5097),
.B(n_365),
.Y(n_5321)
);

A2O1A1Ixp33_ASAP7_75t_L g5322 ( 
.A1(n_5085),
.A2(n_368),
.B(n_366),
.C(n_367),
.Y(n_5322)
);

AND2x2_ASAP7_75t_L g5323 ( 
.A(n_5082),
.B(n_366),
.Y(n_5323)
);

OAI21x1_ASAP7_75t_L g5324 ( 
.A1(n_5013),
.A2(n_367),
.B(n_368),
.Y(n_5324)
);

OAI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_5094),
.A2(n_369),
.B(n_370),
.Y(n_5325)
);

OAI21x1_ASAP7_75t_L g5326 ( 
.A1(n_5031),
.A2(n_5129),
.B(n_5108),
.Y(n_5326)
);

OAI21x1_ASAP7_75t_L g5327 ( 
.A1(n_5133),
.A2(n_369),
.B(n_373),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_5053),
.B(n_373),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_5017),
.B(n_374),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5021),
.Y(n_5330)
);

OAI21xp5_ASAP7_75t_L g5331 ( 
.A1(n_5127),
.A2(n_375),
.B(n_376),
.Y(n_5331)
);

AND2x2_ASAP7_75t_L g5332 ( 
.A(n_5083),
.B(n_376),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_L g5333 ( 
.A(n_5069),
.B(n_377),
.Y(n_5333)
);

NOR4xp25_ASAP7_75t_L g5334 ( 
.A(n_5090),
.B(n_379),
.C(n_377),
.D(n_378),
.Y(n_5334)
);

AO31x2_ASAP7_75t_L g5335 ( 
.A1(n_5103),
.A2(n_381),
.A3(n_378),
.B(n_380),
.Y(n_5335)
);

AOI21xp5_ASAP7_75t_L g5336 ( 
.A1(n_5123),
.A2(n_381),
.B(n_382),
.Y(n_5336)
);

BUFx6f_ASAP7_75t_L g5337 ( 
.A(n_5128),
.Y(n_5337)
);

BUFx2_ASAP7_75t_L g5338 ( 
.A(n_5058),
.Y(n_5338)
);

OA22x2_ASAP7_75t_L g5339 ( 
.A1(n_5130),
.A2(n_386),
.B1(n_383),
.B2(n_385),
.Y(n_5339)
);

AND2x2_ASAP7_75t_L g5340 ( 
.A(n_4943),
.B(n_383),
.Y(n_5340)
);

AOI21xp5_ASAP7_75t_L g5341 ( 
.A1(n_5156),
.A2(n_385),
.B(n_386),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_5048),
.B(n_5078),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_5110),
.B(n_387),
.Y(n_5343)
);

O2A1O1Ixp5_ASAP7_75t_L g5344 ( 
.A1(n_4948),
.A2(n_389),
.B(n_387),
.C(n_388),
.Y(n_5344)
);

OAI22xp5_ASAP7_75t_L g5345 ( 
.A1(n_5163),
.A2(n_390),
.B1(n_388),
.B2(n_389),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5194),
.Y(n_5346)
);

BUFx6f_ASAP7_75t_L g5347 ( 
.A(n_5337),
.Y(n_5347)
);

AND2x4_ASAP7_75t_L g5348 ( 
.A(n_5220),
.B(n_5128),
.Y(n_5348)
);

AOI21xp5_ASAP7_75t_L g5349 ( 
.A1(n_5233),
.A2(n_4946),
.B(n_4962),
.Y(n_5349)
);

BUFx2_ASAP7_75t_SL g5350 ( 
.A(n_5256),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5229),
.Y(n_5351)
);

AOI21xp5_ASAP7_75t_L g5352 ( 
.A1(n_5283),
.A2(n_4975),
.B(n_5144),
.Y(n_5352)
);

BUFx6f_ASAP7_75t_L g5353 ( 
.A(n_5337),
.Y(n_5353)
);

AND2x2_ASAP7_75t_L g5354 ( 
.A(n_5193),
.B(n_5125),
.Y(n_5354)
);

BUFx10_ASAP7_75t_L g5355 ( 
.A(n_5176),
.Y(n_5355)
);

INVx4_ASAP7_75t_L g5356 ( 
.A(n_5314),
.Y(n_5356)
);

OAI21xp33_ASAP7_75t_L g5357 ( 
.A1(n_5170),
.A2(n_5189),
.B(n_5201),
.Y(n_5357)
);

NAND2xp5_ASAP7_75t_L g5358 ( 
.A(n_5191),
.B(n_5115),
.Y(n_5358)
);

INVx2_ASAP7_75t_SL g5359 ( 
.A(n_5236),
.Y(n_5359)
);

AND2x2_ASAP7_75t_L g5360 ( 
.A(n_5290),
.B(n_5088),
.Y(n_5360)
);

OAI22xp5_ASAP7_75t_L g5361 ( 
.A1(n_5277),
.A2(n_5130),
.B1(n_4991),
.B2(n_5140),
.Y(n_5361)
);

INVx3_ASAP7_75t_L g5362 ( 
.A(n_5221),
.Y(n_5362)
);

AND2x2_ASAP7_75t_L g5363 ( 
.A(n_5174),
.B(n_5230),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_5305),
.A2(n_5274),
.B(n_5263),
.Y(n_5364)
);

INVx2_ASAP7_75t_SL g5365 ( 
.A(n_5317),
.Y(n_5365)
);

INVx2_ASAP7_75t_SL g5366 ( 
.A(n_5262),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_5309),
.B(n_5132),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5229),
.Y(n_5368)
);

INVx3_ASAP7_75t_L g5369 ( 
.A(n_5292),
.Y(n_5369)
);

INVx2_ASAP7_75t_SL g5370 ( 
.A(n_5304),
.Y(n_5370)
);

AND2x2_ASAP7_75t_L g5371 ( 
.A(n_5198),
.B(n_5056),
.Y(n_5371)
);

OAI21x1_ASAP7_75t_SL g5372 ( 
.A1(n_5195),
.A2(n_5145),
.B(n_5141),
.Y(n_5372)
);

INVx2_ASAP7_75t_SL g5373 ( 
.A(n_5173),
.Y(n_5373)
);

BUFx6f_ASAP7_75t_L g5374 ( 
.A(n_5338),
.Y(n_5374)
);

BUFx3_ASAP7_75t_L g5375 ( 
.A(n_5306),
.Y(n_5375)
);

AOI22xp33_ASAP7_75t_SL g5376 ( 
.A1(n_5187),
.A2(n_4978),
.B1(n_4957),
.B2(n_5077),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_5192),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_L g5378 ( 
.A(n_5250),
.B(n_5147),
.Y(n_5378)
);

INVx4_ASAP7_75t_L g5379 ( 
.A(n_5254),
.Y(n_5379)
);

BUFx3_ASAP7_75t_L g5380 ( 
.A(n_5225),
.Y(n_5380)
);

INVx2_ASAP7_75t_SL g5381 ( 
.A(n_5310),
.Y(n_5381)
);

INVxp67_ASAP7_75t_L g5382 ( 
.A(n_5313),
.Y(n_5382)
);

AOI22xp5_ASAP7_75t_L g5383 ( 
.A1(n_5241),
.A2(n_5142),
.B1(n_5143),
.B2(n_5067),
.Y(n_5383)
);

HB1xp67_ASAP7_75t_L g5384 ( 
.A(n_5330),
.Y(n_5384)
);

INVx2_ASAP7_75t_SL g5385 ( 
.A(n_5248),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_5276),
.B(n_5050),
.Y(n_5386)
);

AND2x4_ASAP7_75t_L g5387 ( 
.A(n_5218),
.B(n_5100),
.Y(n_5387)
);

BUFx12f_ASAP7_75t_L g5388 ( 
.A(n_5231),
.Y(n_5388)
);

AOI21xp5_ASAP7_75t_L g5389 ( 
.A1(n_5171),
.A2(n_5146),
.B(n_5107),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_SL g5390 ( 
.A(n_5258),
.B(n_5081),
.Y(n_5390)
);

INVx1_ASAP7_75t_L g5391 ( 
.A(n_5234),
.Y(n_5391)
);

INVx2_ASAP7_75t_L g5392 ( 
.A(n_5196),
.Y(n_5392)
);

INVx2_ASAP7_75t_SL g5393 ( 
.A(n_5272),
.Y(n_5393)
);

CKINVDCx20_ASAP7_75t_R g5394 ( 
.A(n_5323),
.Y(n_5394)
);

INVxp67_ASAP7_75t_SL g5395 ( 
.A(n_5280),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_5207),
.Y(n_5396)
);

AOI22xp33_ASAP7_75t_L g5397 ( 
.A1(n_5294),
.A2(n_5102),
.B1(n_5136),
.B2(n_5116),
.Y(n_5397)
);

BUFx2_ASAP7_75t_L g5398 ( 
.A(n_5181),
.Y(n_5398)
);

INVx2_ASAP7_75t_SL g5399 ( 
.A(n_5271),
.Y(n_5399)
);

INVx4_ASAP7_75t_L g5400 ( 
.A(n_5231),
.Y(n_5400)
);

BUFx3_ASAP7_75t_L g5401 ( 
.A(n_5190),
.Y(n_5401)
);

INVx1_ASAP7_75t_L g5402 ( 
.A(n_5216),
.Y(n_5402)
);

A2O1A1Ixp33_ASAP7_75t_L g5403 ( 
.A1(n_5186),
.A2(n_5137),
.B(n_5120),
.C(n_5167),
.Y(n_5403)
);

OAI22xp5_ASAP7_75t_L g5404 ( 
.A1(n_5279),
.A2(n_5063),
.B1(n_4981),
.B2(n_5159),
.Y(n_5404)
);

INVx3_ASAP7_75t_L g5405 ( 
.A(n_5289),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5182),
.Y(n_5406)
);

OR2x2_ASAP7_75t_L g5407 ( 
.A(n_5188),
.B(n_5018),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_5169),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5169),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5179),
.Y(n_5410)
);

AND2x2_ASAP7_75t_L g5411 ( 
.A(n_5268),
.B(n_5206),
.Y(n_5411)
);

BUFx8_ASAP7_75t_SL g5412 ( 
.A(n_5342),
.Y(n_5412)
);

NOR2xp67_ASAP7_75t_L g5413 ( 
.A(n_5208),
.B(n_5111),
.Y(n_5413)
);

BUFx6f_ASAP7_75t_L g5414 ( 
.A(n_5295),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5179),
.Y(n_5415)
);

BUFx5_ASAP7_75t_L g5416 ( 
.A(n_5332),
.Y(n_5416)
);

AND2x4_ASAP7_75t_L g5417 ( 
.A(n_5232),
.B(n_5006),
.Y(n_5417)
);

CKINVDCx5p33_ASAP7_75t_R g5418 ( 
.A(n_5287),
.Y(n_5418)
);

AND2x2_ASAP7_75t_L g5419 ( 
.A(n_5340),
.B(n_5319),
.Y(n_5419)
);

INVx1_ASAP7_75t_L g5420 ( 
.A(n_5235),
.Y(n_5420)
);

INVx2_ASAP7_75t_L g5421 ( 
.A(n_5235),
.Y(n_5421)
);

OR2x2_ASAP7_75t_L g5422 ( 
.A(n_5288),
.B(n_5020),
.Y(n_5422)
);

NOR2xp33_ASAP7_75t_L g5423 ( 
.A(n_5328),
.B(n_391),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_5240),
.Y(n_5424)
);

BUFx6f_ASAP7_75t_L g5425 ( 
.A(n_5299),
.Y(n_5425)
);

OAI22xp5_ASAP7_75t_L g5426 ( 
.A1(n_5311),
.A2(n_4990),
.B1(n_4984),
.B2(n_393),
.Y(n_5426)
);

BUFx6f_ASAP7_75t_L g5427 ( 
.A(n_5291),
.Y(n_5427)
);

NAND2xp5_ASAP7_75t_L g5428 ( 
.A(n_5212),
.B(n_391),
.Y(n_5428)
);

CKINVDCx11_ASAP7_75t_R g5429 ( 
.A(n_5243),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_5224),
.B(n_392),
.Y(n_5430)
);

OR2x2_ASAP7_75t_L g5431 ( 
.A(n_5226),
.B(n_392),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_5228),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_5227),
.Y(n_5433)
);

INVx1_ASAP7_75t_SL g5434 ( 
.A(n_5307),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_5296),
.Y(n_5435)
);

AOI222xp33_ASAP7_75t_L g5436 ( 
.A1(n_5333),
.A2(n_395),
.B1(n_397),
.B2(n_393),
.C1(n_394),
.C2(n_396),
.Y(n_5436)
);

AND2x2_ASAP7_75t_L g5437 ( 
.A(n_5343),
.B(n_394),
.Y(n_5437)
);

AOI22xp5_ASAP7_75t_L g5438 ( 
.A1(n_5252),
.A2(n_398),
.B1(n_395),
.B2(n_397),
.Y(n_5438)
);

NAND2x1p5_ASAP7_75t_L g5439 ( 
.A(n_5266),
.B(n_398),
.Y(n_5439)
);

AOI21xp5_ASAP7_75t_SL g5440 ( 
.A1(n_5273),
.A2(n_399),
.B(n_400),
.Y(n_5440)
);

AOI22xp5_ASAP7_75t_SL g5441 ( 
.A1(n_5339),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_5441)
);

AOI21xp5_ASAP7_75t_L g5442 ( 
.A1(n_5204),
.A2(n_401),
.B(n_402),
.Y(n_5442)
);

AOI21xp5_ASAP7_75t_L g5443 ( 
.A1(n_5213),
.A2(n_5331),
.B(n_5325),
.Y(n_5443)
);

INVx2_ASAP7_75t_SL g5444 ( 
.A(n_5239),
.Y(n_5444)
);

NAND2xp5_ASAP7_75t_L g5445 ( 
.A(n_5260),
.B(n_402),
.Y(n_5445)
);

O2A1O1Ixp33_ASAP7_75t_L g5446 ( 
.A1(n_5322),
.A2(n_405),
.B(n_403),
.C(n_404),
.Y(n_5446)
);

AND2x4_ASAP7_75t_L g5447 ( 
.A(n_5238),
.B(n_403),
.Y(n_5447)
);

INVx3_ASAP7_75t_L g5448 ( 
.A(n_5326),
.Y(n_5448)
);

OAI21x1_ASAP7_75t_L g5449 ( 
.A1(n_5178),
.A2(n_406),
.B(n_407),
.Y(n_5449)
);

OAI22xp5_ASAP7_75t_L g5450 ( 
.A1(n_5318),
.A2(n_411),
.B1(n_407),
.B2(n_408),
.Y(n_5450)
);

AND2x4_ASAP7_75t_L g5451 ( 
.A(n_5245),
.B(n_408),
.Y(n_5451)
);

AOI21xp5_ASAP7_75t_L g5452 ( 
.A1(n_5205),
.A2(n_411),
.B(n_412),
.Y(n_5452)
);

NAND2x1p5_ASAP7_75t_L g5453 ( 
.A(n_5269),
.B(n_412),
.Y(n_5453)
);

AND2x4_ASAP7_75t_L g5454 ( 
.A(n_5298),
.B(n_413),
.Y(n_5454)
);

CKINVDCx6p67_ASAP7_75t_R g5455 ( 
.A(n_5202),
.Y(n_5455)
);

BUFx10_ASAP7_75t_L g5456 ( 
.A(n_5264),
.Y(n_5456)
);

A2O1A1Ixp33_ASAP7_75t_L g5457 ( 
.A1(n_5251),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_5457)
);

AND2x4_ASAP7_75t_L g5458 ( 
.A(n_5217),
.B(n_416),
.Y(n_5458)
);

INVx3_ASAP7_75t_L g5459 ( 
.A(n_5199),
.Y(n_5459)
);

INVx3_ASAP7_75t_L g5460 ( 
.A(n_5247),
.Y(n_5460)
);

NAND2xp5_ASAP7_75t_L g5461 ( 
.A(n_5255),
.B(n_417),
.Y(n_5461)
);

AOI21xp5_ASAP7_75t_L g5462 ( 
.A1(n_5259),
.A2(n_418),
.B(n_419),
.Y(n_5462)
);

INVx1_ASAP7_75t_L g5463 ( 
.A(n_5296),
.Y(n_5463)
);

INVxp67_ASAP7_75t_L g5464 ( 
.A(n_5265),
.Y(n_5464)
);

INVx3_ASAP7_75t_L g5465 ( 
.A(n_5244),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5249),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5249),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_L g5468 ( 
.A(n_5270),
.B(n_5267),
.Y(n_5468)
);

NAND2x1p5_ASAP7_75t_L g5469 ( 
.A(n_5185),
.B(n_418),
.Y(n_5469)
);

INVx3_ASAP7_75t_L g5470 ( 
.A(n_5374),
.Y(n_5470)
);

INVx1_ASAP7_75t_L g5471 ( 
.A(n_5384),
.Y(n_5471)
);

INVx2_ASAP7_75t_L g5472 ( 
.A(n_5385),
.Y(n_5472)
);

BUFx2_ASAP7_75t_L g5473 ( 
.A(n_5416),
.Y(n_5473)
);

INVx1_ASAP7_75t_SL g5474 ( 
.A(n_5412),
.Y(n_5474)
);

AOI22xp33_ASAP7_75t_SL g5475 ( 
.A1(n_5435),
.A2(n_5177),
.B1(n_5184),
.B2(n_5297),
.Y(n_5475)
);

BUFx3_ASAP7_75t_L g5476 ( 
.A(n_5373),
.Y(n_5476)
);

INVx1_ASAP7_75t_L g5477 ( 
.A(n_5377),
.Y(n_5477)
);

INVx1_ASAP7_75t_L g5478 ( 
.A(n_5346),
.Y(n_5478)
);

OAI22xp33_ASAP7_75t_L g5479 ( 
.A1(n_5455),
.A2(n_5209),
.B1(n_5242),
.B2(n_5278),
.Y(n_5479)
);

CKINVDCx11_ASAP7_75t_R g5480 ( 
.A(n_5355),
.Y(n_5480)
);

OAI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_5349),
.A2(n_5345),
.B1(n_5222),
.B2(n_5219),
.Y(n_5481)
);

AOI22xp33_ASAP7_75t_L g5482 ( 
.A1(n_5357),
.A2(n_5300),
.B1(n_5215),
.B2(n_5336),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_5391),
.Y(n_5483)
);

AOI22xp33_ASAP7_75t_L g5484 ( 
.A1(n_5463),
.A2(n_5467),
.B1(n_5466),
.B2(n_5429),
.Y(n_5484)
);

CKINVDCx11_ASAP7_75t_R g5485 ( 
.A(n_5394),
.Y(n_5485)
);

BUFx6f_ASAP7_75t_L g5486 ( 
.A(n_5347),
.Y(n_5486)
);

INVx6_ASAP7_75t_L g5487 ( 
.A(n_5356),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_5392),
.Y(n_5488)
);

BUFx12f_ASAP7_75t_L g5489 ( 
.A(n_5388),
.Y(n_5489)
);

OAI21xp33_ASAP7_75t_L g5490 ( 
.A1(n_5440),
.A2(n_5334),
.B(n_5197),
.Y(n_5490)
);

AOI22xp33_ASAP7_75t_L g5491 ( 
.A1(n_5436),
.A2(n_5312),
.B1(n_5183),
.B2(n_5214),
.Y(n_5491)
);

BUFx12f_ASAP7_75t_L g5492 ( 
.A(n_5400),
.Y(n_5492)
);

BUFx2_ASAP7_75t_SL g5493 ( 
.A(n_5375),
.Y(n_5493)
);

CKINVDCx11_ASAP7_75t_R g5494 ( 
.A(n_5456),
.Y(n_5494)
);

INVx3_ASAP7_75t_L g5495 ( 
.A(n_5374),
.Y(n_5495)
);

OAI22xp5_ASAP7_75t_L g5496 ( 
.A1(n_5397),
.A2(n_5293),
.B1(n_5302),
.B2(n_5329),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5363),
.Y(n_5497)
);

BUFx3_ASAP7_75t_L g5498 ( 
.A(n_5369),
.Y(n_5498)
);

BUFx12f_ASAP7_75t_L g5499 ( 
.A(n_5414),
.Y(n_5499)
);

INVx1_ASAP7_75t_L g5500 ( 
.A(n_5382),
.Y(n_5500)
);

BUFx2_ASAP7_75t_R g5501 ( 
.A(n_5380),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5395),
.Y(n_5502)
);

INVx4_ASAP7_75t_L g5503 ( 
.A(n_5379),
.Y(n_5503)
);

OAI22xp33_ASAP7_75t_L g5504 ( 
.A1(n_5361),
.A2(n_5321),
.B1(n_5315),
.B2(n_5275),
.Y(n_5504)
);

HB1xp67_ASAP7_75t_SL g5505 ( 
.A(n_5350),
.Y(n_5505)
);

INVx4_ASAP7_75t_L g5506 ( 
.A(n_5348),
.Y(n_5506)
);

INVx1_ASAP7_75t_L g5507 ( 
.A(n_5408),
.Y(n_5507)
);

OAI21xp5_ASAP7_75t_L g5508 ( 
.A1(n_5443),
.A2(n_5364),
.B(n_5352),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5409),
.Y(n_5509)
);

BUFx3_ASAP7_75t_L g5510 ( 
.A(n_5370),
.Y(n_5510)
);

OAI22xp5_ASAP7_75t_L g5511 ( 
.A1(n_5383),
.A2(n_5172),
.B1(n_5341),
.B2(n_5316),
.Y(n_5511)
);

INVx3_ASAP7_75t_L g5512 ( 
.A(n_5347),
.Y(n_5512)
);

NAND2xp5_ASAP7_75t_L g5513 ( 
.A(n_5406),
.B(n_5335),
.Y(n_5513)
);

AOI22xp33_ASAP7_75t_L g5514 ( 
.A1(n_5452),
.A2(n_5320),
.B1(n_5327),
.B2(n_5284),
.Y(n_5514)
);

AOI22xp33_ASAP7_75t_L g5515 ( 
.A1(n_5413),
.A2(n_5301),
.B1(n_5285),
.B2(n_5303),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5410),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_5415),
.Y(n_5517)
);

INVx1_ASAP7_75t_L g5518 ( 
.A(n_5396),
.Y(n_5518)
);

AOI22xp33_ASAP7_75t_L g5519 ( 
.A1(n_5372),
.A2(n_5427),
.B1(n_5376),
.B2(n_5462),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5402),
.Y(n_5520)
);

OAI22xp5_ASAP7_75t_L g5521 ( 
.A1(n_5438),
.A2(n_5316),
.B1(n_5335),
.B2(n_5344),
.Y(n_5521)
);

INVx3_ASAP7_75t_L g5522 ( 
.A(n_5353),
.Y(n_5522)
);

AOI22xp33_ASAP7_75t_L g5523 ( 
.A1(n_5427),
.A2(n_5286),
.B1(n_5308),
.B2(n_5324),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5420),
.Y(n_5524)
);

AND2x2_ASAP7_75t_L g5525 ( 
.A(n_5354),
.B(n_5175),
.Y(n_5525)
);

INVx6_ASAP7_75t_L g5526 ( 
.A(n_5353),
.Y(n_5526)
);

NAND2xp5_ASAP7_75t_L g5527 ( 
.A(n_5398),
.B(n_5281),
.Y(n_5527)
);

AOI22xp33_ASAP7_75t_L g5528 ( 
.A1(n_5442),
.A2(n_5282),
.B1(n_5223),
.B2(n_5203),
.Y(n_5528)
);

INVx1_ASAP7_75t_L g5529 ( 
.A(n_5351),
.Y(n_5529)
);

OAI22xp5_ASAP7_75t_L g5530 ( 
.A1(n_5453),
.A2(n_5210),
.B1(n_5211),
.B2(n_5261),
.Y(n_5530)
);

AOI22xp33_ASAP7_75t_L g5531 ( 
.A1(n_5424),
.A2(n_5253),
.B1(n_5180),
.B2(n_5257),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_5368),
.Y(n_5532)
);

OAI22xp5_ASAP7_75t_L g5533 ( 
.A1(n_5454),
.A2(n_5237),
.B1(n_5200),
.B2(n_5246),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5421),
.Y(n_5534)
);

BUFx6f_ASAP7_75t_L g5535 ( 
.A(n_5414),
.Y(n_5535)
);

AOI22xp33_ASAP7_75t_L g5536 ( 
.A1(n_5387),
.A2(n_422),
.B1(n_420),
.B2(n_421),
.Y(n_5536)
);

INVx1_ASAP7_75t_L g5537 ( 
.A(n_5381),
.Y(n_5537)
);

BUFx10_ASAP7_75t_L g5538 ( 
.A(n_5423),
.Y(n_5538)
);

INVx2_ASAP7_75t_R g5539 ( 
.A(n_5433),
.Y(n_5539)
);

CKINVDCx11_ASAP7_75t_R g5540 ( 
.A(n_5416),
.Y(n_5540)
);

AOI22xp33_ASAP7_75t_SL g5541 ( 
.A1(n_5441),
.A2(n_424),
.B1(n_420),
.B2(n_423),
.Y(n_5541)
);

AOI22xp33_ASAP7_75t_L g5542 ( 
.A1(n_5389),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_5542)
);

INVx1_ASAP7_75t_L g5543 ( 
.A(n_5432),
.Y(n_5543)
);

AOI22xp33_ASAP7_75t_L g5544 ( 
.A1(n_5378),
.A2(n_428),
.B1(n_425),
.B2(n_426),
.Y(n_5544)
);

INVx3_ASAP7_75t_L g5545 ( 
.A(n_5362),
.Y(n_5545)
);

INVx6_ASAP7_75t_L g5546 ( 
.A(n_5401),
.Y(n_5546)
);

OAI22xp5_ASAP7_75t_L g5547 ( 
.A1(n_5457),
.A2(n_431),
.B1(n_429),
.B2(n_430),
.Y(n_5547)
);

BUFx3_ASAP7_75t_L g5548 ( 
.A(n_5359),
.Y(n_5548)
);

BUFx6f_ASAP7_75t_L g5549 ( 
.A(n_5366),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_5448),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_5367),
.B(n_429),
.Y(n_5551)
);

AOI22xp33_ASAP7_75t_SL g5552 ( 
.A1(n_5434),
.A2(n_432),
.B1(n_430),
.B2(n_431),
.Y(n_5552)
);

OAI22xp5_ASAP7_75t_L g5553 ( 
.A1(n_5426),
.A2(n_434),
.B1(n_432),
.B2(n_433),
.Y(n_5553)
);

INVx2_ASAP7_75t_L g5554 ( 
.A(n_5460),
.Y(n_5554)
);

BUFx3_ASAP7_75t_L g5555 ( 
.A(n_5365),
.Y(n_5555)
);

OAI21xp5_ASAP7_75t_SL g5556 ( 
.A1(n_5450),
.A2(n_434),
.B(n_435),
.Y(n_5556)
);

INVx4_ASAP7_75t_L g5557 ( 
.A(n_5425),
.Y(n_5557)
);

INVx2_ASAP7_75t_L g5558 ( 
.A(n_5459),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5386),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5358),
.Y(n_5560)
);

INVx3_ASAP7_75t_L g5561 ( 
.A(n_5425),
.Y(n_5561)
);

AOI22xp33_ASAP7_75t_L g5562 ( 
.A1(n_5444),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_5562)
);

BUFx2_ASAP7_75t_L g5563 ( 
.A(n_5416),
.Y(n_5563)
);

INVx6_ASAP7_75t_L g5564 ( 
.A(n_5360),
.Y(n_5564)
);

OAI22xp33_ASAP7_75t_L g5565 ( 
.A1(n_5407),
.A2(n_439),
.B1(n_436),
.B2(n_438),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5393),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_5465),
.Y(n_5567)
);

AOI22xp33_ASAP7_75t_L g5568 ( 
.A1(n_5417),
.A2(n_440),
.B1(n_438),
.B2(n_439),
.Y(n_5568)
);

AOI22xp33_ASAP7_75t_L g5569 ( 
.A1(n_5371),
.A2(n_442),
.B1(n_440),
.B2(n_441),
.Y(n_5569)
);

AOI22xp33_ASAP7_75t_L g5570 ( 
.A1(n_5419),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_5570)
);

CKINVDCx11_ASAP7_75t_R g5571 ( 
.A(n_5447),
.Y(n_5571)
);

AOI22xp33_ASAP7_75t_L g5572 ( 
.A1(n_5404),
.A2(n_447),
.B1(n_444),
.B2(n_446),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_5464),
.Y(n_5573)
);

AND2x2_ASAP7_75t_L g5574 ( 
.A(n_5405),
.B(n_5411),
.Y(n_5574)
);

AOI22xp33_ASAP7_75t_L g5575 ( 
.A1(n_5458),
.A2(n_450),
.B1(n_446),
.B2(n_448),
.Y(n_5575)
);

BUFx6f_ASAP7_75t_L g5576 ( 
.A(n_5399),
.Y(n_5576)
);

AOI22xp33_ASAP7_75t_L g5577 ( 
.A1(n_5468),
.A2(n_453),
.B1(n_451),
.B2(n_452),
.Y(n_5577)
);

OA21x2_ASAP7_75t_L g5578 ( 
.A1(n_5508),
.A2(n_5513),
.B(n_5529),
.Y(n_5578)
);

AND2x2_ASAP7_75t_L g5579 ( 
.A(n_5574),
.B(n_5418),
.Y(n_5579)
);

BUFx2_ASAP7_75t_L g5580 ( 
.A(n_5473),
.Y(n_5580)
);

AOI21xp5_ASAP7_75t_L g5581 ( 
.A1(n_5490),
.A2(n_5390),
.B(n_5403),
.Y(n_5581)
);

OAI22xp5_ASAP7_75t_L g5582 ( 
.A1(n_5482),
.A2(n_5439),
.B1(n_5451),
.B2(n_5431),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5502),
.Y(n_5583)
);

O2A1O1Ixp33_ASAP7_75t_L g5584 ( 
.A1(n_5556),
.A2(n_5461),
.B(n_5445),
.C(n_5428),
.Y(n_5584)
);

INVx1_ASAP7_75t_L g5585 ( 
.A(n_5532),
.Y(n_5585)
);

NAND2xp5_ASAP7_75t_L g5586 ( 
.A(n_5559),
.B(n_5430),
.Y(n_5586)
);

CKINVDCx14_ASAP7_75t_R g5587 ( 
.A(n_5485),
.Y(n_5587)
);

INVx1_ASAP7_75t_L g5588 ( 
.A(n_5524),
.Y(n_5588)
);

NAND2xp5_ASAP7_75t_L g5589 ( 
.A(n_5500),
.B(n_5437),
.Y(n_5589)
);

O2A1O1Ixp33_ASAP7_75t_L g5590 ( 
.A1(n_5504),
.A2(n_5479),
.B(n_5496),
.C(n_5511),
.Y(n_5590)
);

AND2x4_ASAP7_75t_L g5591 ( 
.A(n_5548),
.B(n_5422),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5507),
.Y(n_5592)
);

NAND2xp5_ASAP7_75t_L g5593 ( 
.A(n_5471),
.B(n_5449),
.Y(n_5593)
);

INVx2_ASAP7_75t_L g5594 ( 
.A(n_5558),
.Y(n_5594)
);

OR2x2_ASAP7_75t_L g5595 ( 
.A(n_5497),
.B(n_5469),
.Y(n_5595)
);

OAI22xp5_ASAP7_75t_L g5596 ( 
.A1(n_5519),
.A2(n_5446),
.B1(n_453),
.B2(n_451),
.Y(n_5596)
);

O2A1O1Ixp33_ASAP7_75t_L g5597 ( 
.A1(n_5547),
.A2(n_455),
.B(n_452),
.C(n_454),
.Y(n_5597)
);

AND2x2_ASAP7_75t_L g5598 ( 
.A(n_5560),
.B(n_456),
.Y(n_5598)
);

INVxp67_ASAP7_75t_L g5599 ( 
.A(n_5527),
.Y(n_5599)
);

AND2x4_ASAP7_75t_L g5600 ( 
.A(n_5555),
.B(n_456),
.Y(n_5600)
);

HB1xp67_ASAP7_75t_L g5601 ( 
.A(n_5478),
.Y(n_5601)
);

AND2x2_ASAP7_75t_L g5602 ( 
.A(n_5563),
.B(n_5506),
.Y(n_5602)
);

AOI21xp5_ASAP7_75t_L g5603 ( 
.A1(n_5521),
.A2(n_457),
.B(n_458),
.Y(n_5603)
);

AND2x2_ASAP7_75t_L g5604 ( 
.A(n_5498),
.B(n_457),
.Y(n_5604)
);

AND2x4_ASAP7_75t_L g5605 ( 
.A(n_5510),
.B(n_460),
.Y(n_5605)
);

BUFx6f_ASAP7_75t_L g5606 ( 
.A(n_5480),
.Y(n_5606)
);

AND2x2_ASAP7_75t_L g5607 ( 
.A(n_5545),
.B(n_460),
.Y(n_5607)
);

AOI21xp5_ASAP7_75t_SL g5608 ( 
.A1(n_5567),
.A2(n_461),
.B(n_462),
.Y(n_5608)
);

OAI22xp33_ASAP7_75t_L g5609 ( 
.A1(n_5481),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_5609)
);

OR2x2_ASAP7_75t_L g5610 ( 
.A(n_5573),
.B(n_463),
.Y(n_5610)
);

AND2x2_ASAP7_75t_L g5611 ( 
.A(n_5525),
.B(n_464),
.Y(n_5611)
);

OAI22xp5_ASAP7_75t_L g5612 ( 
.A1(n_5475),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_5612)
);

AND2x2_ASAP7_75t_L g5613 ( 
.A(n_5470),
.B(n_465),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5509),
.Y(n_5614)
);

AOI21xp5_ASAP7_75t_SL g5615 ( 
.A1(n_5551),
.A2(n_466),
.B(n_467),
.Y(n_5615)
);

AND2x2_ASAP7_75t_L g5616 ( 
.A(n_5495),
.B(n_467),
.Y(n_5616)
);

AOI22xp33_ASAP7_75t_SL g5617 ( 
.A1(n_5564),
.A2(n_473),
.B1(n_468),
.B2(n_471),
.Y(n_5617)
);

HB1xp67_ASAP7_75t_L g5618 ( 
.A(n_5566),
.Y(n_5618)
);

OA21x2_ASAP7_75t_L g5619 ( 
.A1(n_5484),
.A2(n_468),
.B(n_471),
.Y(n_5619)
);

INVx2_ASAP7_75t_SL g5620 ( 
.A(n_5546),
.Y(n_5620)
);

NAND2xp5_ASAP7_75t_L g5621 ( 
.A(n_5543),
.B(n_5477),
.Y(n_5621)
);

OR2x2_ASAP7_75t_L g5622 ( 
.A(n_5537),
.B(n_473),
.Y(n_5622)
);

NOR2xp33_ASAP7_75t_L g5623 ( 
.A(n_5474),
.B(n_474),
.Y(n_5623)
);

AOI21x1_ASAP7_75t_SL g5624 ( 
.A1(n_5505),
.A2(n_475),
.B(n_476),
.Y(n_5624)
);

OAI22xp5_ASAP7_75t_L g5625 ( 
.A1(n_5491),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5483),
.B(n_477),
.Y(n_5626)
);

CKINVDCx5p33_ASAP7_75t_R g5627 ( 
.A(n_5493),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_5472),
.B(n_478),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5488),
.Y(n_5629)
);

OR2x2_ASAP7_75t_L g5630 ( 
.A(n_5518),
.B(n_479),
.Y(n_5630)
);

OR2x2_ASAP7_75t_L g5631 ( 
.A(n_5520),
.B(n_479),
.Y(n_5631)
);

NAND2xp5_ASAP7_75t_L g5632 ( 
.A(n_5516),
.B(n_480),
.Y(n_5632)
);

AND2x2_ASAP7_75t_L g5633 ( 
.A(n_5540),
.B(n_481),
.Y(n_5633)
);

OA22x2_ASAP7_75t_L g5634 ( 
.A1(n_5557),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_5634)
);

BUFx12f_ASAP7_75t_L g5635 ( 
.A(n_5489),
.Y(n_5635)
);

AND2x2_ASAP7_75t_L g5636 ( 
.A(n_5501),
.B(n_483),
.Y(n_5636)
);

AND2x4_ASAP7_75t_L g5637 ( 
.A(n_5561),
.B(n_484),
.Y(n_5637)
);

O2A1O1Ixp5_ASAP7_75t_L g5638 ( 
.A1(n_5565),
.A2(n_486),
.B(n_484),
.C(n_485),
.Y(n_5638)
);

OAI22xp5_ASAP7_75t_L g5639 ( 
.A1(n_5515),
.A2(n_488),
.B1(n_485),
.B2(n_487),
.Y(n_5639)
);

NAND2xp5_ASAP7_75t_L g5640 ( 
.A(n_5517),
.B(n_487),
.Y(n_5640)
);

AOI21x1_ASAP7_75t_SL g5641 ( 
.A1(n_5539),
.A2(n_488),
.B(n_489),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_5534),
.Y(n_5642)
);

O2A1O1Ixp33_ASAP7_75t_L g5643 ( 
.A1(n_5553),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_5643)
);

AOI221xp5_ASAP7_75t_L g5644 ( 
.A1(n_5541),
.A2(n_494),
.B1(n_490),
.B2(n_492),
.C(n_495),
.Y(n_5644)
);

AND2x2_ASAP7_75t_L g5645 ( 
.A(n_5549),
.B(n_494),
.Y(n_5645)
);

OAI22xp5_ASAP7_75t_L g5646 ( 
.A1(n_5572),
.A2(n_498),
.B1(n_495),
.B2(n_497),
.Y(n_5646)
);

AND2x2_ASAP7_75t_L g5647 ( 
.A(n_5549),
.B(n_499),
.Y(n_5647)
);

OA21x2_ASAP7_75t_L g5648 ( 
.A1(n_5550),
.A2(n_5554),
.B(n_5523),
.Y(n_5648)
);

O2A1O1Ixp33_ASAP7_75t_L g5649 ( 
.A1(n_5530),
.A2(n_5577),
.B(n_5542),
.C(n_5544),
.Y(n_5649)
);

O2A1O1Ixp33_ASAP7_75t_L g5650 ( 
.A1(n_5569),
.A2(n_502),
.B(n_499),
.C(n_501),
.Y(n_5650)
);

OAI211xp5_ASAP7_75t_L g5651 ( 
.A1(n_5552),
.A2(n_503),
.B(n_501),
.C(n_502),
.Y(n_5651)
);

INVx1_ASAP7_75t_L g5652 ( 
.A(n_5576),
.Y(n_5652)
);

AND2x2_ASAP7_75t_L g5653 ( 
.A(n_5576),
.B(n_503),
.Y(n_5653)
);

AND2x2_ASAP7_75t_L g5654 ( 
.A(n_5503),
.B(n_504),
.Y(n_5654)
);

AOI21x1_ASAP7_75t_SL g5655 ( 
.A1(n_5494),
.A2(n_505),
.B(n_507),
.Y(n_5655)
);

NOR2xp67_ASAP7_75t_L g5656 ( 
.A(n_5492),
.B(n_505),
.Y(n_5656)
);

AND2x4_ASAP7_75t_L g5657 ( 
.A(n_5476),
.B(n_507),
.Y(n_5657)
);

O2A1O1Ixp33_ASAP7_75t_L g5658 ( 
.A1(n_5575),
.A2(n_511),
.B(n_509),
.C(n_510),
.Y(n_5658)
);

AND2x2_ASAP7_75t_L g5659 ( 
.A(n_5538),
.B(n_509),
.Y(n_5659)
);

INVx1_ASAP7_75t_SL g5660 ( 
.A(n_5571),
.Y(n_5660)
);

INVx1_ASAP7_75t_L g5661 ( 
.A(n_5601),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5585),
.Y(n_5662)
);

NAND2xp33_ASAP7_75t_L g5663 ( 
.A(n_5606),
.B(n_5486),
.Y(n_5663)
);

NAND2xp33_ASAP7_75t_SL g5664 ( 
.A(n_5606),
.B(n_5486),
.Y(n_5664)
);

INVx2_ASAP7_75t_L g5665 ( 
.A(n_5594),
.Y(n_5665)
);

NOR2xp33_ASAP7_75t_R g5666 ( 
.A(n_5587),
.B(n_5487),
.Y(n_5666)
);

AOI222xp33_ASAP7_75t_L g5667 ( 
.A1(n_5612),
.A2(n_5570),
.B1(n_5568),
.B2(n_5562),
.C1(n_5536),
.C2(n_5514),
.Y(n_5667)
);

AND2x2_ASAP7_75t_SL g5668 ( 
.A(n_5619),
.B(n_5535),
.Y(n_5668)
);

BUFx12f_ASAP7_75t_L g5669 ( 
.A(n_5635),
.Y(n_5669)
);

INVx2_ASAP7_75t_L g5670 ( 
.A(n_5629),
.Y(n_5670)
);

OAI21xp33_ASAP7_75t_L g5671 ( 
.A1(n_5581),
.A2(n_5590),
.B(n_5599),
.Y(n_5671)
);

INVx2_ASAP7_75t_L g5672 ( 
.A(n_5588),
.Y(n_5672)
);

INVx3_ASAP7_75t_L g5673 ( 
.A(n_5627),
.Y(n_5673)
);

OR2x6_ASAP7_75t_L g5674 ( 
.A(n_5608),
.B(n_5499),
.Y(n_5674)
);

INVx2_ASAP7_75t_L g5675 ( 
.A(n_5592),
.Y(n_5675)
);

NOR2xp67_ASAP7_75t_L g5676 ( 
.A(n_5656),
.B(n_5512),
.Y(n_5676)
);

NOR2xp33_ASAP7_75t_R g5677 ( 
.A(n_5660),
.B(n_5522),
.Y(n_5677)
);

AOI22xp33_ASAP7_75t_L g5678 ( 
.A1(n_5596),
.A2(n_5528),
.B1(n_5533),
.B2(n_5531),
.Y(n_5678)
);

INVxp67_ASAP7_75t_L g5679 ( 
.A(n_5618),
.Y(n_5679)
);

AND2x2_ASAP7_75t_L g5680 ( 
.A(n_5602),
.B(n_5526),
.Y(n_5680)
);

NOR3xp33_ASAP7_75t_SL g5681 ( 
.A(n_5609),
.B(n_510),
.C(n_512),
.Y(n_5681)
);

NAND2xp5_ASAP7_75t_L g5682 ( 
.A(n_5583),
.B(n_5535),
.Y(n_5682)
);

BUFx6f_ASAP7_75t_L g5683 ( 
.A(n_5657),
.Y(n_5683)
);

NAND2xp5_ASAP7_75t_L g5684 ( 
.A(n_5586),
.B(n_513),
.Y(n_5684)
);

NAND2xp33_ASAP7_75t_R g5685 ( 
.A(n_5636),
.B(n_514),
.Y(n_5685)
);

AND2x4_ASAP7_75t_L g5686 ( 
.A(n_5579),
.B(n_513),
.Y(n_5686)
);

HB1xp67_ASAP7_75t_L g5687 ( 
.A(n_5578),
.Y(n_5687)
);

CKINVDCx10_ASAP7_75t_R g5688 ( 
.A(n_5623),
.Y(n_5688)
);

CKINVDCx5p33_ASAP7_75t_R g5689 ( 
.A(n_5620),
.Y(n_5689)
);

OAI221xp5_ASAP7_75t_L g5690 ( 
.A1(n_5603),
.A2(n_516),
.B1(n_514),
.B2(n_515),
.C(n_517),
.Y(n_5690)
);

INVx1_ASAP7_75t_L g5691 ( 
.A(n_5614),
.Y(n_5691)
);

AOI22xp33_ASAP7_75t_L g5692 ( 
.A1(n_5634),
.A2(n_519),
.B1(n_517),
.B2(n_518),
.Y(n_5692)
);

NAND2xp5_ASAP7_75t_L g5693 ( 
.A(n_5593),
.B(n_520),
.Y(n_5693)
);

NAND2xp5_ASAP7_75t_L g5694 ( 
.A(n_5598),
.B(n_521),
.Y(n_5694)
);

INVx1_ASAP7_75t_L g5695 ( 
.A(n_5621),
.Y(n_5695)
);

CKINVDCx16_ASAP7_75t_R g5696 ( 
.A(n_5633),
.Y(n_5696)
);

NAND2xp5_ASAP7_75t_L g5697 ( 
.A(n_5611),
.B(n_521),
.Y(n_5697)
);

NAND2xp5_ASAP7_75t_L g5698 ( 
.A(n_5630),
.B(n_522),
.Y(n_5698)
);

INVx2_ASAP7_75t_L g5699 ( 
.A(n_5642),
.Y(n_5699)
);

AND2x2_ASAP7_75t_L g5700 ( 
.A(n_5591),
.B(n_5580),
.Y(n_5700)
);

INVx5_ASAP7_75t_L g5701 ( 
.A(n_5659),
.Y(n_5701)
);

AND2x2_ASAP7_75t_L g5702 ( 
.A(n_5652),
.B(n_523),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_5631),
.B(n_523),
.Y(n_5703)
);

BUFx2_ASAP7_75t_L g5704 ( 
.A(n_5605),
.Y(n_5704)
);

INVx1_ASAP7_75t_L g5705 ( 
.A(n_5632),
.Y(n_5705)
);

CKINVDCx20_ASAP7_75t_R g5706 ( 
.A(n_5604),
.Y(n_5706)
);

NAND2xp33_ASAP7_75t_R g5707 ( 
.A(n_5648),
.B(n_525),
.Y(n_5707)
);

NOR2xp33_ASAP7_75t_R g5708 ( 
.A(n_5654),
.B(n_1817),
.Y(n_5708)
);

OAI21xp33_ASAP7_75t_L g5709 ( 
.A1(n_5615),
.A2(n_524),
.B(n_527),
.Y(n_5709)
);

INVx2_ASAP7_75t_L g5710 ( 
.A(n_5595),
.Y(n_5710)
);

NAND2xp33_ASAP7_75t_R g5711 ( 
.A(n_5600),
.B(n_527),
.Y(n_5711)
);

BUFx2_ASAP7_75t_L g5712 ( 
.A(n_5637),
.Y(n_5712)
);

OR2x2_ASAP7_75t_L g5713 ( 
.A(n_5589),
.B(n_5610),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5640),
.Y(n_5714)
);

NAND2xp33_ASAP7_75t_R g5715 ( 
.A(n_5653),
.B(n_528),
.Y(n_5715)
);

NAND2xp33_ASAP7_75t_R g5716 ( 
.A(n_5607),
.B(n_528),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_5626),
.Y(n_5717)
);

BUFx3_ASAP7_75t_L g5718 ( 
.A(n_5645),
.Y(n_5718)
);

NAND2xp5_ASAP7_75t_L g5719 ( 
.A(n_5628),
.B(n_524),
.Y(n_5719)
);

NOR2xp33_ASAP7_75t_R g5720 ( 
.A(n_5647),
.B(n_1820),
.Y(n_5720)
);

BUFx3_ASAP7_75t_L g5721 ( 
.A(n_5613),
.Y(n_5721)
);

INVx2_ASAP7_75t_SL g5722 ( 
.A(n_5622),
.Y(n_5722)
);

CKINVDCx5p33_ASAP7_75t_R g5723 ( 
.A(n_5616),
.Y(n_5723)
);

CKINVDCx5p33_ASAP7_75t_R g5724 ( 
.A(n_5582),
.Y(n_5724)
);

INVx2_ASAP7_75t_L g5725 ( 
.A(n_5638),
.Y(n_5725)
);

INVx2_ASAP7_75t_L g5726 ( 
.A(n_5639),
.Y(n_5726)
);

CKINVDCx16_ASAP7_75t_R g5727 ( 
.A(n_5625),
.Y(n_5727)
);

AND2x2_ASAP7_75t_L g5728 ( 
.A(n_5584),
.B(n_5649),
.Y(n_5728)
);

AND2x4_ASAP7_75t_L g5729 ( 
.A(n_5624),
.B(n_529),
.Y(n_5729)
);

OR2x6_ASAP7_75t_L g5730 ( 
.A(n_5597),
.B(n_529),
.Y(n_5730)
);

INVx1_ASAP7_75t_L g5731 ( 
.A(n_5643),
.Y(n_5731)
);

AND2x2_ASAP7_75t_L g5732 ( 
.A(n_5617),
.B(n_530),
.Y(n_5732)
);

AND2x2_ASAP7_75t_L g5733 ( 
.A(n_5646),
.B(n_530),
.Y(n_5733)
);

HB1xp67_ASAP7_75t_L g5734 ( 
.A(n_5644),
.Y(n_5734)
);

NAND2xp33_ASAP7_75t_R g5735 ( 
.A(n_5655),
.B(n_532),
.Y(n_5735)
);

AND2x2_ASAP7_75t_L g5736 ( 
.A(n_5658),
.B(n_531),
.Y(n_5736)
);

NOR3xp33_ASAP7_75t_SL g5737 ( 
.A(n_5651),
.B(n_532),
.C(n_533),
.Y(n_5737)
);

INVx2_ASAP7_75t_L g5738 ( 
.A(n_5641),
.Y(n_5738)
);

OAI22xp5_ASAP7_75t_L g5739 ( 
.A1(n_5650),
.A2(n_535),
.B1(n_533),
.B2(n_534),
.Y(n_5739)
);

NOR2x1p5_ASAP7_75t_L g5740 ( 
.A(n_5635),
.B(n_534),
.Y(n_5740)
);

INVx3_ASAP7_75t_L g5741 ( 
.A(n_5606),
.Y(n_5741)
);

AND2x2_ASAP7_75t_L g5742 ( 
.A(n_5602),
.B(n_535),
.Y(n_5742)
);

INVx1_ASAP7_75t_L g5743 ( 
.A(n_5601),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5601),
.Y(n_5744)
);

INVx2_ASAP7_75t_SL g5745 ( 
.A(n_5606),
.Y(n_5745)
);

AND2x2_ASAP7_75t_L g5746 ( 
.A(n_5602),
.B(n_536),
.Y(n_5746)
);

AND2x2_ASAP7_75t_L g5747 ( 
.A(n_5602),
.B(n_536),
.Y(n_5747)
);

AND2x4_ASAP7_75t_L g5748 ( 
.A(n_5579),
.B(n_537),
.Y(n_5748)
);

NAND2xp5_ASAP7_75t_L g5749 ( 
.A(n_5599),
.B(n_537),
.Y(n_5749)
);

INVx1_ASAP7_75t_L g5750 ( 
.A(n_5601),
.Y(n_5750)
);

INVx5_ASAP7_75t_L g5751 ( 
.A(n_5635),
.Y(n_5751)
);

INVx2_ASAP7_75t_L g5752 ( 
.A(n_5594),
.Y(n_5752)
);

OR2x6_ASAP7_75t_L g5753 ( 
.A(n_5606),
.B(n_538),
.Y(n_5753)
);

INVx2_ASAP7_75t_L g5754 ( 
.A(n_5594),
.Y(n_5754)
);

OR2x2_ASAP7_75t_L g5755 ( 
.A(n_5586),
.B(n_538),
.Y(n_5755)
);

AND2x4_ASAP7_75t_L g5756 ( 
.A(n_5579),
.B(n_540),
.Y(n_5756)
);

BUFx6f_ASAP7_75t_L g5757 ( 
.A(n_5606),
.Y(n_5757)
);

NOR2xp33_ASAP7_75t_R g5758 ( 
.A(n_5587),
.B(n_1814),
.Y(n_5758)
);

CKINVDCx16_ASAP7_75t_R g5759 ( 
.A(n_5587),
.Y(n_5759)
);

AND2x2_ASAP7_75t_L g5760 ( 
.A(n_5602),
.B(n_540),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5601),
.Y(n_5761)
);

OAI21xp5_ASAP7_75t_SL g5762 ( 
.A1(n_5590),
.A2(n_541),
.B(n_542),
.Y(n_5762)
);

INVxp67_ASAP7_75t_L g5763 ( 
.A(n_5618),
.Y(n_5763)
);

NAND2xp33_ASAP7_75t_R g5764 ( 
.A(n_5627),
.B(n_542),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5594),
.Y(n_5765)
);

INVx2_ASAP7_75t_L g5766 ( 
.A(n_5594),
.Y(n_5766)
);

INVx2_ASAP7_75t_L g5767 ( 
.A(n_5594),
.Y(n_5767)
);

OR2x6_ASAP7_75t_L g5768 ( 
.A(n_5606),
.B(n_541),
.Y(n_5768)
);

NOR3xp33_ASAP7_75t_SL g5769 ( 
.A(n_5627),
.B(n_543),
.C(n_544),
.Y(n_5769)
);

INVx1_ASAP7_75t_L g5770 ( 
.A(n_5601),
.Y(n_5770)
);

OR2x2_ASAP7_75t_L g5771 ( 
.A(n_5586),
.B(n_543),
.Y(n_5771)
);

BUFx3_ASAP7_75t_L g5772 ( 
.A(n_5606),
.Y(n_5772)
);

NOR2xp33_ASAP7_75t_R g5773 ( 
.A(n_5587),
.B(n_1819),
.Y(n_5773)
);

AOI22xp33_ASAP7_75t_L g5774 ( 
.A1(n_5619),
.A2(n_547),
.B1(n_544),
.B2(n_545),
.Y(n_5774)
);

OR2x6_ASAP7_75t_L g5775 ( 
.A(n_5606),
.B(n_545),
.Y(n_5775)
);

CKINVDCx5p33_ASAP7_75t_R g5776 ( 
.A(n_5587),
.Y(n_5776)
);

AOI22xp33_ASAP7_75t_SL g5777 ( 
.A1(n_5578),
.A2(n_555),
.B1(n_564),
.B2(n_547),
.Y(n_5777)
);

AND2x2_ASAP7_75t_L g5778 ( 
.A(n_5602),
.B(n_548),
.Y(n_5778)
);

BUFx10_ASAP7_75t_L g5779 ( 
.A(n_5606),
.Y(n_5779)
);

AND2x2_ASAP7_75t_L g5780 ( 
.A(n_5602),
.B(n_548),
.Y(n_5780)
);

BUFx3_ASAP7_75t_L g5781 ( 
.A(n_5606),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5601),
.Y(n_5782)
);

HB1xp67_ASAP7_75t_L g5783 ( 
.A(n_5699),
.Y(n_5783)
);

AOI33xp33_ASAP7_75t_L g5784 ( 
.A1(n_5728),
.A2(n_551),
.A3(n_553),
.B1(n_549),
.B2(n_550),
.B3(n_552),
.Y(n_5784)
);

OAI21x1_ASAP7_75t_L g5785 ( 
.A1(n_5687),
.A2(n_549),
.B(n_551),
.Y(n_5785)
);

INVx1_ASAP7_75t_L g5786 ( 
.A(n_5662),
.Y(n_5786)
);

INVx2_ASAP7_75t_L g5787 ( 
.A(n_5710),
.Y(n_5787)
);

OAI22xp33_ASAP7_75t_L g5788 ( 
.A1(n_5727),
.A2(n_555),
.B1(n_553),
.B2(n_554),
.Y(n_5788)
);

AND2x2_ASAP7_75t_L g5789 ( 
.A(n_5700),
.B(n_556),
.Y(n_5789)
);

INVxp67_ASAP7_75t_SL g5790 ( 
.A(n_5711),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5691),
.Y(n_5791)
);

INVx2_ASAP7_75t_L g5792 ( 
.A(n_5665),
.Y(n_5792)
);

OA21x2_ASAP7_75t_L g5793 ( 
.A1(n_5671),
.A2(n_5724),
.B(n_5679),
.Y(n_5793)
);

INVx1_ASAP7_75t_L g5794 ( 
.A(n_5672),
.Y(n_5794)
);

INVx3_ASAP7_75t_L g5795 ( 
.A(n_5759),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5675),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5752),
.Y(n_5797)
);

NAND2xp5_ASAP7_75t_L g5798 ( 
.A(n_5695),
.B(n_556),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5661),
.Y(n_5799)
);

INVx2_ASAP7_75t_L g5800 ( 
.A(n_5754),
.Y(n_5800)
);

INVx4_ASAP7_75t_L g5801 ( 
.A(n_5751),
.Y(n_5801)
);

INVx2_ASAP7_75t_L g5802 ( 
.A(n_5765),
.Y(n_5802)
);

OA21x2_ASAP7_75t_L g5803 ( 
.A1(n_5763),
.A2(n_5744),
.B(n_5743),
.Y(n_5803)
);

INVx2_ASAP7_75t_L g5804 ( 
.A(n_5766),
.Y(n_5804)
);

OR2x2_ASAP7_75t_L g5805 ( 
.A(n_5750),
.B(n_558),
.Y(n_5805)
);

OR2x2_ASAP7_75t_L g5806 ( 
.A(n_5761),
.B(n_558),
.Y(n_5806)
);

INVx2_ASAP7_75t_L g5807 ( 
.A(n_5767),
.Y(n_5807)
);

INVx2_ASAP7_75t_L g5808 ( 
.A(n_5670),
.Y(n_5808)
);

INVx1_ASAP7_75t_SL g5809 ( 
.A(n_5688),
.Y(n_5809)
);

AOI21xp5_ASAP7_75t_SL g5810 ( 
.A1(n_5674),
.A2(n_5709),
.B(n_5676),
.Y(n_5810)
);

INVx1_ASAP7_75t_L g5811 ( 
.A(n_5770),
.Y(n_5811)
);

OA21x2_ASAP7_75t_L g5812 ( 
.A1(n_5782),
.A2(n_1817),
.B(n_1816),
.Y(n_5812)
);

INVx1_ASAP7_75t_L g5813 ( 
.A(n_5705),
.Y(n_5813)
);

OA21x2_ASAP7_75t_L g5814 ( 
.A1(n_5704),
.A2(n_1820),
.B(n_1818),
.Y(n_5814)
);

INVx1_ASAP7_75t_L g5815 ( 
.A(n_5714),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5717),
.Y(n_5816)
);

OA21x2_ASAP7_75t_L g5817 ( 
.A1(n_5712),
.A2(n_1822),
.B(n_1821),
.Y(n_5817)
);

OA21x2_ASAP7_75t_L g5818 ( 
.A1(n_5689),
.A2(n_5693),
.B(n_5682),
.Y(n_5818)
);

INVx2_ASAP7_75t_L g5819 ( 
.A(n_5721),
.Y(n_5819)
);

AND2x2_ASAP7_75t_L g5820 ( 
.A(n_5696),
.B(n_559),
.Y(n_5820)
);

OR2x6_ASAP7_75t_L g5821 ( 
.A(n_5669),
.B(n_560),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5749),
.Y(n_5822)
);

OA21x2_ASAP7_75t_L g5823 ( 
.A1(n_5678),
.A2(n_1824),
.B(n_1822),
.Y(n_5823)
);

OR2x2_ASAP7_75t_L g5824 ( 
.A(n_5713),
.B(n_560),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_5722),
.Y(n_5825)
);

AND2x2_ASAP7_75t_L g5826 ( 
.A(n_5680),
.B(n_561),
.Y(n_5826)
);

INVx2_ASAP7_75t_L g5827 ( 
.A(n_5668),
.Y(n_5827)
);

INVxp67_ASAP7_75t_L g5828 ( 
.A(n_5764),
.Y(n_5828)
);

AOI22xp5_ASAP7_75t_L g5829 ( 
.A1(n_5762),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.Y(n_5829)
);

INVx2_ASAP7_75t_L g5830 ( 
.A(n_5718),
.Y(n_5830)
);

OA21x2_ASAP7_75t_L g5831 ( 
.A1(n_5684),
.A2(n_562),
.B(n_563),
.Y(n_5831)
);

INVx1_ASAP7_75t_L g5832 ( 
.A(n_5755),
.Y(n_5832)
);

INVxp67_ASAP7_75t_L g5833 ( 
.A(n_5716),
.Y(n_5833)
);

INVx1_ASAP7_75t_L g5834 ( 
.A(n_5771),
.Y(n_5834)
);

OAI21xp5_ASAP7_75t_L g5835 ( 
.A1(n_5777),
.A2(n_5734),
.B(n_5725),
.Y(n_5835)
);

OA21x2_ASAP7_75t_L g5836 ( 
.A1(n_5723),
.A2(n_1804),
.B(n_1803),
.Y(n_5836)
);

OA21x2_ASAP7_75t_L g5837 ( 
.A1(n_5742),
.A2(n_1804),
.B(n_1803),
.Y(n_5837)
);

AND2x2_ASAP7_75t_L g5838 ( 
.A(n_5746),
.B(n_5747),
.Y(n_5838)
);

INVx1_ASAP7_75t_L g5839 ( 
.A(n_5726),
.Y(n_5839)
);

INVx1_ASAP7_75t_L g5840 ( 
.A(n_5731),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5698),
.Y(n_5841)
);

INVx1_ASAP7_75t_L g5842 ( 
.A(n_5703),
.Y(n_5842)
);

AND2x4_ASAP7_75t_L g5843 ( 
.A(n_5701),
.B(n_566),
.Y(n_5843)
);

AO21x2_ASAP7_75t_L g5844 ( 
.A1(n_5758),
.A2(n_5773),
.B(n_5708),
.Y(n_5844)
);

INVx1_ASAP7_75t_L g5845 ( 
.A(n_5702),
.Y(n_5845)
);

INVx2_ASAP7_75t_L g5846 ( 
.A(n_5701),
.Y(n_5846)
);

INVx1_ASAP7_75t_SL g5847 ( 
.A(n_5677),
.Y(n_5847)
);

INVx2_ASAP7_75t_L g5848 ( 
.A(n_5760),
.Y(n_5848)
);

INVx1_ASAP7_75t_L g5849 ( 
.A(n_5778),
.Y(n_5849)
);

INVx1_ASAP7_75t_L g5850 ( 
.A(n_5780),
.Y(n_5850)
);

INVx2_ASAP7_75t_L g5851 ( 
.A(n_5683),
.Y(n_5851)
);

AND2x4_ASAP7_75t_SL g5852 ( 
.A(n_5779),
.B(n_568),
.Y(n_5852)
);

OR2x2_ASAP7_75t_L g5853 ( 
.A(n_5697),
.B(n_568),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_5683),
.B(n_569),
.Y(n_5854)
);

NAND2xp5_ASAP7_75t_L g5855 ( 
.A(n_5719),
.B(n_570),
.Y(n_5855)
);

AO21x2_ASAP7_75t_L g5856 ( 
.A1(n_5720),
.A2(n_5694),
.B(n_5707),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5738),
.Y(n_5857)
);

NOR2xp33_ASAP7_75t_L g5858 ( 
.A(n_5751),
.B(n_570),
.Y(n_5858)
);

INVx1_ASAP7_75t_L g5859 ( 
.A(n_5736),
.Y(n_5859)
);

NOR2xp33_ASAP7_75t_L g5860 ( 
.A(n_5776),
.B(n_571),
.Y(n_5860)
);

OAI21xp5_ASAP7_75t_L g5861 ( 
.A1(n_5730),
.A2(n_5774),
.B(n_5681),
.Y(n_5861)
);

AND2x2_ASAP7_75t_L g5862 ( 
.A(n_5673),
.B(n_571),
.Y(n_5862)
);

AO21x2_ASAP7_75t_L g5863 ( 
.A1(n_5666),
.A2(n_572),
.B(n_573),
.Y(n_5863)
);

OAI21xp5_ASAP7_75t_L g5864 ( 
.A1(n_5730),
.A2(n_573),
.B(n_574),
.Y(n_5864)
);

BUFx2_ASAP7_75t_L g5865 ( 
.A(n_5664),
.Y(n_5865)
);

OA21x2_ASAP7_75t_L g5866 ( 
.A1(n_5745),
.A2(n_1821),
.B(n_1815),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_5706),
.Y(n_5867)
);

HB1xp67_ASAP7_75t_L g5868 ( 
.A(n_5686),
.Y(n_5868)
);

NOR2xp33_ASAP7_75t_L g5869 ( 
.A(n_5757),
.B(n_574),
.Y(n_5869)
);

INVx2_ASAP7_75t_L g5870 ( 
.A(n_5748),
.Y(n_5870)
);

OA21x2_ASAP7_75t_L g5871 ( 
.A1(n_5756),
.A2(n_5692),
.B(n_5769),
.Y(n_5871)
);

OR2x2_ASAP7_75t_L g5872 ( 
.A(n_5674),
.B(n_575),
.Y(n_5872)
);

CKINVDCx5p33_ASAP7_75t_R g5873 ( 
.A(n_5685),
.Y(n_5873)
);

INVx2_ASAP7_75t_L g5874 ( 
.A(n_5741),
.Y(n_5874)
);

INVx1_ASAP7_75t_L g5875 ( 
.A(n_5733),
.Y(n_5875)
);

INVx2_ASAP7_75t_L g5876 ( 
.A(n_5772),
.Y(n_5876)
);

OR2x6_ASAP7_75t_L g5877 ( 
.A(n_5757),
.B(n_5781),
.Y(n_5877)
);

BUFx6f_ASAP7_75t_L g5878 ( 
.A(n_5753),
.Y(n_5878)
);

NAND2xp5_ASAP7_75t_L g5879 ( 
.A(n_5732),
.B(n_576),
.Y(n_5879)
);

AND2x2_ASAP7_75t_L g5880 ( 
.A(n_5663),
.B(n_576),
.Y(n_5880)
);

OAI21x1_ASAP7_75t_L g5881 ( 
.A1(n_5740),
.A2(n_577),
.B(n_578),
.Y(n_5881)
);

HB1xp67_ASAP7_75t_L g5882 ( 
.A(n_5753),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5729),
.Y(n_5883)
);

AOI22xp33_ASAP7_75t_L g5884 ( 
.A1(n_5667),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5739),
.Y(n_5885)
);

INVx1_ASAP7_75t_L g5886 ( 
.A(n_5768),
.Y(n_5886)
);

OR2x6_ASAP7_75t_L g5887 ( 
.A(n_5768),
.B(n_579),
.Y(n_5887)
);

NAND2xp5_ASAP7_75t_L g5888 ( 
.A(n_5737),
.B(n_581),
.Y(n_5888)
);

OAI22xp5_ASAP7_75t_L g5889 ( 
.A1(n_5775),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_5889)
);

AND2x2_ASAP7_75t_L g5890 ( 
.A(n_5775),
.B(n_5715),
.Y(n_5890)
);

INVx2_ASAP7_75t_L g5891 ( 
.A(n_5690),
.Y(n_5891)
);

AND2x4_ASAP7_75t_L g5892 ( 
.A(n_5735),
.B(n_583),
.Y(n_5892)
);

AND2x4_ASAP7_75t_L g5893 ( 
.A(n_5718),
.B(n_584),
.Y(n_5893)
);

OR2x6_ASAP7_75t_L g5894 ( 
.A(n_5669),
.B(n_585),
.Y(n_5894)
);

INVx2_ASAP7_75t_L g5895 ( 
.A(n_5710),
.Y(n_5895)
);

INVx3_ASAP7_75t_L g5896 ( 
.A(n_5759),
.Y(n_5896)
);

OR2x6_ASAP7_75t_L g5897 ( 
.A(n_5669),
.B(n_585),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5662),
.Y(n_5898)
);

AO21x1_ASAP7_75t_L g5899 ( 
.A1(n_5728),
.A2(n_586),
.B(n_587),
.Y(n_5899)
);

OR2x2_ASAP7_75t_L g5900 ( 
.A(n_5695),
.B(n_588),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5710),
.Y(n_5901)
);

OA21x2_ASAP7_75t_L g5902 ( 
.A1(n_5671),
.A2(n_1813),
.B(n_1811),
.Y(n_5902)
);

AOI21x1_ASAP7_75t_L g5903 ( 
.A1(n_5687),
.A2(n_588),
.B(n_589),
.Y(n_5903)
);

BUFx2_ASAP7_75t_L g5904 ( 
.A(n_5666),
.Y(n_5904)
);

AND2x2_ASAP7_75t_L g5905 ( 
.A(n_5700),
.B(n_590),
.Y(n_5905)
);

INVx1_ASAP7_75t_L g5906 ( 
.A(n_5662),
.Y(n_5906)
);

AO21x2_ASAP7_75t_L g5907 ( 
.A1(n_5687),
.A2(n_590),
.B(n_591),
.Y(n_5907)
);

INVx2_ASAP7_75t_L g5908 ( 
.A(n_5710),
.Y(n_5908)
);

NAND2xp5_ASAP7_75t_L g5909 ( 
.A(n_5671),
.B(n_591),
.Y(n_5909)
);

INVx2_ASAP7_75t_L g5910 ( 
.A(n_5710),
.Y(n_5910)
);

OR2x2_ASAP7_75t_L g5911 ( 
.A(n_5695),
.B(n_592),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5662),
.Y(n_5912)
);

INVx1_ASAP7_75t_L g5913 ( 
.A(n_5662),
.Y(n_5913)
);

AO21x2_ASAP7_75t_L g5914 ( 
.A1(n_5687),
.A2(n_592),
.B(n_593),
.Y(n_5914)
);

INVx2_ASAP7_75t_L g5915 ( 
.A(n_5710),
.Y(n_5915)
);

INVx1_ASAP7_75t_L g5916 ( 
.A(n_5662),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5662),
.Y(n_5917)
);

INVx3_ASAP7_75t_L g5918 ( 
.A(n_5759),
.Y(n_5918)
);

INVx2_ASAP7_75t_L g5919 ( 
.A(n_5710),
.Y(n_5919)
);

INVx3_ASAP7_75t_L g5920 ( 
.A(n_5759),
.Y(n_5920)
);

AND2x2_ASAP7_75t_L g5921 ( 
.A(n_5700),
.B(n_593),
.Y(n_5921)
);

INVx2_ASAP7_75t_L g5922 ( 
.A(n_5710),
.Y(n_5922)
);

AOI211xp5_ASAP7_75t_L g5923 ( 
.A1(n_5762),
.A2(n_596),
.B(n_594),
.C(n_595),
.Y(n_5923)
);

HB1xp67_ASAP7_75t_L g5924 ( 
.A(n_5699),
.Y(n_5924)
);

AND2x2_ASAP7_75t_L g5925 ( 
.A(n_5700),
.B(n_595),
.Y(n_5925)
);

AND2x2_ASAP7_75t_L g5926 ( 
.A(n_5700),
.B(n_597),
.Y(n_5926)
);

BUFx6f_ASAP7_75t_L g5927 ( 
.A(n_5669),
.Y(n_5927)
);

INVx1_ASAP7_75t_L g5928 ( 
.A(n_5662),
.Y(n_5928)
);

AOI22xp33_ASAP7_75t_L g5929 ( 
.A1(n_5734),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5710),
.Y(n_5930)
);

AND2x2_ASAP7_75t_L g5931 ( 
.A(n_5700),
.B(n_598),
.Y(n_5931)
);

INVx2_ASAP7_75t_L g5932 ( 
.A(n_5710),
.Y(n_5932)
);

AND2x2_ASAP7_75t_L g5933 ( 
.A(n_5700),
.B(n_600),
.Y(n_5933)
);

INVx2_ASAP7_75t_L g5934 ( 
.A(n_5710),
.Y(n_5934)
);

OAI21x1_ASAP7_75t_L g5935 ( 
.A1(n_5687),
.A2(n_601),
.B(n_602),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5710),
.Y(n_5936)
);

AO21x2_ASAP7_75t_L g5937 ( 
.A1(n_5687),
.A2(n_601),
.B(n_603),
.Y(n_5937)
);

BUFx3_ASAP7_75t_L g5938 ( 
.A(n_5669),
.Y(n_5938)
);

AND2x2_ASAP7_75t_L g5939 ( 
.A(n_5700),
.B(n_604),
.Y(n_5939)
);

OA21x2_ASAP7_75t_L g5940 ( 
.A1(n_5671),
.A2(n_1826),
.B(n_1813),
.Y(n_5940)
);

AND2x2_ASAP7_75t_L g5941 ( 
.A(n_5700),
.B(n_604),
.Y(n_5941)
);

OA21x2_ASAP7_75t_L g5942 ( 
.A1(n_5671),
.A2(n_1828),
.B(n_1827),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5662),
.Y(n_5943)
);

AO21x2_ASAP7_75t_L g5944 ( 
.A1(n_5687),
.A2(n_605),
.B(n_606),
.Y(n_5944)
);

INVx2_ASAP7_75t_L g5945 ( 
.A(n_5710),
.Y(n_5945)
);

OR2x2_ASAP7_75t_L g5946 ( 
.A(n_5840),
.B(n_1828),
.Y(n_5946)
);

NAND2x1_ASAP7_75t_L g5947 ( 
.A(n_5865),
.B(n_606),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_5795),
.Y(n_5948)
);

BUFx2_ASAP7_75t_L g5949 ( 
.A(n_5896),
.Y(n_5949)
);

HB1xp67_ASAP7_75t_L g5950 ( 
.A(n_5803),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5786),
.Y(n_5951)
);

BUFx2_ASAP7_75t_L g5952 ( 
.A(n_5918),
.Y(n_5952)
);

BUFx4f_ASAP7_75t_SL g5953 ( 
.A(n_5809),
.Y(n_5953)
);

AND2x4_ASAP7_75t_L g5954 ( 
.A(n_5920),
.B(n_605),
.Y(n_5954)
);

OAI22xp5_ASAP7_75t_L g5955 ( 
.A1(n_5793),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.Y(n_5955)
);

AO22x1_ASAP7_75t_L g5956 ( 
.A1(n_5892),
.A2(n_611),
.B1(n_609),
.B2(n_610),
.Y(n_5956)
);

INVx2_ASAP7_75t_L g5957 ( 
.A(n_5882),
.Y(n_5957)
);

INVx1_ASAP7_75t_L g5958 ( 
.A(n_5791),
.Y(n_5958)
);

NOR2x1_ASAP7_75t_L g5959 ( 
.A(n_5810),
.B(n_613),
.Y(n_5959)
);

NAND2xp5_ASAP7_75t_L g5960 ( 
.A(n_5907),
.B(n_614),
.Y(n_5960)
);

AND2x2_ASAP7_75t_L g5961 ( 
.A(n_5838),
.B(n_614),
.Y(n_5961)
);

AOI22xp33_ASAP7_75t_L g5962 ( 
.A1(n_5856),
.A2(n_617),
.B1(n_615),
.B2(n_616),
.Y(n_5962)
);

OR2x2_ASAP7_75t_L g5963 ( 
.A(n_5839),
.B(n_1802),
.Y(n_5963)
);

NAND2xp5_ASAP7_75t_L g5964 ( 
.A(n_5914),
.B(n_5937),
.Y(n_5964)
);

AND2x2_ASAP7_75t_L g5965 ( 
.A(n_5868),
.B(n_615),
.Y(n_5965)
);

AND2x2_ASAP7_75t_L g5966 ( 
.A(n_5904),
.B(n_616),
.Y(n_5966)
);

HB1xp67_ASAP7_75t_L g5967 ( 
.A(n_5812),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5818),
.B(n_617),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5824),
.B(n_1809),
.Y(n_5969)
);

INVx1_ASAP7_75t_L g5970 ( 
.A(n_5898),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5906),
.Y(n_5971)
);

OAI22xp5_ASAP7_75t_L g5972 ( 
.A1(n_5859),
.A2(n_620),
.B1(n_618),
.B2(n_619),
.Y(n_5972)
);

AND2x2_ASAP7_75t_L g5973 ( 
.A(n_5819),
.B(n_619),
.Y(n_5973)
);

INVx2_ASAP7_75t_L g5974 ( 
.A(n_5866),
.Y(n_5974)
);

INVx5_ASAP7_75t_L g5975 ( 
.A(n_5927),
.Y(n_5975)
);

INVx1_ASAP7_75t_L g5976 ( 
.A(n_5912),
.Y(n_5976)
);

INVx1_ASAP7_75t_L g5977 ( 
.A(n_5913),
.Y(n_5977)
);

INVx2_ASAP7_75t_L g5978 ( 
.A(n_5848),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5916),
.Y(n_5979)
);

INVx1_ASAP7_75t_L g5980 ( 
.A(n_5917),
.Y(n_5980)
);

AOI22xp5_ASAP7_75t_L g5981 ( 
.A1(n_5899),
.A2(n_622),
.B1(n_620),
.B2(n_621),
.Y(n_5981)
);

INVx1_ASAP7_75t_SL g5982 ( 
.A(n_5847),
.Y(n_5982)
);

BUFx3_ASAP7_75t_L g5983 ( 
.A(n_5927),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5928),
.Y(n_5984)
);

BUFx2_ASAP7_75t_L g5985 ( 
.A(n_5877),
.Y(n_5985)
);

NAND2xp5_ASAP7_75t_L g5986 ( 
.A(n_5944),
.B(n_623),
.Y(n_5986)
);

BUFx2_ASAP7_75t_L g5987 ( 
.A(n_5801),
.Y(n_5987)
);

AND2x2_ASAP7_75t_L g5988 ( 
.A(n_5874),
.B(n_625),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5817),
.Y(n_5989)
);

INVx1_ASAP7_75t_L g5990 ( 
.A(n_5943),
.Y(n_5990)
);

INVx1_ASAP7_75t_L g5991 ( 
.A(n_5813),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_5846),
.B(n_626),
.Y(n_5992)
);

AND2x2_ASAP7_75t_L g5993 ( 
.A(n_5857),
.B(n_627),
.Y(n_5993)
);

NOR2x1_ASAP7_75t_SL g5994 ( 
.A(n_5863),
.B(n_628),
.Y(n_5994)
);

INVx1_ASAP7_75t_L g5995 ( 
.A(n_5815),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5816),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5814),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5799),
.Y(n_5998)
);

OR2x2_ASAP7_75t_L g5999 ( 
.A(n_5822),
.B(n_5841),
.Y(n_5999)
);

INVxp67_ASAP7_75t_SL g6000 ( 
.A(n_5828),
.Y(n_6000)
);

INVx1_ASAP7_75t_L g6001 ( 
.A(n_5811),
.Y(n_6001)
);

AOI22xp33_ASAP7_75t_L g6002 ( 
.A1(n_5790),
.A2(n_630),
.B1(n_628),
.B2(n_629),
.Y(n_6002)
);

NAND2xp5_ASAP7_75t_L g6003 ( 
.A(n_5832),
.B(n_629),
.Y(n_6003)
);

AND2x4_ASAP7_75t_L g6004 ( 
.A(n_5867),
.B(n_630),
.Y(n_6004)
);

INVxp67_ASAP7_75t_SL g6005 ( 
.A(n_5902),
.Y(n_6005)
);

OR2x2_ASAP7_75t_L g6006 ( 
.A(n_5842),
.B(n_1801),
.Y(n_6006)
);

OR2x2_ASAP7_75t_L g6007 ( 
.A(n_5825),
.B(n_1801),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5783),
.Y(n_6008)
);

AND2x2_ASAP7_75t_L g6009 ( 
.A(n_5849),
.B(n_631),
.Y(n_6009)
);

INVx2_ASAP7_75t_SL g6010 ( 
.A(n_5938),
.Y(n_6010)
);

OR2x2_ASAP7_75t_L g6011 ( 
.A(n_5834),
.B(n_1806),
.Y(n_6011)
);

AND2x2_ASAP7_75t_L g6012 ( 
.A(n_5850),
.B(n_5851),
.Y(n_6012)
);

AND2x2_ASAP7_75t_L g6013 ( 
.A(n_5876),
.B(n_632),
.Y(n_6013)
);

INVx1_ASAP7_75t_L g6014 ( 
.A(n_5924),
.Y(n_6014)
);

INVxp67_ASAP7_75t_L g6015 ( 
.A(n_5890),
.Y(n_6015)
);

INVx1_ASAP7_75t_L g6016 ( 
.A(n_5794),
.Y(n_6016)
);

AND2x2_ASAP7_75t_L g6017 ( 
.A(n_5883),
.B(n_632),
.Y(n_6017)
);

INVx2_ASAP7_75t_L g6018 ( 
.A(n_5837),
.Y(n_6018)
);

INVx2_ASAP7_75t_L g6019 ( 
.A(n_5878),
.Y(n_6019)
);

INVxp67_ASAP7_75t_SL g6020 ( 
.A(n_5940),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5796),
.Y(n_6021)
);

NAND2xp5_ASAP7_75t_L g6022 ( 
.A(n_5831),
.B(n_633),
.Y(n_6022)
);

INVx1_ASAP7_75t_SL g6023 ( 
.A(n_5844),
.Y(n_6023)
);

INVx2_ASAP7_75t_L g6024 ( 
.A(n_5878),
.Y(n_6024)
);

AOI22xp33_ASAP7_75t_SL g6025 ( 
.A1(n_5827),
.A2(n_635),
.B1(n_633),
.B2(n_634),
.Y(n_6025)
);

HB1xp67_ASAP7_75t_L g6026 ( 
.A(n_5903),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_5875),
.Y(n_6027)
);

AND2x2_ASAP7_75t_L g6028 ( 
.A(n_5789),
.B(n_5905),
.Y(n_6028)
);

AND2x2_ASAP7_75t_L g6029 ( 
.A(n_5921),
.B(n_634),
.Y(n_6029)
);

NAND2xp5_ASAP7_75t_L g6030 ( 
.A(n_5885),
.B(n_636),
.Y(n_6030)
);

AND2x2_ASAP7_75t_L g6031 ( 
.A(n_5925),
.B(n_636),
.Y(n_6031)
);

INVx2_ASAP7_75t_L g6032 ( 
.A(n_5836),
.Y(n_6032)
);

AND2x2_ASAP7_75t_L g6033 ( 
.A(n_5926),
.B(n_637),
.Y(n_6033)
);

AND2x2_ASAP7_75t_L g6034 ( 
.A(n_5931),
.B(n_637),
.Y(n_6034)
);

AND2x2_ASAP7_75t_L g6035 ( 
.A(n_5933),
.B(n_639),
.Y(n_6035)
);

AND2x2_ASAP7_75t_L g6036 ( 
.A(n_5939),
.B(n_639),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5830),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_5785),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5941),
.B(n_640),
.Y(n_6039)
);

NOR2x1_ASAP7_75t_L g6040 ( 
.A(n_5872),
.B(n_640),
.Y(n_6040)
);

AND2x2_ASAP7_75t_L g6041 ( 
.A(n_5870),
.B(n_5845),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5935),
.Y(n_6042)
);

AND2x2_ASAP7_75t_L g6043 ( 
.A(n_5826),
.B(n_641),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5805),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5806),
.Y(n_6045)
);

INVxp67_ASAP7_75t_L g6046 ( 
.A(n_5909),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5900),
.Y(n_6047)
);

OR2x2_ASAP7_75t_L g6048 ( 
.A(n_5798),
.B(n_5911),
.Y(n_6048)
);

OR2x2_ASAP7_75t_L g6049 ( 
.A(n_5787),
.B(n_1795),
.Y(n_6049)
);

AND2x2_ASAP7_75t_L g6050 ( 
.A(n_5820),
.B(n_642),
.Y(n_6050)
);

NOR2xp67_ASAP7_75t_L g6051 ( 
.A(n_5833),
.B(n_642),
.Y(n_6051)
);

INVx1_ASAP7_75t_L g6052 ( 
.A(n_5895),
.Y(n_6052)
);

NOR2xp33_ASAP7_75t_L g6053 ( 
.A(n_5843),
.B(n_643),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5862),
.B(n_644),
.Y(n_6054)
);

INVx2_ASAP7_75t_L g6055 ( 
.A(n_5886),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5901),
.Y(n_6056)
);

INVx1_ASAP7_75t_L g6057 ( 
.A(n_5908),
.Y(n_6057)
);

INVx1_ASAP7_75t_L g6058 ( 
.A(n_5910),
.Y(n_6058)
);

OR2x2_ASAP7_75t_L g6059 ( 
.A(n_5915),
.B(n_5919),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5922),
.Y(n_6060)
);

INVx1_ASAP7_75t_L g6061 ( 
.A(n_5930),
.Y(n_6061)
);

OR2x2_ASAP7_75t_L g6062 ( 
.A(n_5932),
.B(n_1797),
.Y(n_6062)
);

BUFx6f_ASAP7_75t_L g6063 ( 
.A(n_5821),
.Y(n_6063)
);

AOI22xp33_ASAP7_75t_SL g6064 ( 
.A1(n_5823),
.A2(n_647),
.B1(n_644),
.B2(n_645),
.Y(n_6064)
);

AND2x2_ASAP7_75t_L g6065 ( 
.A(n_5871),
.B(n_645),
.Y(n_6065)
);

INVx2_ASAP7_75t_L g6066 ( 
.A(n_5942),
.Y(n_6066)
);

AOI22xp33_ASAP7_75t_L g6067 ( 
.A1(n_5891),
.A2(n_649),
.B1(n_647),
.B2(n_648),
.Y(n_6067)
);

INVxp67_ASAP7_75t_SL g6068 ( 
.A(n_5835),
.Y(n_6068)
);

AND2x4_ASAP7_75t_L g6069 ( 
.A(n_5893),
.B(n_651),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5934),
.Y(n_6070)
);

INVx2_ASAP7_75t_L g6071 ( 
.A(n_5936),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_5784),
.B(n_651),
.Y(n_6072)
);

INVx2_ASAP7_75t_L g6073 ( 
.A(n_5945),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5853),
.Y(n_6074)
);

INVxp67_ASAP7_75t_SL g6075 ( 
.A(n_5788),
.Y(n_6075)
);

INVxp67_ASAP7_75t_L g6076 ( 
.A(n_5858),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_5880),
.B(n_652),
.Y(n_6077)
);

INVx1_ASAP7_75t_L g6078 ( 
.A(n_5855),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_5792),
.Y(n_6079)
);

AOI22xp33_ASAP7_75t_L g6080 ( 
.A1(n_5861),
.A2(n_655),
.B1(n_653),
.B2(n_654),
.Y(n_6080)
);

NOR2xp67_ASAP7_75t_L g6081 ( 
.A(n_5873),
.B(n_653),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_5797),
.Y(n_6082)
);

NAND2xp5_ASAP7_75t_L g6083 ( 
.A(n_5884),
.B(n_656),
.Y(n_6083)
);

INVx2_ASAP7_75t_L g6084 ( 
.A(n_5800),
.Y(n_6084)
);

INVx1_ASAP7_75t_L g6085 ( 
.A(n_5802),
.Y(n_6085)
);

INVx1_ASAP7_75t_L g6086 ( 
.A(n_5804),
.Y(n_6086)
);

INVx1_ASAP7_75t_L g6087 ( 
.A(n_5807),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5808),
.Y(n_6088)
);

INVxp67_ASAP7_75t_SL g6089 ( 
.A(n_5923),
.Y(n_6089)
);

AOI22xp33_ASAP7_75t_L g6090 ( 
.A1(n_5829),
.A2(n_5864),
.B1(n_5888),
.B2(n_5879),
.Y(n_6090)
);

AND2x2_ASAP7_75t_L g6091 ( 
.A(n_5852),
.B(n_656),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5854),
.Y(n_6092)
);

INVx1_ASAP7_75t_L g6093 ( 
.A(n_5881),
.Y(n_6093)
);

INVx2_ASAP7_75t_L g6094 ( 
.A(n_5887),
.Y(n_6094)
);

INVx2_ASAP7_75t_L g6095 ( 
.A(n_5894),
.Y(n_6095)
);

NOR2x1_ASAP7_75t_L g6096 ( 
.A(n_5897),
.B(n_657),
.Y(n_6096)
);

INVx1_ASAP7_75t_SL g6097 ( 
.A(n_5860),
.Y(n_6097)
);

AND2x4_ASAP7_75t_L g6098 ( 
.A(n_5869),
.B(n_657),
.Y(n_6098)
);

HB1xp67_ASAP7_75t_L g6099 ( 
.A(n_5889),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_5929),
.B(n_658),
.Y(n_6100)
);

INVx3_ASAP7_75t_L g6101 ( 
.A(n_5795),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_5786),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_5795),
.B(n_658),
.Y(n_6103)
);

AND2x2_ASAP7_75t_L g6104 ( 
.A(n_5795),
.B(n_659),
.Y(n_6104)
);

OAI21xp33_ASAP7_75t_L g6105 ( 
.A1(n_5829),
.A2(n_659),
.B(n_660),
.Y(n_6105)
);

NAND2xp5_ASAP7_75t_L g6106 ( 
.A(n_5907),
.B(n_660),
.Y(n_6106)
);

INVx1_ASAP7_75t_L g6107 ( 
.A(n_5786),
.Y(n_6107)
);

AND2x2_ASAP7_75t_L g6108 ( 
.A(n_5795),
.B(n_661),
.Y(n_6108)
);

AND2x4_ASAP7_75t_L g6109 ( 
.A(n_5795),
.B(n_661),
.Y(n_6109)
);

NOR2x1_ASAP7_75t_L g6110 ( 
.A(n_5810),
.B(n_662),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5786),
.Y(n_6111)
);

BUFx12f_ASAP7_75t_L g6112 ( 
.A(n_5927),
.Y(n_6112)
);

OR2x2_ASAP7_75t_L g6113 ( 
.A(n_5840),
.B(n_1797),
.Y(n_6113)
);

INVxp67_ASAP7_75t_L g6114 ( 
.A(n_5890),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_5786),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_5786),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5786),
.Y(n_6117)
);

AND2x2_ASAP7_75t_L g6118 ( 
.A(n_5795),
.B(n_662),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5786),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_5786),
.Y(n_6120)
);

HB1xp67_ASAP7_75t_L g6121 ( 
.A(n_5803),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5786),
.Y(n_6122)
);

INVx2_ASAP7_75t_SL g6123 ( 
.A(n_5795),
.Y(n_6123)
);

OAI22xp5_ASAP7_75t_SL g6124 ( 
.A1(n_5793),
.A2(n_665),
.B1(n_663),
.B2(n_664),
.Y(n_6124)
);

NOR2x1_ASAP7_75t_L g6125 ( 
.A(n_5810),
.B(n_664),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5786),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_5786),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5786),
.Y(n_6128)
);

AND2x2_ASAP7_75t_L g6129 ( 
.A(n_5795),
.B(n_665),
.Y(n_6129)
);

INVx1_ASAP7_75t_L g6130 ( 
.A(n_5786),
.Y(n_6130)
);

INVx1_ASAP7_75t_L g6131 ( 
.A(n_5786),
.Y(n_6131)
);

AOI21xp33_ASAP7_75t_L g6132 ( 
.A1(n_5793),
.A2(n_666),
.B(n_667),
.Y(n_6132)
);

INVx1_ASAP7_75t_L g6133 ( 
.A(n_5786),
.Y(n_6133)
);

BUFx2_ASAP7_75t_L g6134 ( 
.A(n_5795),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_5795),
.B(n_667),
.Y(n_6135)
);

NAND2xp5_ASAP7_75t_L g6136 ( 
.A(n_5907),
.B(n_668),
.Y(n_6136)
);

INVx1_ASAP7_75t_L g6137 ( 
.A(n_5786),
.Y(n_6137)
);

INVx2_ASAP7_75t_L g6138 ( 
.A(n_5795),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_5786),
.Y(n_6139)
);

AND2x2_ASAP7_75t_L g6140 ( 
.A(n_5795),
.B(n_668),
.Y(n_6140)
);

OAI22xp5_ASAP7_75t_L g6141 ( 
.A1(n_5793),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.Y(n_6141)
);

AOI22xp33_ASAP7_75t_L g6142 ( 
.A1(n_5892),
.A2(n_671),
.B1(n_669),
.B2(n_670),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5786),
.Y(n_6143)
);

NAND2xp5_ASAP7_75t_L g6144 ( 
.A(n_5907),
.B(n_672),
.Y(n_6144)
);

INVx1_ASAP7_75t_L g6145 ( 
.A(n_5786),
.Y(n_6145)
);

INVx2_ASAP7_75t_SL g6146 ( 
.A(n_5795),
.Y(n_6146)
);

OAI22xp5_ASAP7_75t_L g6147 ( 
.A1(n_6068),
.A2(n_675),
.B1(n_672),
.B2(n_673),
.Y(n_6147)
);

AND2x2_ASAP7_75t_L g6148 ( 
.A(n_5985),
.B(n_673),
.Y(n_6148)
);

INVx2_ASAP7_75t_L g6149 ( 
.A(n_5949),
.Y(n_6149)
);

NAND3xp33_ASAP7_75t_L g6150 ( 
.A(n_5967),
.B(n_675),
.C(n_676),
.Y(n_6150)
);

AND2x2_ASAP7_75t_L g6151 ( 
.A(n_5952),
.B(n_677),
.Y(n_6151)
);

INVx1_ASAP7_75t_L g6152 ( 
.A(n_5999),
.Y(n_6152)
);

CKINVDCx20_ASAP7_75t_R g6153 ( 
.A(n_5953),
.Y(n_6153)
);

BUFx3_ASAP7_75t_L g6154 ( 
.A(n_6112),
.Y(n_6154)
);

AND2x2_ASAP7_75t_SL g6155 ( 
.A(n_6134),
.B(n_677),
.Y(n_6155)
);

INVx3_ASAP7_75t_L g6156 ( 
.A(n_5983),
.Y(n_6156)
);

OAI33xp33_ASAP7_75t_L g6157 ( 
.A1(n_6124),
.A2(n_680),
.A3(n_682),
.B1(n_678),
.B2(n_679),
.B3(n_681),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_6027),
.Y(n_6158)
);

NOR2xp33_ASAP7_75t_L g6159 ( 
.A(n_5975),
.B(n_678),
.Y(n_6159)
);

INVx2_ASAP7_75t_L g6160 ( 
.A(n_5994),
.Y(n_6160)
);

AOI22xp33_ASAP7_75t_L g6161 ( 
.A1(n_6005),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_6161)
);

INVx2_ASAP7_75t_L g6162 ( 
.A(n_6028),
.Y(n_6162)
);

OAI31xp33_ASAP7_75t_L g6163 ( 
.A1(n_5955),
.A2(n_684),
.A3(n_682),
.B(n_683),
.Y(n_6163)
);

NAND2xp5_ASAP7_75t_L g6164 ( 
.A(n_6065),
.B(n_683),
.Y(n_6164)
);

INVx2_ASAP7_75t_L g6165 ( 
.A(n_5948),
.Y(n_6165)
);

AOI22xp33_ASAP7_75t_L g6166 ( 
.A1(n_6020),
.A2(n_687),
.B1(n_685),
.B2(n_686),
.Y(n_6166)
);

INVx1_ASAP7_75t_L g6167 ( 
.A(n_5951),
.Y(n_6167)
);

BUFx3_ASAP7_75t_L g6168 ( 
.A(n_5975),
.Y(n_6168)
);

NAND3xp33_ASAP7_75t_L g6169 ( 
.A(n_6141),
.B(n_685),
.C(n_688),
.Y(n_6169)
);

INVx1_ASAP7_75t_L g6170 ( 
.A(n_5958),
.Y(n_6170)
);

OAI211xp5_ASAP7_75t_SL g6171 ( 
.A1(n_5950),
.A2(n_691),
.B(n_689),
.C(n_690),
.Y(n_6171)
);

AND2x2_ASAP7_75t_L g6172 ( 
.A(n_6101),
.B(n_689),
.Y(n_6172)
);

INVx2_ASAP7_75t_L g6173 ( 
.A(n_6138),
.Y(n_6173)
);

NAND4xp25_ASAP7_75t_SL g6174 ( 
.A(n_5959),
.B(n_692),
.C(n_690),
.D(n_691),
.Y(n_6174)
);

CKINVDCx14_ASAP7_75t_R g6175 ( 
.A(n_5975),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_6123),
.Y(n_6176)
);

OAI33xp33_ASAP7_75t_L g6177 ( 
.A1(n_6008),
.A2(n_694),
.A3(n_696),
.B1(n_692),
.B2(n_693),
.B3(n_695),
.Y(n_6177)
);

INVx2_ASAP7_75t_L g6178 ( 
.A(n_6146),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_6063),
.Y(n_6179)
);

NOR3xp33_ASAP7_75t_L g6180 ( 
.A(n_6023),
.B(n_694),
.C(n_695),
.Y(n_6180)
);

AND2x4_ASAP7_75t_L g6181 ( 
.A(n_5982),
.B(n_696),
.Y(n_6181)
);

AOI211xp5_ASAP7_75t_L g6182 ( 
.A1(n_6132),
.A2(n_699),
.B(n_700),
.C(n_698),
.Y(n_6182)
);

OR2x6_ASAP7_75t_L g6183 ( 
.A(n_6063),
.B(n_697),
.Y(n_6183)
);

NAND2xp5_ASAP7_75t_L g6184 ( 
.A(n_6000),
.B(n_698),
.Y(n_6184)
);

NAND2xp5_ASAP7_75t_L g6185 ( 
.A(n_6074),
.B(n_699),
.Y(n_6185)
);

AND2x2_ASAP7_75t_L g6186 ( 
.A(n_5987),
.B(n_700),
.Y(n_6186)
);

INVx4_ASAP7_75t_L g6187 ( 
.A(n_6004),
.Y(n_6187)
);

NAND2xp5_ASAP7_75t_L g6188 ( 
.A(n_5989),
.B(n_701),
.Y(n_6188)
);

AND2x2_ASAP7_75t_L g6189 ( 
.A(n_6097),
.B(n_702),
.Y(n_6189)
);

INVx2_ASAP7_75t_SL g6190 ( 
.A(n_6010),
.Y(n_6190)
);

OAI22xp5_ASAP7_75t_L g6191 ( 
.A1(n_6121),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_6191)
);

AOI21xp5_ASAP7_75t_L g6192 ( 
.A1(n_6110),
.A2(n_704),
.B(n_705),
.Y(n_6192)
);

NOR4xp25_ASAP7_75t_SL g6193 ( 
.A(n_6014),
.B(n_707),
.C(n_705),
.D(n_706),
.Y(n_6193)
);

AOI22xp33_ASAP7_75t_L g6194 ( 
.A1(n_6066),
.A2(n_710),
.B1(n_706),
.B2(n_708),
.Y(n_6194)
);

OR2x2_ASAP7_75t_L g6195 ( 
.A(n_5957),
.B(n_6078),
.Y(n_6195)
);

INVx2_ASAP7_75t_L g6196 ( 
.A(n_6019),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_5970),
.Y(n_6197)
);

OAI21xp33_ASAP7_75t_SL g6198 ( 
.A1(n_6125),
.A2(n_708),
.B(n_711),
.Y(n_6198)
);

AND2x2_ASAP7_75t_L g6199 ( 
.A(n_6012),
.B(n_712),
.Y(n_6199)
);

OR2x2_ASAP7_75t_L g6200 ( 
.A(n_6044),
.B(n_712),
.Y(n_6200)
);

OAI31xp33_ASAP7_75t_L g6201 ( 
.A1(n_6026),
.A2(n_715),
.A3(n_713),
.B(n_714),
.Y(n_6201)
);

CKINVDCx5p33_ASAP7_75t_R g6202 ( 
.A(n_5954),
.Y(n_6202)
);

NAND2xp33_ASAP7_75t_R g6203 ( 
.A(n_5968),
.B(n_713),
.Y(n_6203)
);

INVxp67_ASAP7_75t_L g6204 ( 
.A(n_6081),
.Y(n_6204)
);

AOI222xp33_ASAP7_75t_L g6205 ( 
.A1(n_5964),
.A2(n_717),
.B1(n_719),
.B2(n_715),
.C1(n_716),
.C2(n_718),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5971),
.Y(n_6206)
);

OAI221xp5_ASAP7_75t_L g6207 ( 
.A1(n_5997),
.A2(n_720),
.B1(n_716),
.B2(n_719),
.C(n_721),
.Y(n_6207)
);

OAI21xp5_ASAP7_75t_SL g6208 ( 
.A1(n_5981),
.A2(n_720),
.B(n_721),
.Y(n_6208)
);

A2O1A1Ixp33_ASAP7_75t_L g6209 ( 
.A1(n_6018),
.A2(n_730),
.B(n_739),
.C(n_722),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_5976),
.Y(n_6210)
);

INVx2_ASAP7_75t_L g6211 ( 
.A(n_6024),
.Y(n_6211)
);

INVx2_ASAP7_75t_SL g6212 ( 
.A(n_5947),
.Y(n_6212)
);

AND2x2_ASAP7_75t_SL g6213 ( 
.A(n_6032),
.B(n_722),
.Y(n_6213)
);

NAND2xp5_ASAP7_75t_L g6214 ( 
.A(n_6099),
.B(n_723),
.Y(n_6214)
);

AOI21x1_ASAP7_75t_L g6215 ( 
.A1(n_6051),
.A2(n_723),
.B(n_724),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_5966),
.B(n_724),
.Y(n_6216)
);

OAI221xp5_ASAP7_75t_SL g6217 ( 
.A1(n_6089),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.C(n_728),
.Y(n_6217)
);

NOR2xp33_ASAP7_75t_L g6218 ( 
.A(n_6015),
.B(n_725),
.Y(n_6218)
);

OAI221xp5_ASAP7_75t_L g6219 ( 
.A1(n_5962),
.A2(n_728),
.B1(n_726),
.B2(n_727),
.C(n_729),
.Y(n_6219)
);

AOI22xp33_ASAP7_75t_L g6220 ( 
.A1(n_6046),
.A2(n_732),
.B1(n_729),
.B2(n_731),
.Y(n_6220)
);

OR2x6_ASAP7_75t_L g6221 ( 
.A(n_5956),
.B(n_732),
.Y(n_6221)
);

HB1xp67_ASAP7_75t_L g6222 ( 
.A(n_6114),
.Y(n_6222)
);

OR2x2_ASAP7_75t_L g6223 ( 
.A(n_6045),
.B(n_733),
.Y(n_6223)
);

INVx1_ASAP7_75t_L g6224 ( 
.A(n_5977),
.Y(n_6224)
);

NAND2xp5_ASAP7_75t_L g6225 ( 
.A(n_6047),
.B(n_733),
.Y(n_6225)
);

NAND2xp5_ASAP7_75t_L g6226 ( 
.A(n_5974),
.B(n_734),
.Y(n_6226)
);

NOR2xp33_ASAP7_75t_L g6227 ( 
.A(n_6048),
.B(n_736),
.Y(n_6227)
);

BUFx2_ASAP7_75t_L g6228 ( 
.A(n_6095),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_5979),
.Y(n_6229)
);

INVx2_ASAP7_75t_L g6230 ( 
.A(n_6094),
.Y(n_6230)
);

AND2x2_ASAP7_75t_L g6231 ( 
.A(n_5961),
.B(n_736),
.Y(n_6231)
);

AOI221xp5_ASAP7_75t_L g6232 ( 
.A1(n_6075),
.A2(n_739),
.B1(n_737),
.B2(n_738),
.C(n_740),
.Y(n_6232)
);

OAI211xp5_ASAP7_75t_SL g6233 ( 
.A1(n_6090),
.A2(n_742),
.B(n_738),
.C(n_741),
.Y(n_6233)
);

HB1xp67_ASAP7_75t_L g6234 ( 
.A(n_6037),
.Y(n_6234)
);

BUFx3_ASAP7_75t_L g6235 ( 
.A(n_6043),
.Y(n_6235)
);

NOR4xp25_ASAP7_75t_SL g6236 ( 
.A(n_6093),
.B(n_743),
.C(n_741),
.D(n_742),
.Y(n_6236)
);

AO21x2_ASAP7_75t_L g6237 ( 
.A1(n_6022),
.A2(n_743),
.B(n_744),
.Y(n_6237)
);

INVx1_ASAP7_75t_L g6238 ( 
.A(n_5980),
.Y(n_6238)
);

AND2x2_ASAP7_75t_L g6239 ( 
.A(n_6041),
.B(n_744),
.Y(n_6239)
);

OAI33xp33_ASAP7_75t_L g6240 ( 
.A1(n_5998),
.A2(n_747),
.A3(n_749),
.B1(n_745),
.B2(n_746),
.B3(n_748),
.Y(n_6240)
);

INVx3_ASAP7_75t_L g6241 ( 
.A(n_6109),
.Y(n_6241)
);

OAI211xp5_ASAP7_75t_L g6242 ( 
.A1(n_6105),
.A2(n_750),
.B(n_747),
.C(n_748),
.Y(n_6242)
);

OAI321xp33_ASAP7_75t_L g6243 ( 
.A1(n_6080),
.A2(n_752),
.A3(n_754),
.B1(n_750),
.B2(n_751),
.C(n_753),
.Y(n_6243)
);

AOI22xp33_ASAP7_75t_L g6244 ( 
.A1(n_6055),
.A2(n_753),
.B1(n_751),
.B2(n_752),
.Y(n_6244)
);

OAI31xp33_ASAP7_75t_L g6245 ( 
.A1(n_5960),
.A2(n_757),
.A3(n_755),
.B(n_756),
.Y(n_6245)
);

OA21x2_ASAP7_75t_L g6246 ( 
.A1(n_6076),
.A2(n_755),
.B(n_756),
.Y(n_6246)
);

HB1xp67_ASAP7_75t_L g6247 ( 
.A(n_6038),
.Y(n_6247)
);

NAND2xp33_ASAP7_75t_SL g6248 ( 
.A(n_6103),
.B(n_758),
.Y(n_6248)
);

AOI22xp33_ASAP7_75t_L g6249 ( 
.A1(n_6052),
.A2(n_760),
.B1(n_758),
.B2(n_759),
.Y(n_6249)
);

NAND4xp25_ASAP7_75t_L g6250 ( 
.A(n_5991),
.B(n_762),
.C(n_760),
.D(n_761),
.Y(n_6250)
);

AOI31xp33_ASAP7_75t_L g6251 ( 
.A1(n_6096),
.A2(n_765),
.A3(n_763),
.B(n_764),
.Y(n_6251)
);

AOI22xp33_ASAP7_75t_L g6252 ( 
.A1(n_6056),
.A2(n_766),
.B1(n_763),
.B2(n_765),
.Y(n_6252)
);

HB1xp67_ASAP7_75t_L g6253 ( 
.A(n_6042),
.Y(n_6253)
);

BUFx2_ASAP7_75t_L g6254 ( 
.A(n_5965),
.Y(n_6254)
);

AOI22xp33_ASAP7_75t_L g6255 ( 
.A1(n_6057),
.A2(n_769),
.B1(n_767),
.B2(n_768),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_5984),
.Y(n_6256)
);

INVx2_ASAP7_75t_SL g6257 ( 
.A(n_6104),
.Y(n_6257)
);

AOI21xp5_ASAP7_75t_L g6258 ( 
.A1(n_5986),
.A2(n_768),
.B(n_770),
.Y(n_6258)
);

OAI22xp33_ASAP7_75t_L g6259 ( 
.A1(n_5963),
.A2(n_773),
.B1(n_771),
.B2(n_772),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_5990),
.Y(n_6260)
);

NAND3xp33_ASAP7_75t_L g6261 ( 
.A(n_6064),
.B(n_771),
.C(n_772),
.Y(n_6261)
);

AOI221xp5_ASAP7_75t_L g6262 ( 
.A1(n_6106),
.A2(n_776),
.B1(n_774),
.B2(n_775),
.C(n_777),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_6102),
.Y(n_6263)
);

OAI33xp33_ASAP7_75t_L g6264 ( 
.A1(n_6001),
.A2(n_777),
.A3(n_780),
.B1(n_775),
.B2(n_776),
.B3(n_779),
.Y(n_6264)
);

NAND2xp5_ASAP7_75t_L g6265 ( 
.A(n_5993),
.B(n_780),
.Y(n_6265)
);

NAND4xp25_ASAP7_75t_L g6266 ( 
.A(n_5995),
.B(n_783),
.C(n_781),
.D(n_782),
.Y(n_6266)
);

NAND2xp5_ASAP7_75t_L g6267 ( 
.A(n_6009),
.B(n_783),
.Y(n_6267)
);

AND2x2_ASAP7_75t_L g6268 ( 
.A(n_6108),
.B(n_784),
.Y(n_6268)
);

INVx2_ASAP7_75t_L g6269 ( 
.A(n_6049),
.Y(n_6269)
);

AND2x2_ASAP7_75t_L g6270 ( 
.A(n_6118),
.B(n_784),
.Y(n_6270)
);

OR2x2_ASAP7_75t_L g6271 ( 
.A(n_5978),
.B(n_785),
.Y(n_6271)
);

AOI21xp5_ASAP7_75t_L g6272 ( 
.A1(n_6136),
.A2(n_785),
.B(n_786),
.Y(n_6272)
);

NAND2xp33_ASAP7_75t_R g6273 ( 
.A(n_6144),
.B(n_787),
.Y(n_6273)
);

NOR2x1_ASAP7_75t_L g6274 ( 
.A(n_5946),
.B(n_787),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_6129),
.B(n_788),
.Y(n_6275)
);

AOI221xp5_ASAP7_75t_L g6276 ( 
.A1(n_6072),
.A2(n_5972),
.B1(n_6083),
.B2(n_6002),
.C(n_6021),
.Y(n_6276)
);

INVx1_ASAP7_75t_SL g6277 ( 
.A(n_6050),
.Y(n_6277)
);

AND2x2_ASAP7_75t_L g6278 ( 
.A(n_6135),
.B(n_789),
.Y(n_6278)
);

AND2x2_ASAP7_75t_L g6279 ( 
.A(n_6140),
.B(n_5992),
.Y(n_6279)
);

AOI221xp5_ASAP7_75t_L g6280 ( 
.A1(n_6016),
.A2(n_791),
.B1(n_789),
.B2(n_790),
.C(n_792),
.Y(n_6280)
);

AOI22xp5_ASAP7_75t_L g6281 ( 
.A1(n_6040),
.A2(n_6100),
.B1(n_6017),
.B2(n_6092),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_6107),
.Y(n_6282)
);

AOI221xp5_ASAP7_75t_L g6283 ( 
.A1(n_6003),
.A2(n_792),
.B1(n_790),
.B2(n_791),
.C(n_793),
.Y(n_6283)
);

INVx1_ASAP7_75t_L g6284 ( 
.A(n_6111),
.Y(n_6284)
);

INVx1_ASAP7_75t_L g6285 ( 
.A(n_6115),
.Y(n_6285)
);

OAI22xp5_ASAP7_75t_L g6286 ( 
.A1(n_6030),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_6286)
);

BUFx2_ASAP7_75t_L g6287 ( 
.A(n_6007),
.Y(n_6287)
);

INVx1_ASAP7_75t_L g6288 ( 
.A(n_6116),
.Y(n_6288)
);

AOI22xp5_ASAP7_75t_L g6289 ( 
.A1(n_6062),
.A2(n_797),
.B1(n_795),
.B2(n_796),
.Y(n_6289)
);

INVx2_ASAP7_75t_SL g6290 ( 
.A(n_6054),
.Y(n_6290)
);

AOI22xp33_ASAP7_75t_L g6291 ( 
.A1(n_6058),
.A2(n_799),
.B1(n_797),
.B2(n_798),
.Y(n_6291)
);

OAI21x1_ASAP7_75t_L g6292 ( 
.A1(n_6070),
.A2(n_799),
.B(n_800),
.Y(n_6292)
);

INVxp67_ASAP7_75t_SL g6293 ( 
.A(n_6006),
.Y(n_6293)
);

AND2x2_ASAP7_75t_L g6294 ( 
.A(n_6175),
.B(n_5996),
.Y(n_6294)
);

AND2x2_ASAP7_75t_L g6295 ( 
.A(n_6156),
.B(n_6117),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_6222),
.Y(n_6296)
);

BUFx2_ASAP7_75t_SL g6297 ( 
.A(n_6153),
.Y(n_6297)
);

INVx2_ASAP7_75t_L g6298 ( 
.A(n_6235),
.Y(n_6298)
);

INVx1_ASAP7_75t_L g6299 ( 
.A(n_6189),
.Y(n_6299)
);

NAND2xp5_ASAP7_75t_L g6300 ( 
.A(n_6277),
.B(n_6113),
.Y(n_6300)
);

AND2x4_ASAP7_75t_L g6301 ( 
.A(n_6168),
.B(n_6013),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_6184),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_6187),
.B(n_6119),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_6228),
.Y(n_6304)
);

OR2x2_ASAP7_75t_L g6305 ( 
.A(n_6254),
.B(n_6195),
.Y(n_6305)
);

HB1xp67_ASAP7_75t_L g6306 ( 
.A(n_6149),
.Y(n_6306)
);

AND2x2_ASAP7_75t_L g6307 ( 
.A(n_6190),
.B(n_6120),
.Y(n_6307)
);

INVx2_ASAP7_75t_L g6308 ( 
.A(n_6279),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_6183),
.Y(n_6309)
);

OR2x2_ASAP7_75t_L g6310 ( 
.A(n_6214),
.B(n_6152),
.Y(n_6310)
);

AND2x4_ASAP7_75t_L g6311 ( 
.A(n_6290),
.B(n_5973),
.Y(n_6311)
);

NAND2xp5_ASAP7_75t_SL g6312 ( 
.A(n_6212),
.B(n_6011),
.Y(n_6312)
);

AND2x2_ASAP7_75t_L g6313 ( 
.A(n_6162),
.B(n_6122),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_6188),
.Y(n_6314)
);

AND2x2_ASAP7_75t_L g6315 ( 
.A(n_6241),
.B(n_6126),
.Y(n_6315)
);

INVx1_ASAP7_75t_L g6316 ( 
.A(n_6200),
.Y(n_6316)
);

BUFx2_ASAP7_75t_SL g6317 ( 
.A(n_6154),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6223),
.Y(n_6318)
);

OR2x2_ASAP7_75t_L g6319 ( 
.A(n_6287),
.B(n_6127),
.Y(n_6319)
);

AND2x2_ASAP7_75t_L g6320 ( 
.A(n_6176),
.B(n_6178),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_6247),
.Y(n_6321)
);

INVx1_ASAP7_75t_L g6322 ( 
.A(n_6253),
.Y(n_6322)
);

INVx2_ASAP7_75t_L g6323 ( 
.A(n_6183),
.Y(n_6323)
);

INVx1_ASAP7_75t_SL g6324 ( 
.A(n_6155),
.Y(n_6324)
);

NOR2x1_ASAP7_75t_L g6325 ( 
.A(n_6150),
.B(n_6091),
.Y(n_6325)
);

OR2x2_ASAP7_75t_L g6326 ( 
.A(n_6226),
.B(n_6128),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_6148),
.Y(n_6327)
);

NAND2x1p5_ASAP7_75t_L g6328 ( 
.A(n_6172),
.B(n_6181),
.Y(n_6328)
);

HB1xp67_ASAP7_75t_L g6329 ( 
.A(n_6179),
.Y(n_6329)
);

OR2x2_ASAP7_75t_L g6330 ( 
.A(n_6185),
.B(n_6130),
.Y(n_6330)
);

INVx1_ASAP7_75t_L g6331 ( 
.A(n_6225),
.Y(n_6331)
);

AND2x2_ASAP7_75t_L g6332 ( 
.A(n_6151),
.B(n_6202),
.Y(n_6332)
);

AND2x4_ASAP7_75t_L g6333 ( 
.A(n_6257),
.B(n_6160),
.Y(n_6333)
);

HB1xp67_ASAP7_75t_L g6334 ( 
.A(n_6165),
.Y(n_6334)
);

NAND2xp5_ASAP7_75t_L g6335 ( 
.A(n_6293),
.B(n_6029),
.Y(n_6335)
);

OR2x2_ASAP7_75t_L g6336 ( 
.A(n_6173),
.B(n_6196),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_6167),
.Y(n_6337)
);

INVxp33_ASAP7_75t_SL g6338 ( 
.A(n_6216),
.Y(n_6338)
);

AND2x2_ASAP7_75t_L g6339 ( 
.A(n_6186),
.B(n_6131),
.Y(n_6339)
);

INVx1_ASAP7_75t_L g6340 ( 
.A(n_6170),
.Y(n_6340)
);

AND2x2_ASAP7_75t_L g6341 ( 
.A(n_6199),
.B(n_6133),
.Y(n_6341)
);

NAND2xp5_ASAP7_75t_L g6342 ( 
.A(n_6180),
.B(n_6031),
.Y(n_6342)
);

AND2x2_ASAP7_75t_L g6343 ( 
.A(n_6218),
.B(n_6137),
.Y(n_6343)
);

NAND2xp5_ASAP7_75t_L g6344 ( 
.A(n_6227),
.B(n_6033),
.Y(n_6344)
);

INVx1_ASAP7_75t_L g6345 ( 
.A(n_6197),
.Y(n_6345)
);

AND2x4_ASAP7_75t_L g6346 ( 
.A(n_6239),
.B(n_6069),
.Y(n_6346)
);

HB1xp67_ASAP7_75t_L g6347 ( 
.A(n_6211),
.Y(n_6347)
);

NOR2xp33_ASAP7_75t_L g6348 ( 
.A(n_6251),
.B(n_5969),
.Y(n_6348)
);

INVxp67_ASAP7_75t_SL g6349 ( 
.A(n_6203),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_6206),
.Y(n_6350)
);

AND2x2_ASAP7_75t_L g6351 ( 
.A(n_6159),
.B(n_6231),
.Y(n_6351)
);

INVx1_ASAP7_75t_L g6352 ( 
.A(n_6210),
.Y(n_6352)
);

INVx1_ASAP7_75t_L g6353 ( 
.A(n_6224),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_6158),
.B(n_6139),
.Y(n_6354)
);

INVx2_ASAP7_75t_L g6355 ( 
.A(n_6215),
.Y(n_6355)
);

INVx2_ASAP7_75t_L g6356 ( 
.A(n_6221),
.Y(n_6356)
);

NOR2x1_ASAP7_75t_L g6357 ( 
.A(n_6147),
.B(n_6034),
.Y(n_6357)
);

AND2x4_ASAP7_75t_L g6358 ( 
.A(n_6268),
.B(n_5988),
.Y(n_6358)
);

INVx1_ASAP7_75t_L g6359 ( 
.A(n_6229),
.Y(n_6359)
);

AND2x2_ASAP7_75t_L g6360 ( 
.A(n_6270),
.B(n_6143),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_6238),
.Y(n_6361)
);

INVxp67_ASAP7_75t_L g6362 ( 
.A(n_6273),
.Y(n_6362)
);

AND2x4_ASAP7_75t_L g6363 ( 
.A(n_6275),
.B(n_6035),
.Y(n_6363)
);

INVx2_ASAP7_75t_L g6364 ( 
.A(n_6221),
.Y(n_6364)
);

INVx1_ASAP7_75t_L g6365 ( 
.A(n_6256),
.Y(n_6365)
);

INVx3_ASAP7_75t_L g6366 ( 
.A(n_6278),
.Y(n_6366)
);

INVx1_ASAP7_75t_L g6367 ( 
.A(n_6260),
.Y(n_6367)
);

INVx2_ASAP7_75t_L g6368 ( 
.A(n_6213),
.Y(n_6368)
);

NAND2xp5_ASAP7_75t_L g6369 ( 
.A(n_6258),
.B(n_6036),
.Y(n_6369)
);

INVx1_ASAP7_75t_L g6370 ( 
.A(n_6263),
.Y(n_6370)
);

AND2x2_ASAP7_75t_L g6371 ( 
.A(n_6282),
.B(n_6145),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_6284),
.Y(n_6372)
);

NAND2xp5_ASAP7_75t_L g6373 ( 
.A(n_6272),
.B(n_6205),
.Y(n_6373)
);

HB1xp67_ASAP7_75t_L g6374 ( 
.A(n_6246),
.Y(n_6374)
);

INVx1_ASAP7_75t_L g6375 ( 
.A(n_6285),
.Y(n_6375)
);

AND2x2_ASAP7_75t_L g6376 ( 
.A(n_6288),
.B(n_6039),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_6234),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_6230),
.Y(n_6378)
);

OAI33xp33_ASAP7_75t_L g6379 ( 
.A1(n_6191),
.A2(n_6286),
.A3(n_6259),
.B1(n_6250),
.B2(n_6266),
.B3(n_6171),
.Y(n_6379)
);

INVx2_ASAP7_75t_L g6380 ( 
.A(n_6271),
.Y(n_6380)
);

NAND2xp5_ASAP7_75t_L g6381 ( 
.A(n_6161),
.B(n_6077),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6164),
.Y(n_6382)
);

HB1xp67_ASAP7_75t_L g6383 ( 
.A(n_6246),
.Y(n_6383)
);

INVxp67_ASAP7_75t_SL g6384 ( 
.A(n_6274),
.Y(n_6384)
);

INVx2_ASAP7_75t_L g6385 ( 
.A(n_6237),
.Y(n_6385)
);

AND2x2_ASAP7_75t_L g6386 ( 
.A(n_6276),
.B(n_6053),
.Y(n_6386)
);

NAND2xp5_ASAP7_75t_L g6387 ( 
.A(n_6166),
.B(n_6025),
.Y(n_6387)
);

OR2x2_ASAP7_75t_SL g6388 ( 
.A(n_6169),
.B(n_6059),
.Y(n_6388)
);

INVx2_ASAP7_75t_L g6389 ( 
.A(n_6204),
.Y(n_6389)
);

NAND2xp5_ASAP7_75t_L g6390 ( 
.A(n_6245),
.B(n_6142),
.Y(n_6390)
);

INVx1_ASAP7_75t_L g6391 ( 
.A(n_6265),
.Y(n_6391)
);

INVx1_ASAP7_75t_L g6392 ( 
.A(n_6267),
.Y(n_6392)
);

BUFx2_ASAP7_75t_L g6393 ( 
.A(n_6198),
.Y(n_6393)
);

NAND2xp5_ASAP7_75t_L g6394 ( 
.A(n_6362),
.B(n_6208),
.Y(n_6394)
);

AND2x2_ASAP7_75t_L g6395 ( 
.A(n_6297),
.B(n_6281),
.Y(n_6395)
);

INVx1_ASAP7_75t_L g6396 ( 
.A(n_6374),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_6383),
.Y(n_6397)
);

OR2x2_ASAP7_75t_L g6398 ( 
.A(n_6305),
.B(n_6209),
.Y(n_6398)
);

AND2x2_ASAP7_75t_L g6399 ( 
.A(n_6317),
.B(n_6232),
.Y(n_6399)
);

AND2x4_ASAP7_75t_L g6400 ( 
.A(n_6346),
.B(n_6098),
.Y(n_6400)
);

INVx2_ASAP7_75t_L g6401 ( 
.A(n_6363),
.Y(n_6401)
);

OR2x2_ASAP7_75t_L g6402 ( 
.A(n_6304),
.B(n_6201),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_6328),
.Y(n_6403)
);

AND2x2_ASAP7_75t_L g6404 ( 
.A(n_6332),
.B(n_6194),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_L g6405 ( 
.A(n_6338),
.B(n_6192),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6335),
.Y(n_6406)
);

AND2x2_ASAP7_75t_L g6407 ( 
.A(n_6301),
.B(n_6269),
.Y(n_6407)
);

AND2x2_ASAP7_75t_L g6408 ( 
.A(n_6376),
.B(n_6289),
.Y(n_6408)
);

AND2x2_ASAP7_75t_L g6409 ( 
.A(n_6339),
.B(n_6283),
.Y(n_6409)
);

NOR2xp33_ASAP7_75t_L g6410 ( 
.A(n_6379),
.B(n_6177),
.Y(n_6410)
);

NOR2xp33_ASAP7_75t_L g6411 ( 
.A(n_6324),
.B(n_6174),
.Y(n_6411)
);

INVx2_ASAP7_75t_L g6412 ( 
.A(n_6358),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_6306),
.Y(n_6413)
);

AND2x2_ASAP7_75t_L g6414 ( 
.A(n_6308),
.B(n_6163),
.Y(n_6414)
);

AND2x2_ASAP7_75t_L g6415 ( 
.A(n_6341),
.B(n_6193),
.Y(n_6415)
);

HB1xp67_ASAP7_75t_L g6416 ( 
.A(n_6329),
.Y(n_6416)
);

OR2x2_ASAP7_75t_L g6417 ( 
.A(n_6319),
.B(n_6217),
.Y(n_6417)
);

AND2x2_ASAP7_75t_L g6418 ( 
.A(n_6298),
.B(n_6236),
.Y(n_6418)
);

OR2x2_ASAP7_75t_L g6419 ( 
.A(n_6377),
.B(n_6207),
.Y(n_6419)
);

INVx4_ASAP7_75t_L g6420 ( 
.A(n_6389),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_6366),
.B(n_6262),
.Y(n_6421)
);

NOR2xp33_ASAP7_75t_L g6422 ( 
.A(n_6344),
.B(n_6240),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_6334),
.Y(n_6423)
);

INVx1_ASAP7_75t_L g6424 ( 
.A(n_6347),
.Y(n_6424)
);

HB1xp67_ASAP7_75t_L g6425 ( 
.A(n_6311),
.Y(n_6425)
);

NAND2xp5_ASAP7_75t_L g6426 ( 
.A(n_6360),
.B(n_6327),
.Y(n_6426)
);

HB1xp67_ASAP7_75t_L g6427 ( 
.A(n_6320),
.Y(n_6427)
);

AND2x2_ASAP7_75t_L g6428 ( 
.A(n_6333),
.B(n_6182),
.Y(n_6428)
);

AOI22xp5_ASAP7_75t_L g6429 ( 
.A1(n_6393),
.A2(n_6157),
.B1(n_6261),
.B2(n_6248),
.Y(n_6429)
);

AND2x2_ASAP7_75t_L g6430 ( 
.A(n_6294),
.B(n_6220),
.Y(n_6430)
);

INVx1_ASAP7_75t_L g6431 ( 
.A(n_6296),
.Y(n_6431)
);

AOI211xp5_ASAP7_75t_L g6432 ( 
.A1(n_6384),
.A2(n_6242),
.B(n_6280),
.C(n_6233),
.Y(n_6432)
);

INVxp67_ASAP7_75t_L g6433 ( 
.A(n_6349),
.Y(n_6433)
);

INVx1_ASAP7_75t_L g6434 ( 
.A(n_6310),
.Y(n_6434)
);

AND2x2_ASAP7_75t_L g6435 ( 
.A(n_6303),
.B(n_6060),
.Y(n_6435)
);

NOR2x1_ASAP7_75t_R g6436 ( 
.A(n_6312),
.B(n_6264),
.Y(n_6436)
);

HB1xp67_ASAP7_75t_L g6437 ( 
.A(n_6369),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_6351),
.Y(n_6438)
);

NAND2xp5_ASAP7_75t_L g6439 ( 
.A(n_6299),
.B(n_6244),
.Y(n_6439)
);

INVx1_ASAP7_75t_SL g6440 ( 
.A(n_6342),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6321),
.Y(n_6441)
);

INVx1_ASAP7_75t_L g6442 ( 
.A(n_6322),
.Y(n_6442)
);

AND2x2_ASAP7_75t_L g6443 ( 
.A(n_6343),
.B(n_6061),
.Y(n_6443)
);

INVx1_ASAP7_75t_L g6444 ( 
.A(n_6391),
.Y(n_6444)
);

AND2x4_ASAP7_75t_L g6445 ( 
.A(n_6307),
.B(n_6292),
.Y(n_6445)
);

AND2x2_ASAP7_75t_L g6446 ( 
.A(n_6295),
.B(n_6071),
.Y(n_6446)
);

AND2x2_ASAP7_75t_L g6447 ( 
.A(n_6315),
.B(n_6073),
.Y(n_6447)
);

OR2x2_ASAP7_75t_L g6448 ( 
.A(n_6300),
.B(n_6330),
.Y(n_6448)
);

AND2x2_ASAP7_75t_L g6449 ( 
.A(n_6313),
.B(n_6354),
.Y(n_6449)
);

OR2x2_ASAP7_75t_L g6450 ( 
.A(n_6326),
.B(n_6082),
.Y(n_6450)
);

HB1xp67_ASAP7_75t_L g6451 ( 
.A(n_6357),
.Y(n_6451)
);

OR2x2_ASAP7_75t_L g6452 ( 
.A(n_6302),
.B(n_6085),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_6416),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_6427),
.Y(n_6454)
);

AND2x2_ASAP7_75t_L g6455 ( 
.A(n_6449),
.B(n_6371),
.Y(n_6455)
);

NOR2x1p5_ASAP7_75t_L g6456 ( 
.A(n_6420),
.B(n_6438),
.Y(n_6456)
);

INVx1_ASAP7_75t_L g6457 ( 
.A(n_6425),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6448),
.Y(n_6458)
);

NAND2xp33_ASAP7_75t_L g6459 ( 
.A(n_6451),
.B(n_6325),
.Y(n_6459)
);

AND2x2_ASAP7_75t_L g6460 ( 
.A(n_6395),
.B(n_6348),
.Y(n_6460)
);

NAND2xp5_ASAP7_75t_L g6461 ( 
.A(n_6437),
.B(n_6316),
.Y(n_6461)
);

INVx1_ASAP7_75t_SL g6462 ( 
.A(n_6415),
.Y(n_6462)
);

INVxp67_ASAP7_75t_L g6463 ( 
.A(n_6436),
.Y(n_6463)
);

NAND2xp5_ASAP7_75t_L g6464 ( 
.A(n_6408),
.B(n_6407),
.Y(n_6464)
);

AND2x2_ASAP7_75t_SL g6465 ( 
.A(n_6399),
.B(n_6418),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_6409),
.B(n_6318),
.Y(n_6466)
);

NOR2xp33_ASAP7_75t_R g6467 ( 
.A(n_6413),
.B(n_6337),
.Y(n_6467)
);

INVx2_ASAP7_75t_L g6468 ( 
.A(n_6400),
.Y(n_6468)
);

INVx1_ASAP7_75t_L g6469 ( 
.A(n_6396),
.Y(n_6469)
);

INVx2_ASAP7_75t_L g6470 ( 
.A(n_6447),
.Y(n_6470)
);

NAND2xp5_ASAP7_75t_L g6471 ( 
.A(n_6429),
.B(n_6443),
.Y(n_6471)
);

AND2x2_ASAP7_75t_L g6472 ( 
.A(n_6401),
.B(n_6340),
.Y(n_6472)
);

OAI22xp5_ASAP7_75t_L g6473 ( 
.A1(n_6433),
.A2(n_6373),
.B1(n_6387),
.B2(n_6388),
.Y(n_6473)
);

INVx1_ASAP7_75t_L g6474 ( 
.A(n_6397),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_6426),
.Y(n_6475)
);

OAI31xp33_ASAP7_75t_L g6476 ( 
.A1(n_6410),
.A2(n_6355),
.A3(n_6385),
.B(n_6386),
.Y(n_6476)
);

AND2x2_ASAP7_75t_L g6477 ( 
.A(n_6435),
.B(n_6345),
.Y(n_6477)
);

NAND2xp5_ASAP7_75t_SL g6478 ( 
.A(n_6398),
.B(n_6368),
.Y(n_6478)
);

INVx1_ASAP7_75t_L g6479 ( 
.A(n_6450),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_6423),
.Y(n_6480)
);

INVx1_ASAP7_75t_L g6481 ( 
.A(n_6424),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_6446),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6412),
.B(n_6350),
.Y(n_6483)
);

NOR2xp33_ASAP7_75t_L g6484 ( 
.A(n_6394),
.B(n_6392),
.Y(n_6484)
);

OR2x2_ASAP7_75t_L g6485 ( 
.A(n_6440),
.B(n_6331),
.Y(n_6485)
);

AND2x2_ASAP7_75t_L g6486 ( 
.A(n_6434),
.B(n_6352),
.Y(n_6486)
);

INVx2_ASAP7_75t_L g6487 ( 
.A(n_6428),
.Y(n_6487)
);

INVxp67_ASAP7_75t_L g6488 ( 
.A(n_6411),
.Y(n_6488)
);

INVxp67_ASAP7_75t_SL g6489 ( 
.A(n_6405),
.Y(n_6489)
);

BUFx3_ASAP7_75t_L g6490 ( 
.A(n_6403),
.Y(n_6490)
);

INVxp67_ASAP7_75t_L g6491 ( 
.A(n_6422),
.Y(n_6491)
);

NAND2xp5_ASAP7_75t_L g6492 ( 
.A(n_6414),
.B(n_6382),
.Y(n_6492)
);

INVx1_ASAP7_75t_L g6493 ( 
.A(n_6452),
.Y(n_6493)
);

NOR2xp33_ASAP7_75t_L g6494 ( 
.A(n_6417),
.B(n_6336),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6406),
.B(n_6353),
.Y(n_6495)
);

INVx1_ASAP7_75t_SL g6496 ( 
.A(n_6402),
.Y(n_6496)
);

NOR2xp33_ASAP7_75t_L g6497 ( 
.A(n_6404),
.B(n_6314),
.Y(n_6497)
);

NAND4xp25_ASAP7_75t_L g6498 ( 
.A(n_6490),
.B(n_6431),
.C(n_6442),
.D(n_6441),
.Y(n_6498)
);

CKINVDCx16_ASAP7_75t_R g6499 ( 
.A(n_6460),
.Y(n_6499)
);

INVx1_ASAP7_75t_L g6500 ( 
.A(n_6464),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_6455),
.Y(n_6501)
);

NAND2xp5_ASAP7_75t_L g6502 ( 
.A(n_6477),
.B(n_6432),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_6492),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6457),
.Y(n_6504)
);

INVx2_ASAP7_75t_SL g6505 ( 
.A(n_6456),
.Y(n_6505)
);

AND2x2_ASAP7_75t_L g6506 ( 
.A(n_6468),
.B(n_6430),
.Y(n_6506)
);

OR2x2_ASAP7_75t_L g6507 ( 
.A(n_6458),
.B(n_6444),
.Y(n_6507)
);

NAND2xp5_ASAP7_75t_L g6508 ( 
.A(n_6470),
.B(n_6482),
.Y(n_6508)
);

AND2x4_ASAP7_75t_L g6509 ( 
.A(n_6472),
.B(n_6309),
.Y(n_6509)
);

INVx2_ASAP7_75t_L g6510 ( 
.A(n_6485),
.Y(n_6510)
);

AND2x2_ASAP7_75t_L g6511 ( 
.A(n_6483),
.B(n_6359),
.Y(n_6511)
);

INVxp67_ASAP7_75t_L g6512 ( 
.A(n_6494),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_6466),
.Y(n_6513)
);

AND2x4_ASAP7_75t_L g6514 ( 
.A(n_6454),
.B(n_6323),
.Y(n_6514)
);

NAND2xp5_ASAP7_75t_L g6515 ( 
.A(n_6497),
.B(n_6381),
.Y(n_6515)
);

INVx2_ASAP7_75t_L g6516 ( 
.A(n_6465),
.Y(n_6516)
);

INVxp33_ASAP7_75t_L g6517 ( 
.A(n_6478),
.Y(n_6517)
);

HB1xp67_ASAP7_75t_L g6518 ( 
.A(n_6463),
.Y(n_6518)
);

INVx1_ASAP7_75t_L g6519 ( 
.A(n_6486),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_6461),
.Y(n_6520)
);

NOR3x1_ASAP7_75t_L g6521 ( 
.A(n_6489),
.B(n_6421),
.C(n_6419),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_6479),
.Y(n_6522)
);

NAND2xp5_ASAP7_75t_L g6523 ( 
.A(n_6493),
.B(n_6445),
.Y(n_6523)
);

AND2x2_ASAP7_75t_L g6524 ( 
.A(n_6475),
.B(n_6361),
.Y(n_6524)
);

AND2x4_ASAP7_75t_L g6525 ( 
.A(n_6487),
.B(n_6356),
.Y(n_6525)
);

INVx2_ASAP7_75t_L g6526 ( 
.A(n_6495),
.Y(n_6526)
);

INVx2_ASAP7_75t_L g6527 ( 
.A(n_6496),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_L g6528 ( 
.A(n_6462),
.B(n_6484),
.Y(n_6528)
);

AND2x2_ASAP7_75t_L g6529 ( 
.A(n_6453),
.B(n_6365),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_6469),
.Y(n_6530)
);

OAI21xp5_ASAP7_75t_L g6531 ( 
.A1(n_6473),
.A2(n_6390),
.B(n_6439),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6459),
.B(n_6367),
.Y(n_6532)
);

OR2x2_ASAP7_75t_L g6533 ( 
.A(n_6491),
.B(n_6370),
.Y(n_6533)
);

AOI22xp5_ASAP7_75t_L g6534 ( 
.A1(n_6471),
.A2(n_6364),
.B1(n_6380),
.B2(n_6378),
.Y(n_6534)
);

INVx2_ASAP7_75t_L g6535 ( 
.A(n_6474),
.Y(n_6535)
);

INVx1_ASAP7_75t_SL g6536 ( 
.A(n_6467),
.Y(n_6536)
);

OAI21xp5_ASAP7_75t_L g6537 ( 
.A1(n_6476),
.A2(n_6375),
.B(n_6372),
.Y(n_6537)
);

OAI22xp33_ASAP7_75t_L g6538 ( 
.A1(n_6488),
.A2(n_6219),
.B1(n_6243),
.B2(n_6087),
.Y(n_6538)
);

NAND2xp5_ASAP7_75t_L g6539 ( 
.A(n_6480),
.B(n_6249),
.Y(n_6539)
);

AOI31xp33_ASAP7_75t_L g6540 ( 
.A1(n_6481),
.A2(n_6252),
.A3(n_6291),
.B(n_6255),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6464),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_6464),
.Y(n_6542)
);

NAND2xp5_ASAP7_75t_L g6543 ( 
.A(n_6455),
.B(n_6086),
.Y(n_6543)
);

AOI311xp33_ASAP7_75t_L g6544 ( 
.A1(n_6457),
.A2(n_6067),
.A3(n_6084),
.B(n_6088),
.C(n_6079),
.Y(n_6544)
);

INVx1_ASAP7_75t_L g6545 ( 
.A(n_6464),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_6518),
.Y(n_6546)
);

NAND2xp5_ASAP7_75t_L g6547 ( 
.A(n_6499),
.B(n_6506),
.Y(n_6547)
);

AOI22xp33_ASAP7_75t_L g6548 ( 
.A1(n_6516),
.A2(n_803),
.B1(n_801),
.B2(n_802),
.Y(n_6548)
);

BUFx3_ASAP7_75t_L g6549 ( 
.A(n_6509),
.Y(n_6549)
);

INVx1_ASAP7_75t_L g6550 ( 
.A(n_6511),
.Y(n_6550)
);

AND2x2_ASAP7_75t_L g6551 ( 
.A(n_6510),
.B(n_801),
.Y(n_6551)
);

BUFx6f_ASAP7_75t_L g6552 ( 
.A(n_6527),
.Y(n_6552)
);

INVx1_ASAP7_75t_L g6553 ( 
.A(n_6501),
.Y(n_6553)
);

INVx5_ASAP7_75t_L g6554 ( 
.A(n_6505),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_6526),
.B(n_802),
.Y(n_6555)
);

INVx1_ASAP7_75t_L g6556 ( 
.A(n_6525),
.Y(n_6556)
);

INVx1_ASAP7_75t_SL g6557 ( 
.A(n_6528),
.Y(n_6557)
);

NAND2xp5_ASAP7_75t_L g6558 ( 
.A(n_6512),
.B(n_804),
.Y(n_6558)
);

INVx1_ASAP7_75t_L g6559 ( 
.A(n_6519),
.Y(n_6559)
);

HB1xp67_ASAP7_75t_L g6560 ( 
.A(n_6536),
.Y(n_6560)
);

NAND2xp5_ASAP7_75t_L g6561 ( 
.A(n_6517),
.B(n_805),
.Y(n_6561)
);

INVx2_ASAP7_75t_L g6562 ( 
.A(n_6507),
.Y(n_6562)
);

CKINVDCx16_ASAP7_75t_R g6563 ( 
.A(n_6531),
.Y(n_6563)
);

INVx1_ASAP7_75t_SL g6564 ( 
.A(n_6533),
.Y(n_6564)
);

NAND3xp33_ASAP7_75t_SL g6565 ( 
.A(n_6537),
.B(n_6534),
.C(n_6515),
.Y(n_6565)
);

OAI21x1_ASAP7_75t_L g6566 ( 
.A1(n_6523),
.A2(n_805),
.B(n_807),
.Y(n_6566)
);

NOR2xp33_ASAP7_75t_L g6567 ( 
.A(n_6500),
.B(n_807),
.Y(n_6567)
);

INVx1_ASAP7_75t_L g6568 ( 
.A(n_6541),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6542),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_6545),
.Y(n_6570)
);

INVx1_ASAP7_75t_L g6571 ( 
.A(n_6543),
.Y(n_6571)
);

NOR2xp33_ASAP7_75t_L g6572 ( 
.A(n_6513),
.B(n_808),
.Y(n_6572)
);

INVx1_ASAP7_75t_L g6573 ( 
.A(n_6503),
.Y(n_6573)
);

INVxp33_ASAP7_75t_L g6574 ( 
.A(n_6498),
.Y(n_6574)
);

INVx4_ASAP7_75t_L g6575 ( 
.A(n_6514),
.Y(n_6575)
);

OAI21x1_ASAP7_75t_L g6576 ( 
.A1(n_6502),
.A2(n_808),
.B(n_810),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6524),
.Y(n_6577)
);

AND2x2_ASAP7_75t_L g6578 ( 
.A(n_6520),
.B(n_811),
.Y(n_6578)
);

NAND2xp5_ASAP7_75t_L g6579 ( 
.A(n_6521),
.B(n_6532),
.Y(n_6579)
);

OR2x2_ASAP7_75t_L g6580 ( 
.A(n_6508),
.B(n_811),
.Y(n_6580)
);

INVx1_ASAP7_75t_SL g6581 ( 
.A(n_6529),
.Y(n_6581)
);

AND2x2_ASAP7_75t_L g6582 ( 
.A(n_6522),
.B(n_812),
.Y(n_6582)
);

AOI22xp33_ASAP7_75t_L g6583 ( 
.A1(n_6538),
.A2(n_6539),
.B1(n_6530),
.B2(n_6535),
.Y(n_6583)
);

NOR2xp33_ASAP7_75t_SL g6584 ( 
.A(n_6504),
.B(n_812),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_SL g6585 ( 
.A(n_6544),
.B(n_813),
.Y(n_6585)
);

NAND2xp5_ASAP7_75t_L g6586 ( 
.A(n_6540),
.B(n_813),
.Y(n_6586)
);

OR2x2_ASAP7_75t_L g6587 ( 
.A(n_6499),
.B(n_814),
.Y(n_6587)
);

OAI21x1_ASAP7_75t_L g6588 ( 
.A1(n_6516),
.A2(n_814),
.B(n_815),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_6518),
.Y(n_6589)
);

HB1xp67_ASAP7_75t_L g6590 ( 
.A(n_6499),
.Y(n_6590)
);

NOR2x1_ASAP7_75t_L g6591 ( 
.A(n_6528),
.B(n_815),
.Y(n_6591)
);

INVx2_ASAP7_75t_L g6592 ( 
.A(n_6499),
.Y(n_6592)
);

NOR2xp33_ASAP7_75t_SL g6593 ( 
.A(n_6499),
.B(n_816),
.Y(n_6593)
);

INVx1_ASAP7_75t_SL g6594 ( 
.A(n_6499),
.Y(n_6594)
);

INVxp67_ASAP7_75t_L g6595 ( 
.A(n_6518),
.Y(n_6595)
);

AND2x2_ASAP7_75t_L g6596 ( 
.A(n_6499),
.B(n_816),
.Y(n_6596)
);

NOR2xp33_ASAP7_75t_L g6597 ( 
.A(n_6499),
.B(n_817),
.Y(n_6597)
);

NAND2xp5_ASAP7_75t_L g6598 ( 
.A(n_6499),
.B(n_818),
.Y(n_6598)
);

OAI221xp5_ASAP7_75t_L g6599 ( 
.A1(n_6531),
.A2(n_820),
.B1(n_818),
.B2(n_819),
.C(n_821),
.Y(n_6599)
);

OR2x2_ASAP7_75t_L g6600 ( 
.A(n_6499),
.B(n_820),
.Y(n_6600)
);

CKINVDCx16_ASAP7_75t_R g6601 ( 
.A(n_6499),
.Y(n_6601)
);

OR2x2_ASAP7_75t_L g6602 ( 
.A(n_6499),
.B(n_822),
.Y(n_6602)
);

HB1xp67_ASAP7_75t_L g6603 ( 
.A(n_6499),
.Y(n_6603)
);

NAND2xp5_ASAP7_75t_L g6604 ( 
.A(n_6499),
.B(n_823),
.Y(n_6604)
);

INVx1_ASAP7_75t_L g6605 ( 
.A(n_6518),
.Y(n_6605)
);

INVx2_ASAP7_75t_SL g6606 ( 
.A(n_6601),
.Y(n_6606)
);

OAI21xp33_ASAP7_75t_L g6607 ( 
.A1(n_6594),
.A2(n_823),
.B(n_824),
.Y(n_6607)
);

INVx1_ASAP7_75t_L g6608 ( 
.A(n_6590),
.Y(n_6608)
);

NOR2xp33_ASAP7_75t_SL g6609 ( 
.A(n_6575),
.B(n_824),
.Y(n_6609)
);

NOR3xp33_ASAP7_75t_L g6610 ( 
.A(n_6563),
.B(n_6603),
.C(n_6565),
.Y(n_6610)
);

NOR2xp33_ASAP7_75t_L g6611 ( 
.A(n_6547),
.B(n_825),
.Y(n_6611)
);

OAI22xp5_ASAP7_75t_L g6612 ( 
.A1(n_6595),
.A2(n_827),
.B1(n_825),
.B2(n_826),
.Y(n_6612)
);

AND2x2_ASAP7_75t_SL g6613 ( 
.A(n_6596),
.B(n_828),
.Y(n_6613)
);

AO21x1_ASAP7_75t_L g6614 ( 
.A1(n_6585),
.A2(n_828),
.B(n_829),
.Y(n_6614)
);

AOI332xp33_ASAP7_75t_L g6615 ( 
.A1(n_6546),
.A2(n_6589),
.A3(n_6605),
.B1(n_6592),
.B2(n_6553),
.B3(n_6550),
.C1(n_6559),
.C2(n_6577),
.Y(n_6615)
);

INVx1_ASAP7_75t_L g6616 ( 
.A(n_6587),
.Y(n_6616)
);

AOI22x1_ASAP7_75t_L g6617 ( 
.A1(n_6560),
.A2(n_831),
.B1(n_829),
.B2(n_830),
.Y(n_6617)
);

INVx1_ASAP7_75t_SL g6618 ( 
.A(n_6600),
.Y(n_6618)
);

OAI322xp33_ASAP7_75t_L g6619 ( 
.A1(n_6579),
.A2(n_835),
.A3(n_834),
.B1(n_832),
.B2(n_830),
.C1(n_831),
.C2(n_833),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_L g6620 ( 
.A(n_6549),
.B(n_833),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_6602),
.Y(n_6621)
);

OAI31xp33_ASAP7_75t_SL g6622 ( 
.A1(n_6581),
.A2(n_836),
.A3(n_834),
.B(n_835),
.Y(n_6622)
);

INVxp33_ASAP7_75t_L g6623 ( 
.A(n_6597),
.Y(n_6623)
);

NAND2xp5_ASAP7_75t_L g6624 ( 
.A(n_6591),
.B(n_836),
.Y(n_6624)
);

XNOR2x1_ASAP7_75t_L g6625 ( 
.A(n_6557),
.B(n_837),
.Y(n_6625)
);

NAND2xp5_ASAP7_75t_L g6626 ( 
.A(n_6593),
.B(n_839),
.Y(n_6626)
);

NOR2x1_ASAP7_75t_L g6627 ( 
.A(n_6598),
.B(n_839),
.Y(n_6627)
);

OAI21xp33_ASAP7_75t_L g6628 ( 
.A1(n_6574),
.A2(n_840),
.B(n_841),
.Y(n_6628)
);

AND2x4_ASAP7_75t_L g6629 ( 
.A(n_6554),
.B(n_840),
.Y(n_6629)
);

OAI221xp5_ASAP7_75t_L g6630 ( 
.A1(n_6583),
.A2(n_843),
.B1(n_841),
.B2(n_842),
.C(n_844),
.Y(n_6630)
);

OAI221xp5_ASAP7_75t_L g6631 ( 
.A1(n_6604),
.A2(n_845),
.B1(n_843),
.B2(n_844),
.C(n_846),
.Y(n_6631)
);

INVx1_ASAP7_75t_L g6632 ( 
.A(n_6556),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_6552),
.Y(n_6633)
);

AOI221xp5_ASAP7_75t_L g6634 ( 
.A1(n_6586),
.A2(n_847),
.B1(n_845),
.B2(n_846),
.C(n_848),
.Y(n_6634)
);

AOI22xp33_ASAP7_75t_SL g6635 ( 
.A1(n_6562),
.A2(n_856),
.B1(n_864),
.B2(n_847),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_6552),
.Y(n_6636)
);

AOI21xp5_ASAP7_75t_L g6637 ( 
.A1(n_6561),
.A2(n_849),
.B(n_850),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_6551),
.B(n_849),
.Y(n_6638)
);

NOR3xp33_ASAP7_75t_SL g6639 ( 
.A(n_6568),
.B(n_850),
.C(n_851),
.Y(n_6639)
);

NAND2xp5_ASAP7_75t_L g6640 ( 
.A(n_6555),
.B(n_851),
.Y(n_6640)
);

NOR4xp25_ASAP7_75t_SL g6641 ( 
.A(n_6569),
.B(n_854),
.C(n_852),
.D(n_853),
.Y(n_6641)
);

AOI22xp33_ASAP7_75t_L g6642 ( 
.A1(n_6572),
.A2(n_855),
.B1(n_853),
.B2(n_854),
.Y(n_6642)
);

INVx1_ASAP7_75t_L g6643 ( 
.A(n_6578),
.Y(n_6643)
);

A2O1A1Ixp33_ASAP7_75t_L g6644 ( 
.A1(n_6567),
.A2(n_857),
.B(n_855),
.C(n_856),
.Y(n_6644)
);

OAI221xp5_ASAP7_75t_L g6645 ( 
.A1(n_6584),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.C(n_860),
.Y(n_6645)
);

O2A1O1Ixp33_ASAP7_75t_L g6646 ( 
.A1(n_6564),
.A2(n_860),
.B(n_858),
.C(n_859),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6582),
.Y(n_6647)
);

INVx1_ASAP7_75t_L g6648 ( 
.A(n_6580),
.Y(n_6648)
);

NAND3xp33_ASAP7_75t_SL g6649 ( 
.A(n_6571),
.B(n_861),
.C(n_862),
.Y(n_6649)
);

AOI21xp33_ASAP7_75t_L g6650 ( 
.A1(n_6573),
.A2(n_1799),
.B(n_1798),
.Y(n_6650)
);

INVx2_ASAP7_75t_L g6651 ( 
.A(n_6576),
.Y(n_6651)
);

AND2x2_ASAP7_75t_L g6652 ( 
.A(n_6554),
.B(n_861),
.Y(n_6652)
);

OAI21xp33_ASAP7_75t_L g6653 ( 
.A1(n_6570),
.A2(n_862),
.B(n_863),
.Y(n_6653)
);

INVx2_ASAP7_75t_L g6654 ( 
.A(n_6588),
.Y(n_6654)
);

INVx2_ASAP7_75t_L g6655 ( 
.A(n_6554),
.Y(n_6655)
);

AOI211x1_ASAP7_75t_L g6656 ( 
.A1(n_6599),
.A2(n_865),
.B(n_863),
.C(n_864),
.Y(n_6656)
);

O2A1O1Ixp33_ASAP7_75t_L g6657 ( 
.A1(n_6558),
.A2(n_868),
.B(n_866),
.C(n_867),
.Y(n_6657)
);

INVx2_ASAP7_75t_L g6658 ( 
.A(n_6566),
.Y(n_6658)
);

INVx1_ASAP7_75t_L g6659 ( 
.A(n_6548),
.Y(n_6659)
);

INVx1_ASAP7_75t_L g6660 ( 
.A(n_6590),
.Y(n_6660)
);

OAI32xp33_ASAP7_75t_L g6661 ( 
.A1(n_6601),
.A2(n_868),
.A3(n_866),
.B1(n_867),
.B2(n_869),
.Y(n_6661)
);

NOR2xp67_ASAP7_75t_L g6662 ( 
.A(n_6575),
.B(n_871),
.Y(n_6662)
);

NAND2xp5_ASAP7_75t_SL g6663 ( 
.A(n_6601),
.B(n_871),
.Y(n_6663)
);

NAND2xp5_ASAP7_75t_L g6664 ( 
.A(n_6601),
.B(n_872),
.Y(n_6664)
);

INVx4_ASAP7_75t_L g6665 ( 
.A(n_6554),
.Y(n_6665)
);

OAI21xp33_ASAP7_75t_L g6666 ( 
.A1(n_6594),
.A2(n_872),
.B(n_873),
.Y(n_6666)
);

HB1xp67_ASAP7_75t_L g6667 ( 
.A(n_6601),
.Y(n_6667)
);

OA21x2_ASAP7_75t_L g6668 ( 
.A1(n_6585),
.A2(n_873),
.B(n_874),
.Y(n_6668)
);

INVx1_ASAP7_75t_L g6669 ( 
.A(n_6590),
.Y(n_6669)
);

NAND3xp33_ASAP7_75t_L g6670 ( 
.A(n_6590),
.B(n_885),
.C(n_875),
.Y(n_6670)
);

NOR3xp33_ASAP7_75t_SL g6671 ( 
.A(n_6601),
.B(n_875),
.C(n_876),
.Y(n_6671)
);

OAI221xp5_ASAP7_75t_L g6672 ( 
.A1(n_6594),
.A2(n_880),
.B1(n_878),
.B2(n_879),
.C(n_881),
.Y(n_6672)
);

AND2x2_ASAP7_75t_L g6673 ( 
.A(n_6601),
.B(n_878),
.Y(n_6673)
);

AND2x2_ASAP7_75t_L g6674 ( 
.A(n_6601),
.B(n_879),
.Y(n_6674)
);

OAI21xp33_ASAP7_75t_L g6675 ( 
.A1(n_6594),
.A2(n_881),
.B(n_882),
.Y(n_6675)
);

OAI22xp33_ASAP7_75t_L g6676 ( 
.A1(n_6601),
.A2(n_885),
.B1(n_882),
.B2(n_884),
.Y(n_6676)
);

NOR2xp33_ASAP7_75t_SL g6677 ( 
.A(n_6601),
.B(n_884),
.Y(n_6677)
);

INVxp33_ASAP7_75t_L g6678 ( 
.A(n_6590),
.Y(n_6678)
);

AOI221xp5_ASAP7_75t_L g6679 ( 
.A1(n_6565),
.A2(n_888),
.B1(n_886),
.B2(n_887),
.C(n_889),
.Y(n_6679)
);

AOI211xp5_ASAP7_75t_L g6680 ( 
.A1(n_6594),
.A2(n_888),
.B(n_886),
.C(n_887),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_6590),
.Y(n_6681)
);

AOI21xp5_ASAP7_75t_L g6682 ( 
.A1(n_6547),
.A2(n_889),
.B(n_890),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_6590),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6590),
.Y(n_6684)
);

INVx2_ASAP7_75t_L g6685 ( 
.A(n_6601),
.Y(n_6685)
);

AND2x4_ASAP7_75t_L g6686 ( 
.A(n_6575),
.B(n_890),
.Y(n_6686)
);

NAND2xp5_ASAP7_75t_L g6687 ( 
.A(n_6601),
.B(n_891),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_SL g6688 ( 
.A(n_6601),
.B(n_892),
.Y(n_6688)
);

OAI22xp5_ASAP7_75t_L g6689 ( 
.A1(n_6601),
.A2(n_894),
.B1(n_892),
.B2(n_893),
.Y(n_6689)
);

NAND2xp5_ASAP7_75t_L g6690 ( 
.A(n_6601),
.B(n_893),
.Y(n_6690)
);

OAI222xp33_ASAP7_75t_L g6691 ( 
.A1(n_6594),
.A2(n_896),
.B1(n_898),
.B2(n_894),
.C1(n_895),
.C2(n_897),
.Y(n_6691)
);

NAND2xp5_ASAP7_75t_L g6692 ( 
.A(n_6601),
.B(n_895),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6590),
.Y(n_6693)
);

NAND2xp5_ASAP7_75t_L g6694 ( 
.A(n_6601),
.B(n_896),
.Y(n_6694)
);

INVx2_ASAP7_75t_L g6695 ( 
.A(n_6601),
.Y(n_6695)
);

NAND2xp5_ASAP7_75t_SL g6696 ( 
.A(n_6601),
.B(n_897),
.Y(n_6696)
);

AO22x1_ASAP7_75t_L g6697 ( 
.A1(n_6590),
.A2(n_900),
.B1(n_898),
.B2(n_899),
.Y(n_6697)
);

NAND2x1_ASAP7_75t_L g6698 ( 
.A(n_6575),
.B(n_900),
.Y(n_6698)
);

INVx2_ASAP7_75t_SL g6699 ( 
.A(n_6601),
.Y(n_6699)
);

NAND3xp33_ASAP7_75t_L g6700 ( 
.A(n_6590),
.B(n_910),
.C(n_901),
.Y(n_6700)
);

INVx1_ASAP7_75t_SL g6701 ( 
.A(n_6601),
.Y(n_6701)
);

OAI322xp33_ASAP7_75t_L g6702 ( 
.A1(n_6701),
.A2(n_6699),
.A3(n_6606),
.B1(n_6695),
.B2(n_6685),
.C1(n_6669),
.C2(n_6660),
.Y(n_6702)
);

OAI221xp5_ASAP7_75t_L g6703 ( 
.A1(n_6667),
.A2(n_903),
.B1(n_901),
.B2(n_902),
.C(n_905),
.Y(n_6703)
);

OAI222xp33_ASAP7_75t_L g6704 ( 
.A1(n_6618),
.A2(n_906),
.B1(n_908),
.B2(n_902),
.C1(n_903),
.C2(n_907),
.Y(n_6704)
);

AND2x2_ASAP7_75t_L g6705 ( 
.A(n_6673),
.B(n_6674),
.Y(n_6705)
);

HB1xp67_ASAP7_75t_L g6706 ( 
.A(n_6662),
.Y(n_6706)
);

AND2x4_ASAP7_75t_L g6707 ( 
.A(n_6652),
.B(n_6665),
.Y(n_6707)
);

AOI21xp5_ASAP7_75t_L g6708 ( 
.A1(n_6698),
.A2(n_907),
.B(n_908),
.Y(n_6708)
);

OAI21xp33_ASAP7_75t_SL g6709 ( 
.A1(n_6633),
.A2(n_909),
.B(n_911),
.Y(n_6709)
);

AOI22xp33_ASAP7_75t_L g6710 ( 
.A1(n_6614),
.A2(n_912),
.B1(n_909),
.B2(n_911),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6610),
.B(n_912),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_6625),
.Y(n_6712)
);

NAND3xp33_ASAP7_75t_L g6713 ( 
.A(n_6677),
.B(n_913),
.C(n_914),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_6629),
.Y(n_6714)
);

NAND2xp5_ASAP7_75t_L g6715 ( 
.A(n_6697),
.B(n_913),
.Y(n_6715)
);

AOI221xp5_ASAP7_75t_L g6716 ( 
.A1(n_6616),
.A2(n_916),
.B1(n_914),
.B2(n_915),
.C(n_917),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6678),
.B(n_915),
.Y(n_6717)
);

OAI22xp5_ASAP7_75t_L g6718 ( 
.A1(n_6664),
.A2(n_919),
.B1(n_916),
.B2(n_918),
.Y(n_6718)
);

OAI22xp33_ASAP7_75t_L g6719 ( 
.A1(n_6687),
.A2(n_921),
.B1(n_918),
.B2(n_920),
.Y(n_6719)
);

AND2x2_ASAP7_75t_L g6720 ( 
.A(n_6636),
.B(n_920),
.Y(n_6720)
);

INVx1_ASAP7_75t_L g6721 ( 
.A(n_6629),
.Y(n_6721)
);

INVx1_ASAP7_75t_L g6722 ( 
.A(n_6613),
.Y(n_6722)
);

NOR3xp33_ASAP7_75t_L g6723 ( 
.A(n_6690),
.B(n_921),
.C(n_922),
.Y(n_6723)
);

NOR2xp33_ASAP7_75t_L g6724 ( 
.A(n_6691),
.B(n_1790),
.Y(n_6724)
);

NOR2x1_ASAP7_75t_L g6725 ( 
.A(n_6692),
.B(n_922),
.Y(n_6725)
);

NAND2xp5_ASAP7_75t_L g6726 ( 
.A(n_6622),
.B(n_923),
.Y(n_6726)
);

OAI21xp33_ASAP7_75t_SL g6727 ( 
.A1(n_6608),
.A2(n_923),
.B(n_924),
.Y(n_6727)
);

INVx1_ASAP7_75t_L g6728 ( 
.A(n_6694),
.Y(n_6728)
);

INVxp67_ASAP7_75t_L g6729 ( 
.A(n_6609),
.Y(n_6729)
);

NAND2xp5_ASAP7_75t_L g6730 ( 
.A(n_6686),
.B(n_6671),
.Y(n_6730)
);

NAND2x1p5_ASAP7_75t_L g6731 ( 
.A(n_6663),
.B(n_926),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6627),
.Y(n_6732)
);

AOI22xp5_ASAP7_75t_L g6733 ( 
.A1(n_6621),
.A2(n_927),
.B1(n_925),
.B2(n_926),
.Y(n_6733)
);

INVx2_ASAP7_75t_L g6734 ( 
.A(n_6617),
.Y(n_6734)
);

AOI22xp33_ASAP7_75t_L g6735 ( 
.A1(n_6658),
.A2(n_928),
.B1(n_925),
.B2(n_927),
.Y(n_6735)
);

AOI221xp5_ASAP7_75t_L g6736 ( 
.A1(n_6623),
.A2(n_930),
.B1(n_928),
.B2(n_929),
.C(n_931),
.Y(n_6736)
);

INVx2_ASAP7_75t_L g6737 ( 
.A(n_6655),
.Y(n_6737)
);

AOI31xp33_ASAP7_75t_L g6738 ( 
.A1(n_6681),
.A2(n_932),
.A3(n_930),
.B(n_931),
.Y(n_6738)
);

AOI22xp5_ASAP7_75t_L g6739 ( 
.A1(n_6668),
.A2(n_935),
.B1(n_933),
.B2(n_934),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6624),
.Y(n_6740)
);

AOI22xp33_ASAP7_75t_L g6741 ( 
.A1(n_6651),
.A2(n_936),
.B1(n_933),
.B2(n_935),
.Y(n_6741)
);

AND2x2_ASAP7_75t_L g6742 ( 
.A(n_6683),
.B(n_936),
.Y(n_6742)
);

NAND2xp5_ASAP7_75t_L g6743 ( 
.A(n_6641),
.B(n_937),
.Y(n_6743)
);

INVxp33_ASAP7_75t_L g6744 ( 
.A(n_6611),
.Y(n_6744)
);

AOI22xp33_ASAP7_75t_L g6745 ( 
.A1(n_6654),
.A2(n_939),
.B1(n_937),
.B2(n_938),
.Y(n_6745)
);

HB1xp67_ASAP7_75t_L g6746 ( 
.A(n_6668),
.Y(n_6746)
);

NAND2xp5_ASAP7_75t_L g6747 ( 
.A(n_6639),
.B(n_6656),
.Y(n_6747)
);

AOI21xp5_ASAP7_75t_L g6748 ( 
.A1(n_6688),
.A2(n_6696),
.B(n_6646),
.Y(n_6748)
);

NAND2xp5_ASAP7_75t_L g6749 ( 
.A(n_6635),
.B(n_6643),
.Y(n_6749)
);

INVx1_ASAP7_75t_SL g6750 ( 
.A(n_6640),
.Y(n_6750)
);

INVx1_ASAP7_75t_L g6751 ( 
.A(n_6638),
.Y(n_6751)
);

NAND2xp5_ASAP7_75t_L g6752 ( 
.A(n_6648),
.B(n_939),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_6626),
.Y(n_6753)
);

NAND2xp5_ASAP7_75t_SL g6754 ( 
.A(n_6676),
.B(n_940),
.Y(n_6754)
);

NOR2xp33_ASAP7_75t_L g6755 ( 
.A(n_6619),
.B(n_1794),
.Y(n_6755)
);

A2O1A1Ixp33_ASAP7_75t_L g6756 ( 
.A1(n_6682),
.A2(n_943),
.B(n_941),
.C(n_942),
.Y(n_6756)
);

NAND2xp5_ASAP7_75t_L g6757 ( 
.A(n_6647),
.B(n_941),
.Y(n_6757)
);

INVx1_ASAP7_75t_L g6758 ( 
.A(n_6620),
.Y(n_6758)
);

AND2x4_ASAP7_75t_L g6759 ( 
.A(n_6684),
.B(n_6693),
.Y(n_6759)
);

AOI221xp5_ASAP7_75t_L g6760 ( 
.A1(n_6632),
.A2(n_944),
.B1(n_942),
.B2(n_943),
.C(n_945),
.Y(n_6760)
);

NOR2xp33_ASAP7_75t_L g6761 ( 
.A(n_6661),
.B(n_1805),
.Y(n_6761)
);

OR2x2_ASAP7_75t_L g6762 ( 
.A(n_6649),
.B(n_946),
.Y(n_6762)
);

NOR2xp33_ASAP7_75t_L g6763 ( 
.A(n_6630),
.B(n_1805),
.Y(n_6763)
);

NAND2xp5_ASAP7_75t_L g6764 ( 
.A(n_6680),
.B(n_946),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_6657),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_6670),
.Y(n_6766)
);

OAI21xp5_ASAP7_75t_SL g6767 ( 
.A1(n_6679),
.A2(n_947),
.B(n_948),
.Y(n_6767)
);

AOI21xp33_ASAP7_75t_SL g6768 ( 
.A1(n_6650),
.A2(n_1810),
.B(n_1809),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_6700),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6689),
.Y(n_6770)
);

AND2x2_ASAP7_75t_L g6771 ( 
.A(n_6607),
.B(n_947),
.Y(n_6771)
);

AND2x2_ASAP7_75t_L g6772 ( 
.A(n_6666),
.B(n_948),
.Y(n_6772)
);

OAI22xp33_ASAP7_75t_L g6773 ( 
.A1(n_6659),
.A2(n_952),
.B1(n_949),
.B2(n_951),
.Y(n_6773)
);

OAI221xp5_ASAP7_75t_L g6774 ( 
.A1(n_6628),
.A2(n_953),
.B1(n_949),
.B2(n_951),
.C(n_954),
.Y(n_6774)
);

OR2x2_ASAP7_75t_L g6775 ( 
.A(n_6675),
.B(n_953),
.Y(n_6775)
);

INVx1_ASAP7_75t_SL g6776 ( 
.A(n_6637),
.Y(n_6776)
);

AOI21xp5_ASAP7_75t_L g6777 ( 
.A1(n_6653),
.A2(n_954),
.B(n_956),
.Y(n_6777)
);

NAND2xp5_ASAP7_75t_SL g6778 ( 
.A(n_6634),
.B(n_957),
.Y(n_6778)
);

AND2x2_ASAP7_75t_L g6779 ( 
.A(n_6642),
.B(n_6644),
.Y(n_6779)
);

INVx1_ASAP7_75t_L g6780 ( 
.A(n_6612),
.Y(n_6780)
);

AOI22xp5_ASAP7_75t_L g6781 ( 
.A1(n_6631),
.A2(n_960),
.B1(n_958),
.B2(n_959),
.Y(n_6781)
);

AOI222xp33_ASAP7_75t_L g6782 ( 
.A1(n_6672),
.A2(n_963),
.B1(n_965),
.B2(n_966),
.C1(n_962),
.C2(n_964),
.Y(n_6782)
);

BUFx2_ASAP7_75t_L g6783 ( 
.A(n_6615),
.Y(n_6783)
);

AOI322xp5_ASAP7_75t_L g6784 ( 
.A1(n_6645),
.A2(n_967),
.A3(n_966),
.B1(n_964),
.B2(n_961),
.C1(n_963),
.C2(n_965),
.Y(n_6784)
);

NOR2xp33_ASAP7_75t_L g6785 ( 
.A(n_6701),
.B(n_961),
.Y(n_6785)
);

NAND2xp5_ASAP7_75t_L g6786 ( 
.A(n_6701),
.B(n_968),
.Y(n_6786)
);

NAND2xp33_ASAP7_75t_SL g6787 ( 
.A(n_6667),
.B(n_969),
.Y(n_6787)
);

OAI322xp33_ASAP7_75t_L g6788 ( 
.A1(n_6701),
.A2(n_974),
.A3(n_973),
.B1(n_971),
.B2(n_969),
.C1(n_970),
.C2(n_972),
.Y(n_6788)
);

AOI322xp5_ASAP7_75t_L g6789 ( 
.A1(n_6701),
.A2(n_975),
.A3(n_974),
.B1(n_972),
.B2(n_970),
.C1(n_971),
.C2(n_973),
.Y(n_6789)
);

AND2x2_ASAP7_75t_L g6790 ( 
.A(n_6667),
.B(n_975),
.Y(n_6790)
);

INVx1_ASAP7_75t_L g6791 ( 
.A(n_6667),
.Y(n_6791)
);

AOI332xp33_ASAP7_75t_L g6792 ( 
.A1(n_6608),
.A2(n_982),
.A3(n_980),
.B1(n_978),
.B2(n_983),
.B3(n_976),
.C1(n_977),
.C2(n_979),
.Y(n_6792)
);

OAI222xp33_ASAP7_75t_L g6793 ( 
.A1(n_6701),
.A2(n_980),
.B1(n_984),
.B2(n_976),
.C1(n_977),
.C2(n_982),
.Y(n_6793)
);

OAI32xp33_ASAP7_75t_L g6794 ( 
.A1(n_6701),
.A2(n_988),
.A3(n_985),
.B1(n_987),
.B2(n_989),
.Y(n_6794)
);

AOI22xp5_ASAP7_75t_L g6795 ( 
.A1(n_6701),
.A2(n_988),
.B1(n_985),
.B2(n_987),
.Y(n_6795)
);

INVxp67_ASAP7_75t_L g6796 ( 
.A(n_6667),
.Y(n_6796)
);

OAI22xp33_ASAP7_75t_L g6797 ( 
.A1(n_6701),
.A2(n_991),
.B1(n_989),
.B2(n_990),
.Y(n_6797)
);

INVx1_ASAP7_75t_SL g6798 ( 
.A(n_6701),
.Y(n_6798)
);

AOI32xp33_ASAP7_75t_L g6799 ( 
.A1(n_6701),
.A2(n_993),
.A3(n_990),
.B1(n_992),
.B2(n_994),
.Y(n_6799)
);

INVxp67_ASAP7_75t_SL g6800 ( 
.A(n_6667),
.Y(n_6800)
);

AOI22xp33_ASAP7_75t_L g6801 ( 
.A1(n_6706),
.A2(n_995),
.B1(n_992),
.B2(n_994),
.Y(n_6801)
);

NOR2xp33_ASAP7_75t_L g6802 ( 
.A(n_6709),
.B(n_995),
.Y(n_6802)
);

INVxp67_ASAP7_75t_L g6803 ( 
.A(n_6746),
.Y(n_6803)
);

NAND2xp5_ASAP7_75t_L g6804 ( 
.A(n_6798),
.B(n_996),
.Y(n_6804)
);

NOR2xp33_ASAP7_75t_L g6805 ( 
.A(n_6727),
.B(n_996),
.Y(n_6805)
);

AND2x2_ASAP7_75t_L g6806 ( 
.A(n_6800),
.B(n_6790),
.Y(n_6806)
);

INVx2_ASAP7_75t_SL g6807 ( 
.A(n_6707),
.Y(n_6807)
);

NAND2xp5_ASAP7_75t_L g6808 ( 
.A(n_6705),
.B(n_997),
.Y(n_6808)
);

INVx2_ASAP7_75t_L g6809 ( 
.A(n_6731),
.Y(n_6809)
);

OR2x2_ASAP7_75t_L g6810 ( 
.A(n_6783),
.B(n_997),
.Y(n_6810)
);

AND2x2_ASAP7_75t_L g6811 ( 
.A(n_6796),
.B(n_1807),
.Y(n_6811)
);

NOR2xp33_ASAP7_75t_L g6812 ( 
.A(n_6793),
.B(n_999),
.Y(n_6812)
);

AOI22xp33_ASAP7_75t_L g6813 ( 
.A1(n_6740),
.A2(n_1002),
.B1(n_1000),
.B2(n_1001),
.Y(n_6813)
);

BUFx2_ASAP7_75t_L g6814 ( 
.A(n_6787),
.Y(n_6814)
);

NAND2xp5_ASAP7_75t_L g6815 ( 
.A(n_6707),
.B(n_1000),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_6759),
.B(n_1002),
.Y(n_6816)
);

NOR2xp33_ASAP7_75t_L g6817 ( 
.A(n_6704),
.B(n_1003),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_L g6818 ( 
.A(n_6708),
.B(n_1003),
.Y(n_6818)
);

INVx1_ASAP7_75t_L g6819 ( 
.A(n_6743),
.Y(n_6819)
);

OR2x2_ASAP7_75t_L g6820 ( 
.A(n_6714),
.B(n_1004),
.Y(n_6820)
);

INVx2_ASAP7_75t_SL g6821 ( 
.A(n_6759),
.Y(n_6821)
);

NOR2xp33_ASAP7_75t_L g6822 ( 
.A(n_6744),
.B(n_1004),
.Y(n_6822)
);

AOI221xp5_ASAP7_75t_L g6823 ( 
.A1(n_6728),
.A2(n_1007),
.B1(n_1005),
.B2(n_1006),
.C(n_1008),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6732),
.Y(n_6824)
);

HB1xp67_ASAP7_75t_L g6825 ( 
.A(n_6721),
.Y(n_6825)
);

INVx2_ASAP7_75t_L g6826 ( 
.A(n_6725),
.Y(n_6826)
);

HB1xp67_ASAP7_75t_L g6827 ( 
.A(n_6730),
.Y(n_6827)
);

INVx1_ASAP7_75t_SL g6828 ( 
.A(n_6747),
.Y(n_6828)
);

AND2x4_ASAP7_75t_L g6829 ( 
.A(n_6791),
.B(n_1005),
.Y(n_6829)
);

INVx1_ASAP7_75t_L g6830 ( 
.A(n_6738),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_6720),
.Y(n_6831)
);

NAND2xp5_ASAP7_75t_L g6832 ( 
.A(n_6710),
.B(n_1006),
.Y(n_6832)
);

NAND2xp5_ASAP7_75t_L g6833 ( 
.A(n_6776),
.B(n_1007),
.Y(n_6833)
);

AND2x2_ASAP7_75t_L g6834 ( 
.A(n_6734),
.B(n_1792),
.Y(n_6834)
);

INVx2_ASAP7_75t_SL g6835 ( 
.A(n_6742),
.Y(n_6835)
);

AND2x2_ASAP7_75t_L g6836 ( 
.A(n_6717),
.B(n_1792),
.Y(n_6836)
);

AND2x2_ASAP7_75t_L g6837 ( 
.A(n_6711),
.B(n_1793),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6724),
.B(n_1008),
.Y(n_6838)
);

INVx1_ASAP7_75t_L g6839 ( 
.A(n_6715),
.Y(n_6839)
);

INVx1_ASAP7_75t_L g6840 ( 
.A(n_6726),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_6739),
.B(n_1009),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6785),
.B(n_1794),
.Y(n_6842)
);

NAND2xp5_ASAP7_75t_L g6843 ( 
.A(n_6799),
.B(n_1009),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_6722),
.Y(n_6844)
);

AOI22xp33_ASAP7_75t_L g6845 ( 
.A1(n_6750),
.A2(n_1012),
.B1(n_1010),
.B2(n_1011),
.Y(n_6845)
);

AND2x2_ASAP7_75t_L g6846 ( 
.A(n_6737),
.B(n_1800),
.Y(n_6846)
);

NAND2xp5_ASAP7_75t_L g6847 ( 
.A(n_6723),
.B(n_1011),
.Y(n_6847)
);

OR2x2_ASAP7_75t_L g6848 ( 
.A(n_6786),
.B(n_1013),
.Y(n_6848)
);

NAND2xp33_ASAP7_75t_L g6849 ( 
.A(n_6795),
.B(n_1013),
.Y(n_6849)
);

AND2x2_ASAP7_75t_L g6850 ( 
.A(n_6771),
.B(n_1826),
.Y(n_6850)
);

INVx2_ASAP7_75t_L g6851 ( 
.A(n_6762),
.Y(n_6851)
);

NAND2xp5_ASAP7_75t_L g6852 ( 
.A(n_6789),
.B(n_1014),
.Y(n_6852)
);

NAND2xp5_ASAP7_75t_L g6853 ( 
.A(n_6748),
.B(n_1014),
.Y(n_6853)
);

NAND2xp5_ASAP7_75t_L g6854 ( 
.A(n_6712),
.B(n_1015),
.Y(n_6854)
);

AND2x2_ASAP7_75t_L g6855 ( 
.A(n_6772),
.B(n_6766),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6702),
.Y(n_6856)
);

INVx1_ASAP7_75t_L g6857 ( 
.A(n_6752),
.Y(n_6857)
);

NOR2xp33_ASAP7_75t_L g6858 ( 
.A(n_6729),
.B(n_1015),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_L g6859 ( 
.A(n_6765),
.B(n_1016),
.Y(n_6859)
);

AND2x2_ASAP7_75t_L g6860 ( 
.A(n_6769),
.B(n_1783),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6755),
.B(n_1783),
.Y(n_6861)
);

INVx2_ASAP7_75t_L g6862 ( 
.A(n_6775),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_L g6863 ( 
.A(n_6756),
.B(n_1016),
.Y(n_6863)
);

INVxp67_ASAP7_75t_L g6864 ( 
.A(n_6761),
.Y(n_6864)
);

NAND2xp5_ASAP7_75t_L g6865 ( 
.A(n_6751),
.B(n_1017),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6757),
.Y(n_6866)
);

NAND2xp5_ASAP7_75t_L g6867 ( 
.A(n_6768),
.B(n_1017),
.Y(n_6867)
);

AND2x2_ASAP7_75t_L g6868 ( 
.A(n_6782),
.B(n_1786),
.Y(n_6868)
);

INVx1_ASAP7_75t_SL g6869 ( 
.A(n_6749),
.Y(n_6869)
);

NAND2xp33_ASAP7_75t_L g6870 ( 
.A(n_6764),
.B(n_1018),
.Y(n_6870)
);

AOI22xp33_ASAP7_75t_L g6871 ( 
.A1(n_6758),
.A2(n_1020),
.B1(n_1018),
.B2(n_1019),
.Y(n_6871)
);

HB1xp67_ASAP7_75t_SL g6872 ( 
.A(n_6703),
.Y(n_6872)
);

NAND2xp5_ASAP7_75t_L g6873 ( 
.A(n_6784),
.B(n_1019),
.Y(n_6873)
);

NOR2xp33_ASAP7_75t_SL g6874 ( 
.A(n_6788),
.B(n_1021),
.Y(n_6874)
);

INVx1_ASAP7_75t_L g6875 ( 
.A(n_6713),
.Y(n_6875)
);

AND2x2_ASAP7_75t_L g6876 ( 
.A(n_6770),
.B(n_1791),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6779),
.B(n_1022),
.Y(n_6877)
);

NOR2xp33_ASAP7_75t_L g6878 ( 
.A(n_6794),
.B(n_1022),
.Y(n_6878)
);

NOR2xp33_ASAP7_75t_L g6879 ( 
.A(n_6797),
.B(n_1023),
.Y(n_6879)
);

INVx1_ASAP7_75t_SL g6880 ( 
.A(n_6754),
.Y(n_6880)
);

INVx1_ASAP7_75t_SL g6881 ( 
.A(n_6753),
.Y(n_6881)
);

NOR2xp33_ASAP7_75t_L g6882 ( 
.A(n_6719),
.B(n_1023),
.Y(n_6882)
);

AND2x2_ASAP7_75t_L g6883 ( 
.A(n_6780),
.B(n_1796),
.Y(n_6883)
);

OAI222xp33_ASAP7_75t_L g6884 ( 
.A1(n_6778),
.A2(n_1026),
.B1(n_1028),
.B2(n_1024),
.C1(n_1025),
.C2(n_1027),
.Y(n_6884)
);

OR2x2_ASAP7_75t_L g6885 ( 
.A(n_6777),
.B(n_1024),
.Y(n_6885)
);

HB1xp67_ASAP7_75t_L g6886 ( 
.A(n_6718),
.Y(n_6886)
);

INVxp67_ASAP7_75t_L g6887 ( 
.A(n_6763),
.Y(n_6887)
);

NAND2xp33_ASAP7_75t_SL g6888 ( 
.A(n_6735),
.B(n_1025),
.Y(n_6888)
);

INVx1_ASAP7_75t_SL g6889 ( 
.A(n_6733),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6781),
.Y(n_6890)
);

INVx1_ASAP7_75t_SL g6891 ( 
.A(n_6792),
.Y(n_6891)
);

OR2x2_ASAP7_75t_L g6892 ( 
.A(n_6741),
.B(n_1026),
.Y(n_6892)
);

NAND2xp5_ASAP7_75t_L g6893 ( 
.A(n_6745),
.B(n_1027),
.Y(n_6893)
);

NAND2xp5_ASAP7_75t_L g6894 ( 
.A(n_6773),
.B(n_1028),
.Y(n_6894)
);

INVx1_ASAP7_75t_L g6895 ( 
.A(n_6774),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6767),
.B(n_1029),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_L g6897 ( 
.A(n_6716),
.B(n_1029),
.Y(n_6897)
);

INVx1_ASAP7_75t_L g6898 ( 
.A(n_6760),
.Y(n_6898)
);

INVxp67_ASAP7_75t_L g6899 ( 
.A(n_6736),
.Y(n_6899)
);

NAND2xp5_ASAP7_75t_L g6900 ( 
.A(n_6798),
.B(n_1030),
.Y(n_6900)
);

NOR3xp33_ASAP7_75t_SL g6901 ( 
.A(n_6856),
.B(n_1031),
.C(n_1032),
.Y(n_6901)
);

AOI22xp5_ASAP7_75t_L g6902 ( 
.A1(n_6803),
.A2(n_1036),
.B1(n_1033),
.B2(n_1034),
.Y(n_6902)
);

NOR2x1_ASAP7_75t_L g6903 ( 
.A(n_6806),
.B(n_1033),
.Y(n_6903)
);

NAND2xp5_ASAP7_75t_L g6904 ( 
.A(n_6821),
.B(n_1037),
.Y(n_6904)
);

HB1xp67_ASAP7_75t_L g6905 ( 
.A(n_6825),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_6814),
.Y(n_6906)
);

NOR2xp33_ASAP7_75t_L g6907 ( 
.A(n_6891),
.B(n_1034),
.Y(n_6907)
);

NAND4xp25_ASAP7_75t_SL g6908 ( 
.A(n_6881),
.B(n_1042),
.C(n_1038),
.D(n_1039),
.Y(n_6908)
);

AOI21xp5_ASAP7_75t_L g6909 ( 
.A1(n_6807),
.A2(n_1039),
.B(n_1042),
.Y(n_6909)
);

INVx1_ASAP7_75t_L g6910 ( 
.A(n_6816),
.Y(n_6910)
);

NAND4xp25_ASAP7_75t_L g6911 ( 
.A(n_6869),
.B(n_1045),
.C(n_1043),
.D(n_1044),
.Y(n_6911)
);

NAND2xp5_ASAP7_75t_L g6912 ( 
.A(n_6802),
.B(n_1044),
.Y(n_6912)
);

INVx1_ASAP7_75t_L g6913 ( 
.A(n_6846),
.Y(n_6913)
);

NOR4xp25_ASAP7_75t_L g6914 ( 
.A(n_6819),
.B(n_1046),
.C(n_1043),
.D(n_1045),
.Y(n_6914)
);

NOR2xp33_ASAP7_75t_SL g6915 ( 
.A(n_6827),
.B(n_1047),
.Y(n_6915)
);

AOI221xp5_ASAP7_75t_L g6916 ( 
.A1(n_6828),
.A2(n_1050),
.B1(n_1048),
.B2(n_1049),
.C(n_1051),
.Y(n_6916)
);

OAI21xp5_ASAP7_75t_L g6917 ( 
.A1(n_6812),
.A2(n_1048),
.B(n_1050),
.Y(n_6917)
);

NOR2xp33_ASAP7_75t_L g6918 ( 
.A(n_6830),
.B(n_1051),
.Y(n_6918)
);

NAND2xp5_ASAP7_75t_L g6919 ( 
.A(n_6805),
.B(n_1053),
.Y(n_6919)
);

OAI21xp33_ASAP7_75t_L g6920 ( 
.A1(n_6874),
.A2(n_6824),
.B(n_6817),
.Y(n_6920)
);

NAND2xp5_ASAP7_75t_L g6921 ( 
.A(n_6835),
.B(n_1054),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6826),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6829),
.Y(n_6923)
);

INVx1_ASAP7_75t_L g6924 ( 
.A(n_6829),
.Y(n_6924)
);

AOI211xp5_ASAP7_75t_L g6925 ( 
.A1(n_6810),
.A2(n_1055),
.B(n_1052),
.C(n_1054),
.Y(n_6925)
);

NAND2xp5_ASAP7_75t_L g6926 ( 
.A(n_6836),
.B(n_1055),
.Y(n_6926)
);

AOI211xp5_ASAP7_75t_L g6927 ( 
.A1(n_6844),
.A2(n_1058),
.B(n_1052),
.C(n_1057),
.Y(n_6927)
);

NAND2x1_ASAP7_75t_SL g6928 ( 
.A(n_6811),
.B(n_1057),
.Y(n_6928)
);

NAND2xp5_ASAP7_75t_SL g6929 ( 
.A(n_6808),
.B(n_1058),
.Y(n_6929)
);

NOR4xp25_ASAP7_75t_L g6930 ( 
.A(n_6880),
.B(n_6839),
.C(n_6840),
.D(n_6864),
.Y(n_6930)
);

INVx1_ASAP7_75t_L g6931 ( 
.A(n_6820),
.Y(n_6931)
);

NAND3xp33_ASAP7_75t_L g6932 ( 
.A(n_6870),
.B(n_1059),
.C(n_1060),
.Y(n_6932)
);

NOR4xp25_ASAP7_75t_L g6933 ( 
.A(n_6855),
.B(n_1063),
.C(n_1059),
.D(n_1062),
.Y(n_6933)
);

AOI22xp5_ASAP7_75t_L g6934 ( 
.A1(n_6866),
.A2(n_1065),
.B1(n_1063),
.B2(n_1064),
.Y(n_6934)
);

NOR3xp33_ASAP7_75t_L g6935 ( 
.A(n_6804),
.B(n_1064),
.C(n_1065),
.Y(n_6935)
);

AOI32xp33_ASAP7_75t_L g6936 ( 
.A1(n_6849),
.A2(n_6834),
.A3(n_6888),
.B1(n_6879),
.B2(n_6875),
.Y(n_6936)
);

INVx1_ASAP7_75t_L g6937 ( 
.A(n_6842),
.Y(n_6937)
);

NAND2xp5_ASAP7_75t_L g6938 ( 
.A(n_6831),
.B(n_1067),
.Y(n_6938)
);

NAND2xp5_ASAP7_75t_L g6939 ( 
.A(n_6860),
.B(n_1067),
.Y(n_6939)
);

NAND3xp33_ASAP7_75t_SL g6940 ( 
.A(n_6877),
.B(n_1066),
.C(n_1068),
.Y(n_6940)
);

NAND2xp5_ASAP7_75t_L g6941 ( 
.A(n_6837),
.B(n_1068),
.Y(n_6941)
);

NAND3xp33_ASAP7_75t_L g6942 ( 
.A(n_6878),
.B(n_1066),
.C(n_1069),
.Y(n_6942)
);

NOR2xp33_ASAP7_75t_L g6943 ( 
.A(n_6884),
.B(n_1070),
.Y(n_6943)
);

AOI211xp5_ASAP7_75t_SL g6944 ( 
.A1(n_6900),
.A2(n_6853),
.B(n_6815),
.C(n_6852),
.Y(n_6944)
);

INVx1_ASAP7_75t_L g6945 ( 
.A(n_6818),
.Y(n_6945)
);

NAND3xp33_ASAP7_75t_L g6946 ( 
.A(n_6822),
.B(n_1070),
.C(n_1071),
.Y(n_6946)
);

NOR3x1_ASAP7_75t_L g6947 ( 
.A(n_6843),
.B(n_1079),
.C(n_1071),
.Y(n_6947)
);

AOI211x1_ASAP7_75t_SL g6948 ( 
.A1(n_6851),
.A2(n_1074),
.B(n_1072),
.C(n_1073),
.Y(n_6948)
);

NOR2xp33_ASAP7_75t_L g6949 ( 
.A(n_6809),
.B(n_6833),
.Y(n_6949)
);

INVx1_ASAP7_75t_L g6950 ( 
.A(n_6883),
.Y(n_6950)
);

NAND3xp33_ASAP7_75t_L g6951 ( 
.A(n_6858),
.B(n_1073),
.C(n_1074),
.Y(n_6951)
);

NOR2xp33_ASAP7_75t_L g6952 ( 
.A(n_6848),
.B(n_1075),
.Y(n_6952)
);

NAND4xp25_ASAP7_75t_L g6953 ( 
.A(n_6882),
.B(n_1077),
.C(n_1075),
.D(n_1076),
.Y(n_6953)
);

NOR2x1_ASAP7_75t_L g6954 ( 
.A(n_6838),
.B(n_1076),
.Y(n_6954)
);

NAND3xp33_ASAP7_75t_SL g6955 ( 
.A(n_6859),
.B(n_1078),
.C(n_1080),
.Y(n_6955)
);

INVx1_ASAP7_75t_L g6956 ( 
.A(n_6876),
.Y(n_6956)
);

AOI22xp5_ASAP7_75t_L g6957 ( 
.A1(n_6861),
.A2(n_1083),
.B1(n_1081),
.B2(n_1082),
.Y(n_6957)
);

AOI221xp5_ASAP7_75t_L g6958 ( 
.A1(n_6857),
.A2(n_1083),
.B1(n_1081),
.B2(n_1082),
.C(n_1084),
.Y(n_6958)
);

NAND4xp25_ASAP7_75t_L g6959 ( 
.A(n_6889),
.B(n_1088),
.C(n_1086),
.D(n_1087),
.Y(n_6959)
);

AND4x1_ASAP7_75t_L g6960 ( 
.A(n_6845),
.B(n_1089),
.C(n_1086),
.D(n_1087),
.Y(n_6960)
);

NAND2xp5_ASAP7_75t_L g6961 ( 
.A(n_6850),
.B(n_1090),
.Y(n_6961)
);

AOI32xp33_ASAP7_75t_L g6962 ( 
.A1(n_6895),
.A2(n_1092),
.A3(n_1089),
.B1(n_1091),
.B2(n_1095),
.Y(n_6962)
);

NOR2xp33_ASAP7_75t_L g6963 ( 
.A(n_6867),
.B(n_1095),
.Y(n_6963)
);

INVx1_ASAP7_75t_L g6964 ( 
.A(n_6886),
.Y(n_6964)
);

NOR3x1_ASAP7_75t_L g6965 ( 
.A(n_6873),
.B(n_1105),
.C(n_1097),
.Y(n_6965)
);

AOI221x1_ASAP7_75t_L g6966 ( 
.A1(n_6854),
.A2(n_1099),
.B1(n_1097),
.B2(n_1098),
.C(n_1100),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6865),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6868),
.B(n_1101),
.Y(n_6968)
);

A2O1A1Ixp33_ASAP7_75t_L g6969 ( 
.A1(n_6885),
.A2(n_1102),
.B(n_1098),
.C(n_1101),
.Y(n_6969)
);

INVx1_ASAP7_75t_L g6970 ( 
.A(n_6896),
.Y(n_6970)
);

AOI21xp5_ASAP7_75t_L g6971 ( 
.A1(n_6897),
.A2(n_6863),
.B(n_6847),
.Y(n_6971)
);

OAI21xp33_ASAP7_75t_L g6972 ( 
.A1(n_6898),
.A2(n_1102),
.B(n_1103),
.Y(n_6972)
);

INVx1_ASAP7_75t_L g6973 ( 
.A(n_6832),
.Y(n_6973)
);

AOI21xp5_ASAP7_75t_L g6974 ( 
.A1(n_6801),
.A2(n_1104),
.B(n_1107),
.Y(n_6974)
);

INVxp67_ASAP7_75t_L g6975 ( 
.A(n_6872),
.Y(n_6975)
);

INVx1_ASAP7_75t_L g6976 ( 
.A(n_6841),
.Y(n_6976)
);

NOR2xp33_ASAP7_75t_SL g6977 ( 
.A(n_6899),
.B(n_1107),
.Y(n_6977)
);

NAND2xp5_ASAP7_75t_SL g6978 ( 
.A(n_6823),
.B(n_1108),
.Y(n_6978)
);

NOR2xp33_ASAP7_75t_L g6979 ( 
.A(n_6862),
.B(n_1108),
.Y(n_6979)
);

NAND2xp5_ASAP7_75t_L g6980 ( 
.A(n_6813),
.B(n_1110),
.Y(n_6980)
);

AOI21xp5_ASAP7_75t_L g6981 ( 
.A1(n_6894),
.A2(n_1109),
.B(n_1110),
.Y(n_6981)
);

NOR4xp25_ASAP7_75t_L g6982 ( 
.A(n_6887),
.B(n_6890),
.C(n_6893),
.D(n_6892),
.Y(n_6982)
);

INVx1_ASAP7_75t_L g6983 ( 
.A(n_6871),
.Y(n_6983)
);

NAND4xp25_ASAP7_75t_L g6984 ( 
.A(n_6869),
.B(n_1112),
.C(n_1109),
.D(n_1111),
.Y(n_6984)
);

AOI22xp5_ASAP7_75t_L g6985 ( 
.A1(n_6803),
.A2(n_1113),
.B1(n_1111),
.B2(n_1112),
.Y(n_6985)
);

AOI221xp5_ASAP7_75t_L g6986 ( 
.A1(n_6803),
.A2(n_1116),
.B1(n_1114),
.B2(n_1115),
.C(n_1117),
.Y(n_6986)
);

AOI21xp5_ASAP7_75t_L g6987 ( 
.A1(n_6821),
.A2(n_1114),
.B(n_1115),
.Y(n_6987)
);

AOI22xp5_ASAP7_75t_L g6988 ( 
.A1(n_6803),
.A2(n_1118),
.B1(n_1116),
.B2(n_1117),
.Y(n_6988)
);

NAND3xp33_ASAP7_75t_L g6989 ( 
.A(n_6803),
.B(n_1119),
.C(n_1120),
.Y(n_6989)
);

NAND2xp5_ASAP7_75t_L g6990 ( 
.A(n_6821),
.B(n_1122),
.Y(n_6990)
);

NAND4xp25_ASAP7_75t_L g6991 ( 
.A(n_6869),
.B(n_1124),
.C(n_1121),
.D(n_1123),
.Y(n_6991)
);

O2A1O1Ixp5_ASAP7_75t_L g6992 ( 
.A1(n_6824),
.A2(n_1125),
.B(n_1121),
.C(n_1123),
.Y(n_6992)
);

NAND2xp5_ASAP7_75t_L g6993 ( 
.A(n_6821),
.B(n_1126),
.Y(n_6993)
);

NOR3xp33_ASAP7_75t_L g6994 ( 
.A(n_6803),
.B(n_1125),
.C(n_1126),
.Y(n_6994)
);

NAND4xp25_ASAP7_75t_SL g6995 ( 
.A(n_6856),
.B(n_1130),
.C(n_1127),
.D(n_1128),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6821),
.Y(n_6996)
);

AOI221x1_ASAP7_75t_L g6997 ( 
.A1(n_6856),
.A2(n_1133),
.B1(n_1128),
.B2(n_1131),
.C(n_1134),
.Y(n_6997)
);

AOI211xp5_ASAP7_75t_SL g6998 ( 
.A1(n_6803),
.A2(n_1134),
.B(n_1131),
.C(n_1133),
.Y(n_6998)
);

OAI211xp5_ASAP7_75t_L g6999 ( 
.A1(n_6803),
.A2(n_1137),
.B(n_1135),
.C(n_1136),
.Y(n_6999)
);

INVx1_ASAP7_75t_L g7000 ( 
.A(n_6905),
.Y(n_7000)
);

AND2x2_ASAP7_75t_L g7001 ( 
.A(n_6996),
.B(n_1135),
.Y(n_7001)
);

AOI211xp5_ASAP7_75t_L g7002 ( 
.A1(n_6906),
.A2(n_6995),
.B(n_6930),
.C(n_6920),
.Y(n_7002)
);

NAND3xp33_ASAP7_75t_L g7003 ( 
.A(n_6901),
.B(n_1136),
.C(n_1138),
.Y(n_7003)
);

INVx1_ASAP7_75t_L g7004 ( 
.A(n_6928),
.Y(n_7004)
);

NOR2xp33_ASAP7_75t_L g7005 ( 
.A(n_6923),
.B(n_1138),
.Y(n_7005)
);

O2A1O1Ixp33_ASAP7_75t_L g7006 ( 
.A1(n_6975),
.A2(n_1141),
.B(n_1139),
.C(n_1140),
.Y(n_7006)
);

NAND5xp2_ASAP7_75t_L g7007 ( 
.A(n_6944),
.B(n_1141),
.C(n_1139),
.D(n_1140),
.E(n_1142),
.Y(n_7007)
);

AND2x2_ASAP7_75t_L g7008 ( 
.A(n_6964),
.B(n_1143),
.Y(n_7008)
);

INVx2_ASAP7_75t_L g7009 ( 
.A(n_6903),
.Y(n_7009)
);

OA22x2_ASAP7_75t_L g7010 ( 
.A1(n_6997),
.A2(n_1145),
.B1(n_1143),
.B2(n_1144),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6926),
.Y(n_7011)
);

NOR2xp67_ASAP7_75t_L g7012 ( 
.A(n_6908),
.B(n_1145),
.Y(n_7012)
);

NAND2xp5_ASAP7_75t_L g7013 ( 
.A(n_6948),
.B(n_1146),
.Y(n_7013)
);

NOR3xp33_ASAP7_75t_L g7014 ( 
.A(n_6924),
.B(n_1795),
.C(n_1793),
.Y(n_7014)
);

INVx1_ASAP7_75t_L g7015 ( 
.A(n_6954),
.Y(n_7015)
);

AOI22xp5_ASAP7_75t_L g7016 ( 
.A1(n_6949),
.A2(n_1149),
.B1(n_1146),
.B2(n_1148),
.Y(n_7016)
);

NOR2xp33_ASAP7_75t_L g7017 ( 
.A(n_6915),
.B(n_1149),
.Y(n_7017)
);

NAND3xp33_ASAP7_75t_L g7018 ( 
.A(n_6977),
.B(n_1150),
.C(n_1151),
.Y(n_7018)
);

AOI221xp5_ASAP7_75t_L g7019 ( 
.A1(n_6907),
.A2(n_1153),
.B1(n_1151),
.B2(n_1152),
.C(n_1155),
.Y(n_7019)
);

NOR2xp33_ASAP7_75t_L g7020 ( 
.A(n_6911),
.B(n_1153),
.Y(n_7020)
);

OR2x2_ASAP7_75t_L g7021 ( 
.A(n_6914),
.B(n_1155),
.Y(n_7021)
);

NOR2x1_ASAP7_75t_L g7022 ( 
.A(n_6904),
.B(n_1156),
.Y(n_7022)
);

OR2x2_ASAP7_75t_L g7023 ( 
.A(n_6933),
.B(n_1156),
.Y(n_7023)
);

XOR2x2_ASAP7_75t_L g7024 ( 
.A(n_6960),
.B(n_1158),
.Y(n_7024)
);

AOI22xp5_ASAP7_75t_L g7025 ( 
.A1(n_6970),
.A2(n_1159),
.B1(n_1157),
.B2(n_1158),
.Y(n_7025)
);

NAND4xp25_ASAP7_75t_L g7026 ( 
.A(n_6965),
.B(n_1160),
.C(n_1157),
.D(n_1159),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6961),
.Y(n_7027)
);

AND2x2_ASAP7_75t_L g7028 ( 
.A(n_6922),
.B(n_1161),
.Y(n_7028)
);

NAND3xp33_ASAP7_75t_L g7029 ( 
.A(n_6998),
.B(n_1161),
.C(n_1162),
.Y(n_7029)
);

NAND2xp5_ASAP7_75t_L g7030 ( 
.A(n_6966),
.B(n_1162),
.Y(n_7030)
);

AND4x1_ASAP7_75t_L g7031 ( 
.A(n_6918),
.B(n_1165),
.C(n_1163),
.D(n_1164),
.Y(n_7031)
);

OAI22xp5_ASAP7_75t_L g7032 ( 
.A1(n_6990),
.A2(n_1168),
.B1(n_1165),
.B2(n_1166),
.Y(n_7032)
);

NAND2xp5_ASAP7_75t_SL g7033 ( 
.A(n_6925),
.B(n_1166),
.Y(n_7033)
);

AOI22xp5_ASAP7_75t_L g7034 ( 
.A1(n_6912),
.A2(n_1170),
.B1(n_1168),
.B2(n_1169),
.Y(n_7034)
);

OAI211xp5_ASAP7_75t_L g7035 ( 
.A1(n_6962),
.A2(n_1172),
.B(n_1169),
.C(n_1171),
.Y(n_7035)
);

NOR2xp33_ASAP7_75t_SL g7036 ( 
.A(n_6984),
.B(n_1173),
.Y(n_7036)
);

NOR2x1_ASAP7_75t_L g7037 ( 
.A(n_6993),
.B(n_1173),
.Y(n_7037)
);

NOR2xp33_ASAP7_75t_L g7038 ( 
.A(n_6991),
.B(n_6959),
.Y(n_7038)
);

NOR2xp33_ASAP7_75t_L g7039 ( 
.A(n_6940),
.B(n_6999),
.Y(n_7039)
);

NOR2x1_ASAP7_75t_L g7040 ( 
.A(n_6989),
.B(n_1174),
.Y(n_7040)
);

INVxp67_ASAP7_75t_L g7041 ( 
.A(n_6943),
.Y(n_7041)
);

INVx1_ASAP7_75t_L g7042 ( 
.A(n_6941),
.Y(n_7042)
);

AND2x2_ASAP7_75t_L g7043 ( 
.A(n_6910),
.B(n_1174),
.Y(n_7043)
);

NAND2xp5_ASAP7_75t_L g7044 ( 
.A(n_6952),
.B(n_1175),
.Y(n_7044)
);

NOR2xp33_ASAP7_75t_L g7045 ( 
.A(n_6955),
.B(n_1175),
.Y(n_7045)
);

NOR4xp25_ASAP7_75t_L g7046 ( 
.A(n_6917),
.B(n_1179),
.C(n_1176),
.D(n_1178),
.Y(n_7046)
);

NOR3xp33_ASAP7_75t_SL g7047 ( 
.A(n_6942),
.B(n_1179),
.C(n_1181),
.Y(n_7047)
);

OAI21xp5_ASAP7_75t_SL g7048 ( 
.A1(n_6987),
.A2(n_1181),
.B(n_1182),
.Y(n_7048)
);

OAI21x1_ASAP7_75t_L g7049 ( 
.A1(n_6992),
.A2(n_6909),
.B(n_6981),
.Y(n_7049)
);

AOI22xp5_ASAP7_75t_L g7050 ( 
.A1(n_6919),
.A2(n_1186),
.B1(n_1184),
.B2(n_1185),
.Y(n_7050)
);

NOR3xp33_ASAP7_75t_SL g7051 ( 
.A(n_6971),
.B(n_1184),
.C(n_1185),
.Y(n_7051)
);

HAxp5_ASAP7_75t_SL g7052 ( 
.A(n_6937),
.B(n_1186),
.CON(n_7052),
.SN(n_7052)
);

NOR2xp33_ASAP7_75t_L g7053 ( 
.A(n_6953),
.B(n_1187),
.Y(n_7053)
);

NOR2xp33_ASAP7_75t_L g7054 ( 
.A(n_6939),
.B(n_1187),
.Y(n_7054)
);

AOI22xp33_ASAP7_75t_L g7055 ( 
.A1(n_6945),
.A2(n_1190),
.B1(n_1188),
.B2(n_1189),
.Y(n_7055)
);

INVx1_ASAP7_75t_L g7056 ( 
.A(n_6931),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_6947),
.Y(n_7057)
);

NOR2xp33_ASAP7_75t_R g7058 ( 
.A(n_6921),
.B(n_1188),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_6968),
.Y(n_7059)
);

INVx1_ASAP7_75t_L g7060 ( 
.A(n_6913),
.Y(n_7060)
);

AOI22xp5_ASAP7_75t_L g7061 ( 
.A1(n_6963),
.A2(n_1194),
.B1(n_1191),
.B2(n_1193),
.Y(n_7061)
);

AOI22xp5_ASAP7_75t_L g7062 ( 
.A1(n_6967),
.A2(n_1195),
.B1(n_1193),
.B2(n_1194),
.Y(n_7062)
);

NOR2x1_ASAP7_75t_L g7063 ( 
.A(n_6938),
.B(n_1195),
.Y(n_7063)
);

INVxp67_ASAP7_75t_L g7064 ( 
.A(n_6979),
.Y(n_7064)
);

INVxp67_ASAP7_75t_SL g7065 ( 
.A(n_6927),
.Y(n_7065)
);

INVx1_ASAP7_75t_L g7066 ( 
.A(n_6950),
.Y(n_7066)
);

INVx1_ASAP7_75t_L g7067 ( 
.A(n_6956),
.Y(n_7067)
);

AOI21xp5_ASAP7_75t_L g7068 ( 
.A1(n_6916),
.A2(n_1197),
.B(n_1198),
.Y(n_7068)
);

NAND2xp5_ASAP7_75t_L g7069 ( 
.A(n_6935),
.B(n_1197),
.Y(n_7069)
);

NOR2xp33_ASAP7_75t_L g7070 ( 
.A(n_6929),
.B(n_1198),
.Y(n_7070)
);

NOR2xp33_ASAP7_75t_SL g7071 ( 
.A(n_6972),
.B(n_1199),
.Y(n_7071)
);

NAND3xp33_ASAP7_75t_L g7072 ( 
.A(n_6936),
.B(n_1199),
.C(n_1200),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6932),
.Y(n_7073)
);

NOR2xp33_ASAP7_75t_L g7074 ( 
.A(n_6973),
.B(n_1200),
.Y(n_7074)
);

NAND4xp25_ASAP7_75t_L g7075 ( 
.A(n_6974),
.B(n_1204),
.C(n_1201),
.D(n_1203),
.Y(n_7075)
);

NAND2xp33_ASAP7_75t_SL g7076 ( 
.A(n_6980),
.B(n_1203),
.Y(n_7076)
);

OAI221xp5_ASAP7_75t_L g7077 ( 
.A1(n_6994),
.A2(n_1206),
.B1(n_1201),
.B2(n_1205),
.C(n_1207),
.Y(n_7077)
);

NAND2xp5_ASAP7_75t_SL g7078 ( 
.A(n_6986),
.B(n_1205),
.Y(n_7078)
);

NAND3xp33_ASAP7_75t_L g7079 ( 
.A(n_6969),
.B(n_6976),
.C(n_6946),
.Y(n_7079)
);

AOI221xp5_ASAP7_75t_L g7080 ( 
.A1(n_6982),
.A2(n_1209),
.B1(n_1207),
.B2(n_1208),
.C(n_1210),
.Y(n_7080)
);

NOR3x1_ASAP7_75t_L g7081 ( 
.A(n_6951),
.B(n_1208),
.C(n_1209),
.Y(n_7081)
);

NOR2x1_ASAP7_75t_L g7082 ( 
.A(n_6983),
.B(n_1210),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6957),
.Y(n_7083)
);

NAND2xp5_ASAP7_75t_L g7084 ( 
.A(n_6902),
.B(n_1211),
.Y(n_7084)
);

AOI221xp5_ASAP7_75t_SL g7085 ( 
.A1(n_6978),
.A2(n_1213),
.B1(n_1211),
.B2(n_1212),
.C(n_1215),
.Y(n_7085)
);

NOR2xp67_ASAP7_75t_L g7086 ( 
.A(n_6985),
.B(n_1216),
.Y(n_7086)
);

NAND3xp33_ASAP7_75t_L g7087 ( 
.A(n_6988),
.B(n_1216),
.C(n_1217),
.Y(n_7087)
);

OAI21xp5_ASAP7_75t_L g7088 ( 
.A1(n_6934),
.A2(n_6958),
.B(n_1217),
.Y(n_7088)
);

HB1xp67_ASAP7_75t_L g7089 ( 
.A(n_6905),
.Y(n_7089)
);

NAND2xp5_ASAP7_75t_L g7090 ( 
.A(n_6905),
.B(n_1218),
.Y(n_7090)
);

AOI21xp5_ASAP7_75t_L g7091 ( 
.A1(n_6905),
.A2(n_1218),
.B(n_1219),
.Y(n_7091)
);

O2A1O1Ixp5_ASAP7_75t_SL g7092 ( 
.A1(n_6905),
.A2(n_1225),
.B(n_1222),
.C(n_1224),
.Y(n_7092)
);

NAND2xp5_ASAP7_75t_L g7093 ( 
.A(n_6905),
.B(n_1222),
.Y(n_7093)
);

INVx1_ASAP7_75t_SL g7094 ( 
.A(n_6905),
.Y(n_7094)
);

NAND2xp5_ASAP7_75t_L g7095 ( 
.A(n_7089),
.B(n_7094),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_7000),
.B(n_1224),
.Y(n_7096)
);

INVx2_ASAP7_75t_SL g7097 ( 
.A(n_7024),
.Y(n_7097)
);

AOI21xp5_ASAP7_75t_L g7098 ( 
.A1(n_7090),
.A2(n_1225),
.B(n_1226),
.Y(n_7098)
);

NAND2xp5_ASAP7_75t_L g7099 ( 
.A(n_7004),
.B(n_1226),
.Y(n_7099)
);

NOR2x1_ASAP7_75t_L g7100 ( 
.A(n_7093),
.B(n_1227),
.Y(n_7100)
);

NAND5xp2_ASAP7_75t_L g7101 ( 
.A(n_7002),
.B(n_1231),
.C(n_1229),
.D(n_1230),
.E(n_1233),
.Y(n_7101)
);

NAND2xp5_ASAP7_75t_L g7102 ( 
.A(n_7057),
.B(n_1230),
.Y(n_7102)
);

INVx1_ASAP7_75t_L g7103 ( 
.A(n_7010),
.Y(n_7103)
);

INVx1_ASAP7_75t_L g7104 ( 
.A(n_7023),
.Y(n_7104)
);

NOR2xp33_ASAP7_75t_L g7105 ( 
.A(n_7007),
.B(n_1233),
.Y(n_7105)
);

NAND4xp25_ASAP7_75t_L g7106 ( 
.A(n_7003),
.B(n_1237),
.C(n_1235),
.D(n_1236),
.Y(n_7106)
);

OAI221xp5_ASAP7_75t_L g7107 ( 
.A1(n_7048),
.A2(n_1238),
.B1(n_1235),
.B2(n_1236),
.C(n_1239),
.Y(n_7107)
);

AOI211xp5_ASAP7_75t_L g7108 ( 
.A1(n_7080),
.A2(n_1241),
.B(n_1238),
.C(n_1240),
.Y(n_7108)
);

AOI211xp5_ASAP7_75t_L g7109 ( 
.A1(n_7013),
.A2(n_1244),
.B(n_1242),
.C(n_1243),
.Y(n_7109)
);

INVxp67_ASAP7_75t_L g7110 ( 
.A(n_7021),
.Y(n_7110)
);

AND3x1_ASAP7_75t_L g7111 ( 
.A(n_7051),
.B(n_1251),
.C(n_1242),
.Y(n_7111)
);

AOI21xp5_ASAP7_75t_L g7112 ( 
.A1(n_7006),
.A2(n_1243),
.B(n_1245),
.Y(n_7112)
);

OAI211xp5_ASAP7_75t_SL g7113 ( 
.A1(n_7041),
.A2(n_1248),
.B(n_1246),
.C(n_1247),
.Y(n_7113)
);

NAND3xp33_ASAP7_75t_L g7114 ( 
.A(n_7052),
.B(n_1247),
.C(n_1249),
.Y(n_7114)
);

OAI211xp5_ASAP7_75t_L g7115 ( 
.A1(n_7091),
.A2(n_1252),
.B(n_1249),
.C(n_1250),
.Y(n_7115)
);

OAI221xp5_ASAP7_75t_L g7116 ( 
.A1(n_7066),
.A2(n_1253),
.B1(n_1250),
.B2(n_1252),
.C(n_1254),
.Y(n_7116)
);

NOR2x1p5_ASAP7_75t_L g7117 ( 
.A(n_7029),
.B(n_1253),
.Y(n_7117)
);

AND2x2_ASAP7_75t_L g7118 ( 
.A(n_7008),
.B(n_1254),
.Y(n_7118)
);

AOI21x1_ASAP7_75t_L g7119 ( 
.A1(n_7001),
.A2(n_7028),
.B(n_7067),
.Y(n_7119)
);

AND2x2_ASAP7_75t_L g7120 ( 
.A(n_7043),
.B(n_1256),
.Y(n_7120)
);

NOR2xp33_ASAP7_75t_L g7121 ( 
.A(n_7026),
.B(n_7030),
.Y(n_7121)
);

NOR2x1_ASAP7_75t_SL g7122 ( 
.A(n_7035),
.B(n_1257),
.Y(n_7122)
);

INVx1_ASAP7_75t_L g7123 ( 
.A(n_7022),
.Y(n_7123)
);

NAND3xp33_ASAP7_75t_L g7124 ( 
.A(n_7015),
.B(n_1258),
.C(n_1259),
.Y(n_7124)
);

NAND4xp25_ASAP7_75t_SL g7125 ( 
.A(n_7085),
.B(n_1260),
.C(n_1258),
.D(n_1259),
.Y(n_7125)
);

INVxp33_ASAP7_75t_L g7126 ( 
.A(n_7058),
.Y(n_7126)
);

NOR3xp33_ASAP7_75t_L g7127 ( 
.A(n_7056),
.B(n_1261),
.C(n_1262),
.Y(n_7127)
);

AOI221xp5_ASAP7_75t_L g7128 ( 
.A1(n_7060),
.A2(n_1264),
.B1(n_1262),
.B2(n_1263),
.C(n_1265),
.Y(n_7128)
);

OR2x2_ASAP7_75t_L g7129 ( 
.A(n_7046),
.B(n_1263),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_7009),
.Y(n_7130)
);

NOR2xp33_ASAP7_75t_L g7131 ( 
.A(n_7031),
.B(n_1264),
.Y(n_7131)
);

OAI211xp5_ASAP7_75t_L g7132 ( 
.A1(n_7020),
.A2(n_1268),
.B(n_1265),
.C(n_1266),
.Y(n_7132)
);

NOR3xp33_ASAP7_75t_SL g7133 ( 
.A(n_7079),
.B(n_1266),
.C(n_1268),
.Y(n_7133)
);

NOR2xp33_ASAP7_75t_L g7134 ( 
.A(n_7036),
.B(n_1269),
.Y(n_7134)
);

NOR3xp33_ASAP7_75t_L g7135 ( 
.A(n_7011),
.B(n_1270),
.C(n_1271),
.Y(n_7135)
);

NAND4xp25_ASAP7_75t_SL g7136 ( 
.A(n_7072),
.B(n_1272),
.C(n_1270),
.D(n_1271),
.Y(n_7136)
);

AOI211xp5_ASAP7_75t_SL g7137 ( 
.A1(n_7012),
.A2(n_1274),
.B(n_1272),
.C(n_1273),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_7037),
.Y(n_7138)
);

NAND3xp33_ASAP7_75t_L g7139 ( 
.A(n_7082),
.B(n_1273),
.C(n_1275),
.Y(n_7139)
);

NAND2xp33_ASAP7_75t_SL g7140 ( 
.A(n_7047),
.B(n_1275),
.Y(n_7140)
);

NOR2xp33_ASAP7_75t_L g7141 ( 
.A(n_7075),
.B(n_1276),
.Y(n_7141)
);

NAND4xp25_ASAP7_75t_L g7142 ( 
.A(n_7081),
.B(n_1278),
.C(n_1276),
.D(n_1277),
.Y(n_7142)
);

NOR2x1_ASAP7_75t_SL g7143 ( 
.A(n_7032),
.B(n_1277),
.Y(n_7143)
);

XNOR2xp5_ASAP7_75t_L g7144 ( 
.A(n_7063),
.B(n_1278),
.Y(n_7144)
);

NAND3xp33_ASAP7_75t_SL g7145 ( 
.A(n_7092),
.B(n_1288),
.C(n_1279),
.Y(n_7145)
);

NAND4xp75_ASAP7_75t_L g7146 ( 
.A(n_7040),
.B(n_1282),
.C(n_1280),
.D(n_1281),
.Y(n_7146)
);

NOR2xp33_ASAP7_75t_L g7147 ( 
.A(n_7018),
.B(n_1283),
.Y(n_7147)
);

OAI222xp33_ASAP7_75t_L g7148 ( 
.A1(n_7033),
.A2(n_1285),
.B1(n_1288),
.B2(n_1283),
.C1(n_1284),
.C2(n_1287),
.Y(n_7148)
);

INVx1_ASAP7_75t_L g7149 ( 
.A(n_7049),
.Y(n_7149)
);

OAI21xp5_ASAP7_75t_L g7150 ( 
.A1(n_7038),
.A2(n_1285),
.B(n_1287),
.Y(n_7150)
);

INVx1_ASAP7_75t_L g7151 ( 
.A(n_7044),
.Y(n_7151)
);

OAI211xp5_ASAP7_75t_L g7152 ( 
.A1(n_7065),
.A2(n_1291),
.B(n_1289),
.C(n_1290),
.Y(n_7152)
);

A2O1A1Ixp33_ASAP7_75t_L g7153 ( 
.A1(n_7054),
.A2(n_1291),
.B(n_1289),
.C(n_1290),
.Y(n_7153)
);

NAND3xp33_ASAP7_75t_L g7154 ( 
.A(n_7074),
.B(n_1292),
.C(n_1293),
.Y(n_7154)
);

AOI21xp5_ASAP7_75t_L g7155 ( 
.A1(n_7078),
.A2(n_1292),
.B(n_1293),
.Y(n_7155)
);

AND4x1_ASAP7_75t_L g7156 ( 
.A(n_7053),
.B(n_1297),
.C(n_1294),
.D(n_1296),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_L g7157 ( 
.A(n_7017),
.B(n_1296),
.Y(n_7157)
);

NAND4xp25_ASAP7_75t_SL g7158 ( 
.A(n_7068),
.B(n_1300),
.C(n_1298),
.D(n_1299),
.Y(n_7158)
);

AOI32xp33_ASAP7_75t_L g7159 ( 
.A1(n_7071),
.A2(n_1300),
.A3(n_1298),
.B1(n_1299),
.B2(n_1301),
.Y(n_7159)
);

NOR4xp25_ASAP7_75t_L g7160 ( 
.A(n_7064),
.B(n_7073),
.C(n_7059),
.D(n_7027),
.Y(n_7160)
);

NAND4xp25_ASAP7_75t_L g7161 ( 
.A(n_7039),
.B(n_1303),
.C(n_1301),
.D(n_1302),
.Y(n_7161)
);

OAI211xp5_ASAP7_75t_SL g7162 ( 
.A1(n_7088),
.A2(n_1306),
.B(n_1302),
.C(n_1305),
.Y(n_7162)
);

NOR2x1_ASAP7_75t_L g7163 ( 
.A(n_7005),
.B(n_7087),
.Y(n_7163)
);

INVx1_ASAP7_75t_L g7164 ( 
.A(n_7069),
.Y(n_7164)
);

NOR2xp33_ASAP7_75t_L g7165 ( 
.A(n_7042),
.B(n_1305),
.Y(n_7165)
);

AOI22xp5_ASAP7_75t_L g7166 ( 
.A1(n_7086),
.A2(n_1308),
.B1(n_1306),
.B2(n_1307),
.Y(n_7166)
);

OAI221xp5_ASAP7_75t_L g7167 ( 
.A1(n_7084),
.A2(n_1310),
.B1(n_1308),
.B2(n_1309),
.C(n_1311),
.Y(n_7167)
);

OAI211xp5_ASAP7_75t_SL g7168 ( 
.A1(n_7083),
.A2(n_1313),
.B(n_1310),
.C(n_1312),
.Y(n_7168)
);

NOR3xp33_ASAP7_75t_L g7169 ( 
.A(n_7076),
.B(n_1314),
.C(n_1315),
.Y(n_7169)
);

NOR2x1_ASAP7_75t_L g7170 ( 
.A(n_7095),
.B(n_7077),
.Y(n_7170)
);

INVx1_ASAP7_75t_L g7171 ( 
.A(n_7129),
.Y(n_7171)
);

NAND4xp25_ASAP7_75t_L g7172 ( 
.A(n_7137),
.B(n_7045),
.C(n_7070),
.D(n_7014),
.Y(n_7172)
);

NAND3xp33_ASAP7_75t_SL g7173 ( 
.A(n_7160),
.B(n_7019),
.C(n_7034),
.Y(n_7173)
);

OAI311xp33_ASAP7_75t_L g7174 ( 
.A1(n_7110),
.A2(n_7050),
.A3(n_7061),
.B1(n_7016),
.C1(n_7062),
.Y(n_7174)
);

OAI22xp5_ASAP7_75t_L g7175 ( 
.A1(n_7149),
.A2(n_7055),
.B1(n_7025),
.B2(n_1317),
.Y(n_7175)
);

INVx1_ASAP7_75t_L g7176 ( 
.A(n_7119),
.Y(n_7176)
);

NOR3xp33_ASAP7_75t_L g7177 ( 
.A(n_7130),
.B(n_1314),
.C(n_1316),
.Y(n_7177)
);

OAI211xp5_ASAP7_75t_L g7178 ( 
.A1(n_7102),
.A2(n_1320),
.B(n_1318),
.C(n_1319),
.Y(n_7178)
);

A2O1A1Ixp33_ASAP7_75t_L g7179 ( 
.A1(n_7121),
.A2(n_1321),
.B(n_1318),
.C(n_1320),
.Y(n_7179)
);

AOI221x1_ASAP7_75t_L g7180 ( 
.A1(n_7104),
.A2(n_1324),
.B1(n_1322),
.B2(n_1323),
.C(n_1325),
.Y(n_7180)
);

OAI211xp5_ASAP7_75t_SL g7181 ( 
.A1(n_7103),
.A2(n_1325),
.B(n_1322),
.C(n_1323),
.Y(n_7181)
);

NOR2x1_ASAP7_75t_L g7182 ( 
.A(n_7099),
.B(n_1326),
.Y(n_7182)
);

AOI222xp33_ASAP7_75t_L g7183 ( 
.A1(n_7145),
.A2(n_1328),
.B1(n_1331),
.B2(n_1326),
.C1(n_1327),
.C2(n_1330),
.Y(n_7183)
);

NOR2xp67_ASAP7_75t_L g7184 ( 
.A(n_7101),
.B(n_1327),
.Y(n_7184)
);

NOR2x1p5_ASAP7_75t_L g7185 ( 
.A(n_7146),
.B(n_1330),
.Y(n_7185)
);

INVxp67_ASAP7_75t_L g7186 ( 
.A(n_7105),
.Y(n_7186)
);

NOR3x1_ASAP7_75t_L g7187 ( 
.A(n_7107),
.B(n_1331),
.C(n_1332),
.Y(n_7187)
);

NAND4xp75_ASAP7_75t_L g7188 ( 
.A(n_7100),
.B(n_7097),
.C(n_7111),
.D(n_7163),
.Y(n_7188)
);

NAND2xp5_ASAP7_75t_L g7189 ( 
.A(n_7144),
.B(n_1333),
.Y(n_7189)
);

AND4x1_ASAP7_75t_L g7190 ( 
.A(n_7109),
.B(n_1344),
.C(n_1352),
.D(n_1334),
.Y(n_7190)
);

NAND2xp5_ASAP7_75t_SL g7191 ( 
.A(n_7159),
.B(n_1334),
.Y(n_7191)
);

NOR2x1_ASAP7_75t_L g7192 ( 
.A(n_7124),
.B(n_1335),
.Y(n_7192)
);

INVx1_ASAP7_75t_L g7193 ( 
.A(n_7120),
.Y(n_7193)
);

AND2x2_ASAP7_75t_SL g7194 ( 
.A(n_7169),
.B(n_1335),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_7118),
.Y(n_7195)
);

AOI21xp33_ASAP7_75t_L g7196 ( 
.A1(n_7126),
.A2(n_1785),
.B(n_1784),
.Y(n_7196)
);

NOR3xp33_ASAP7_75t_L g7197 ( 
.A(n_7151),
.B(n_7138),
.C(n_7123),
.Y(n_7197)
);

NAND4xp25_ASAP7_75t_L g7198 ( 
.A(n_7114),
.B(n_1340),
.C(n_1337),
.D(n_1338),
.Y(n_7198)
);

NOR2x1_ASAP7_75t_L g7199 ( 
.A(n_7096),
.B(n_1340),
.Y(n_7199)
);

NAND3xp33_ASAP7_75t_L g7200 ( 
.A(n_7134),
.B(n_1341),
.C(n_1342),
.Y(n_7200)
);

OR2x2_ASAP7_75t_L g7201 ( 
.A(n_7142),
.B(n_1341),
.Y(n_7201)
);

INVx1_ASAP7_75t_L g7202 ( 
.A(n_7122),
.Y(n_7202)
);

NAND3xp33_ASAP7_75t_SL g7203 ( 
.A(n_7156),
.B(n_1342),
.C(n_1343),
.Y(n_7203)
);

OAI221xp5_ASAP7_75t_SL g7204 ( 
.A1(n_7112),
.A2(n_1347),
.B1(n_1345),
.B2(n_1346),
.C(n_1348),
.Y(n_7204)
);

AND2x4_ASAP7_75t_L g7205 ( 
.A(n_7117),
.B(n_1346),
.Y(n_7205)
);

NOR3xp33_ASAP7_75t_SL g7206 ( 
.A(n_7162),
.B(n_1348),
.C(n_1349),
.Y(n_7206)
);

NAND3xp33_ASAP7_75t_SL g7207 ( 
.A(n_7135),
.B(n_1350),
.C(n_1351),
.Y(n_7207)
);

NAND3xp33_ASAP7_75t_L g7208 ( 
.A(n_7127),
.B(n_1350),
.C(n_1351),
.Y(n_7208)
);

OAI211xp5_ASAP7_75t_SL g7209 ( 
.A1(n_7164),
.A2(n_1355),
.B(n_1353),
.C(n_1354),
.Y(n_7209)
);

NAND5xp2_ASAP7_75t_L g7210 ( 
.A(n_7133),
.B(n_1355),
.C(n_1353),
.D(n_1354),
.E(n_1356),
.Y(n_7210)
);

AOI322xp5_ASAP7_75t_L g7211 ( 
.A1(n_7140),
.A2(n_1788),
.A3(n_1786),
.B1(n_1789),
.B2(n_1796),
.C1(n_1787),
.C2(n_1785),
.Y(n_7211)
);

NAND4xp75_ASAP7_75t_L g7212 ( 
.A(n_7165),
.B(n_1358),
.C(n_1356),
.D(n_1357),
.Y(n_7212)
);

O2A1O1Ixp33_ASAP7_75t_L g7213 ( 
.A1(n_7148),
.A2(n_1359),
.B(n_1357),
.C(n_1358),
.Y(n_7213)
);

NOR3xp33_ASAP7_75t_L g7214 ( 
.A(n_7139),
.B(n_1360),
.C(n_1362),
.Y(n_7214)
);

NOR2xp33_ASAP7_75t_L g7215 ( 
.A(n_7168),
.B(n_1363),
.Y(n_7215)
);

NOR4xp25_ASAP7_75t_L g7216 ( 
.A(n_7132),
.B(n_1365),
.C(n_1360),
.D(n_1364),
.Y(n_7216)
);

AOI32xp33_ASAP7_75t_L g7217 ( 
.A1(n_7141),
.A2(n_1366),
.A3(n_1364),
.B1(n_1365),
.B2(n_1367),
.Y(n_7217)
);

OR2x2_ASAP7_75t_L g7218 ( 
.A(n_7161),
.B(n_1367),
.Y(n_7218)
);

NAND2xp5_ASAP7_75t_L g7219 ( 
.A(n_7131),
.B(n_1368),
.Y(n_7219)
);

NOR3xp33_ASAP7_75t_SL g7220 ( 
.A(n_7125),
.B(n_7158),
.C(n_7115),
.Y(n_7220)
);

OAI211xp5_ASAP7_75t_SL g7221 ( 
.A1(n_7155),
.A2(n_1371),
.B(n_1368),
.C(n_1370),
.Y(n_7221)
);

AOI221xp5_ASAP7_75t_L g7222 ( 
.A1(n_7106),
.A2(n_1374),
.B1(n_1372),
.B2(n_1373),
.C(n_1375),
.Y(n_7222)
);

NOR2xp33_ASAP7_75t_L g7223 ( 
.A(n_7113),
.B(n_7152),
.Y(n_7223)
);

INVx1_ASAP7_75t_L g7224 ( 
.A(n_7143),
.Y(n_7224)
);

NAND3xp33_ASAP7_75t_SL g7225 ( 
.A(n_7166),
.B(n_1372),
.C(n_1373),
.Y(n_7225)
);

NAND2xp5_ASAP7_75t_SL g7226 ( 
.A(n_7128),
.B(n_1374),
.Y(n_7226)
);

NAND3xp33_ASAP7_75t_SL g7227 ( 
.A(n_7157),
.B(n_1376),
.C(n_1377),
.Y(n_7227)
);

NAND4xp25_ASAP7_75t_SL g7228 ( 
.A(n_7108),
.B(n_1378),
.C(n_1376),
.D(n_1377),
.Y(n_7228)
);

NOR2x1_ASAP7_75t_L g7229 ( 
.A(n_7150),
.B(n_1379),
.Y(n_7229)
);

NOR3xp33_ASAP7_75t_L g7230 ( 
.A(n_7167),
.B(n_7154),
.C(n_7136),
.Y(n_7230)
);

NAND4xp25_ASAP7_75t_L g7231 ( 
.A(n_7147),
.B(n_1381),
.C(n_1379),
.D(n_1380),
.Y(n_7231)
);

AOI221xp5_ASAP7_75t_L g7232 ( 
.A1(n_7098),
.A2(n_1384),
.B1(n_1382),
.B2(n_1383),
.C(n_1385),
.Y(n_7232)
);

OAI22xp5_ASAP7_75t_L g7233 ( 
.A1(n_7153),
.A2(n_1386),
.B1(n_1383),
.B2(n_1384),
.Y(n_7233)
);

NAND2xp5_ASAP7_75t_L g7234 ( 
.A(n_7116),
.B(n_1386),
.Y(n_7234)
);

NAND4xp75_ASAP7_75t_L g7235 ( 
.A(n_7095),
.B(n_1389),
.C(n_1387),
.D(n_1388),
.Y(n_7235)
);

OAI221xp5_ASAP7_75t_L g7236 ( 
.A1(n_7095),
.A2(n_1390),
.B1(n_1387),
.B2(n_1389),
.C(n_1391),
.Y(n_7236)
);

NAND3xp33_ASAP7_75t_SL g7237 ( 
.A(n_7095),
.B(n_1390),
.C(n_1391),
.Y(n_7237)
);

AOI221x1_ASAP7_75t_L g7238 ( 
.A1(n_7095),
.A2(n_1394),
.B1(n_1392),
.B2(n_1393),
.C(n_1395),
.Y(n_7238)
);

AOI221xp5_ASAP7_75t_SL g7239 ( 
.A1(n_7095),
.A2(n_1395),
.B1(n_1392),
.B2(n_1394),
.C(n_1396),
.Y(n_7239)
);

NOR4xp25_ASAP7_75t_L g7240 ( 
.A(n_7095),
.B(n_1398),
.C(n_1396),
.D(n_1397),
.Y(n_7240)
);

OAI21xp5_ASAP7_75t_L g7241 ( 
.A1(n_7095),
.A2(n_1397),
.B(n_1398),
.Y(n_7241)
);

NOR2xp33_ASAP7_75t_L g7242 ( 
.A(n_7110),
.B(n_1400),
.Y(n_7242)
);

NOR2x1_ASAP7_75t_L g7243 ( 
.A(n_7095),
.B(n_1399),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_7110),
.B(n_1399),
.Y(n_7244)
);

A2O1A1Ixp33_ASAP7_75t_L g7245 ( 
.A1(n_7095),
.A2(n_1403),
.B(n_1401),
.C(n_1402),
.Y(n_7245)
);

NAND3xp33_ASAP7_75t_L g7246 ( 
.A(n_7095),
.B(n_1401),
.C(n_1403),
.Y(n_7246)
);

AOI22xp5_ASAP7_75t_L g7247 ( 
.A1(n_7095),
.A2(n_1406),
.B1(n_1404),
.B2(n_1405),
.Y(n_7247)
);

NAND3xp33_ASAP7_75t_L g7248 ( 
.A(n_7095),
.B(n_1404),
.C(n_1405),
.Y(n_7248)
);

AOI21xp5_ASAP7_75t_L g7249 ( 
.A1(n_7095),
.A2(n_1407),
.B(n_1409),
.Y(n_7249)
);

NOR3xp33_ASAP7_75t_L g7250 ( 
.A(n_7095),
.B(n_1407),
.C(n_1409),
.Y(n_7250)
);

XNOR2xp5_ASAP7_75t_L g7251 ( 
.A(n_7184),
.B(n_7188),
.Y(n_7251)
);

OAI22xp33_ASAP7_75t_SL g7252 ( 
.A1(n_7202),
.A2(n_1412),
.B1(n_1410),
.B2(n_1411),
.Y(n_7252)
);

NAND4xp25_ASAP7_75t_SL g7253 ( 
.A(n_7239),
.B(n_1412),
.C(n_1410),
.D(n_1411),
.Y(n_7253)
);

AOI22xp33_ASAP7_75t_SL g7254 ( 
.A1(n_7176),
.A2(n_1415),
.B1(n_1413),
.B2(n_1414),
.Y(n_7254)
);

AOI221x1_ASAP7_75t_L g7255 ( 
.A1(n_7197),
.A2(n_1779),
.B1(n_1780),
.B2(n_1778),
.C(n_1776),
.Y(n_7255)
);

AOI221xp5_ASAP7_75t_L g7256 ( 
.A1(n_7186),
.A2(n_1416),
.B1(n_1413),
.B2(n_1415),
.C(n_1417),
.Y(n_7256)
);

NAND4xp25_ASAP7_75t_L g7257 ( 
.A(n_7210),
.B(n_1419),
.C(n_1417),
.D(n_1418),
.Y(n_7257)
);

NOR2xp33_ASAP7_75t_L g7258 ( 
.A(n_7224),
.B(n_1419),
.Y(n_7258)
);

NAND2xp5_ASAP7_75t_L g7259 ( 
.A(n_7171),
.B(n_7199),
.Y(n_7259)
);

OAI22xp5_ASAP7_75t_L g7260 ( 
.A1(n_7201),
.A2(n_1424),
.B1(n_1422),
.B2(n_1423),
.Y(n_7260)
);

INVx1_ASAP7_75t_L g7261 ( 
.A(n_7243),
.Y(n_7261)
);

NOR2xp33_ASAP7_75t_L g7262 ( 
.A(n_7193),
.B(n_1422),
.Y(n_7262)
);

NAND3xp33_ASAP7_75t_SL g7263 ( 
.A(n_7195),
.B(n_1425),
.C(n_1424),
.Y(n_7263)
);

AOI22xp5_ASAP7_75t_L g7264 ( 
.A1(n_7223),
.A2(n_1426),
.B1(n_1423),
.B2(n_1425),
.Y(n_7264)
);

OAI21xp33_ASAP7_75t_L g7265 ( 
.A1(n_7220),
.A2(n_1427),
.B(n_1428),
.Y(n_7265)
);

NOR2x1_ASAP7_75t_L g7266 ( 
.A(n_7173),
.B(n_7170),
.Y(n_7266)
);

OAI21xp33_ASAP7_75t_SL g7267 ( 
.A1(n_7183),
.A2(n_1427),
.B(n_1428),
.Y(n_7267)
);

AOI221xp5_ASAP7_75t_L g7268 ( 
.A1(n_7240),
.A2(n_1431),
.B1(n_1429),
.B2(n_1430),
.C(n_1433),
.Y(n_7268)
);

NOR2xp33_ASAP7_75t_L g7269 ( 
.A(n_7203),
.B(n_1430),
.Y(n_7269)
);

AOI22xp33_ASAP7_75t_SL g7270 ( 
.A1(n_7205),
.A2(n_1434),
.B1(n_1431),
.B2(n_1433),
.Y(n_7270)
);

AOI21xp33_ASAP7_75t_L g7271 ( 
.A1(n_7182),
.A2(n_1436),
.B(n_1435),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_7205),
.Y(n_7272)
);

AOI22xp5_ASAP7_75t_L g7273 ( 
.A1(n_7175),
.A2(n_1437),
.B1(n_1434),
.B2(n_1436),
.Y(n_7273)
);

NAND2xp5_ASAP7_75t_L g7274 ( 
.A(n_7194),
.B(n_1437),
.Y(n_7274)
);

INVxp67_ASAP7_75t_L g7275 ( 
.A(n_7215),
.Y(n_7275)
);

CKINVDCx20_ASAP7_75t_R g7276 ( 
.A(n_7189),
.Y(n_7276)
);

INVxp67_ASAP7_75t_L g7277 ( 
.A(n_7229),
.Y(n_7277)
);

NOR2x1_ASAP7_75t_L g7278 ( 
.A(n_7244),
.B(n_1438),
.Y(n_7278)
);

HB1xp67_ASAP7_75t_L g7279 ( 
.A(n_7185),
.Y(n_7279)
);

OAI211xp5_ASAP7_75t_L g7280 ( 
.A1(n_7211),
.A2(n_1440),
.B(n_1438),
.C(n_1439),
.Y(n_7280)
);

AND2x4_ASAP7_75t_L g7281 ( 
.A(n_7192),
.B(n_1439),
.Y(n_7281)
);

NOR2x1p5_ASAP7_75t_L g7282 ( 
.A(n_7235),
.B(n_1440),
.Y(n_7282)
);

INVx1_ASAP7_75t_SL g7283 ( 
.A(n_7218),
.Y(n_7283)
);

OAI22xp5_ASAP7_75t_L g7284 ( 
.A1(n_7247),
.A2(n_1443),
.B1(n_1441),
.B2(n_1442),
.Y(n_7284)
);

A2O1A1Ixp33_ASAP7_75t_L g7285 ( 
.A1(n_7213),
.A2(n_1444),
.B(n_1442),
.C(n_1443),
.Y(n_7285)
);

OAI211xp5_ASAP7_75t_L g7286 ( 
.A1(n_7217),
.A2(n_7241),
.B(n_7219),
.C(n_7249),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_7190),
.Y(n_7287)
);

AOI221xp5_ASAP7_75t_L g7288 ( 
.A1(n_7216),
.A2(n_1446),
.B1(n_1444),
.B2(n_1445),
.C(n_1447),
.Y(n_7288)
);

NAND2xp5_ASAP7_75t_L g7289 ( 
.A(n_7206),
.B(n_1446),
.Y(n_7289)
);

NOR2xp33_ASAP7_75t_R g7290 ( 
.A(n_7237),
.B(n_1447),
.Y(n_7290)
);

NAND5xp2_ASAP7_75t_L g7291 ( 
.A(n_7230),
.B(n_1450),
.C(n_1448),
.D(n_1449),
.E(n_1451),
.Y(n_7291)
);

CKINVDCx16_ASAP7_75t_R g7292 ( 
.A(n_7227),
.Y(n_7292)
);

NAND2xp5_ASAP7_75t_L g7293 ( 
.A(n_7177),
.B(n_1448),
.Y(n_7293)
);

AND2x4_ASAP7_75t_L g7294 ( 
.A(n_7214),
.B(n_1449),
.Y(n_7294)
);

NOR3xp33_ASAP7_75t_L g7295 ( 
.A(n_7242),
.B(n_1451),
.C(n_1453),
.Y(n_7295)
);

AOI21xp5_ASAP7_75t_L g7296 ( 
.A1(n_7191),
.A2(n_1454),
.B(n_1456),
.Y(n_7296)
);

O2A1O1Ixp33_ASAP7_75t_L g7297 ( 
.A1(n_7245),
.A2(n_1458),
.B(n_1456),
.C(n_1457),
.Y(n_7297)
);

OAI21xp5_ASAP7_75t_L g7298 ( 
.A1(n_7172),
.A2(n_1457),
.B(n_1458),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_7180),
.Y(n_7299)
);

AOI21xp33_ASAP7_75t_SL g7300 ( 
.A1(n_7196),
.A2(n_1468),
.B(n_1459),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_7212),
.Y(n_7301)
);

INVx1_ASAP7_75t_L g7302 ( 
.A(n_7238),
.Y(n_7302)
);

O2A1O1Ixp33_ASAP7_75t_L g7303 ( 
.A1(n_7250),
.A2(n_1461),
.B(n_1459),
.C(n_1460),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_7187),
.Y(n_7304)
);

A2O1A1Ixp33_ASAP7_75t_L g7305 ( 
.A1(n_7246),
.A2(n_1463),
.B(n_1461),
.C(n_1462),
.Y(n_7305)
);

NOR2xp33_ASAP7_75t_L g7306 ( 
.A(n_7181),
.B(n_1462),
.Y(n_7306)
);

INVx2_ASAP7_75t_L g7307 ( 
.A(n_7234),
.Y(n_7307)
);

BUFx2_ASAP7_75t_L g7308 ( 
.A(n_7198),
.Y(n_7308)
);

NAND2xp5_ASAP7_75t_SL g7309 ( 
.A(n_7222),
.B(n_1463),
.Y(n_7309)
);

AOI22xp5_ASAP7_75t_SL g7310 ( 
.A1(n_7233),
.A2(n_7228),
.B1(n_7209),
.B2(n_7174),
.Y(n_7310)
);

INVx2_ASAP7_75t_SL g7311 ( 
.A(n_7248),
.Y(n_7311)
);

AOI211xp5_ASAP7_75t_L g7312 ( 
.A1(n_7204),
.A2(n_1467),
.B(n_1464),
.C(n_1466),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_7178),
.Y(n_7313)
);

INVxp33_ASAP7_75t_L g7314 ( 
.A(n_7231),
.Y(n_7314)
);

NOR2xp33_ASAP7_75t_R g7315 ( 
.A(n_7207),
.B(n_1464),
.Y(n_7315)
);

AND2x2_ASAP7_75t_L g7316 ( 
.A(n_7179),
.B(n_1467),
.Y(n_7316)
);

INVx1_ASAP7_75t_SL g7317 ( 
.A(n_7226),
.Y(n_7317)
);

OAI21xp33_ASAP7_75t_L g7318 ( 
.A1(n_7221),
.A2(n_1470),
.B(n_1472),
.Y(n_7318)
);

INVx1_ASAP7_75t_SL g7319 ( 
.A(n_7200),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_7232),
.B(n_1470),
.Y(n_7320)
);

INVx3_ASAP7_75t_SL g7321 ( 
.A(n_7225),
.Y(n_7321)
);

AND2x2_ASAP7_75t_L g7322 ( 
.A(n_7208),
.B(n_1472),
.Y(n_7322)
);

NOR2x1_ASAP7_75t_L g7323 ( 
.A(n_7236),
.B(n_1473),
.Y(n_7323)
);

NAND4xp75_ASAP7_75t_L g7324 ( 
.A(n_7266),
.B(n_1475),
.C(n_1473),
.D(n_1474),
.Y(n_7324)
);

NOR2x1_ASAP7_75t_L g7325 ( 
.A(n_7251),
.B(n_1475),
.Y(n_7325)
);

AOI22xp5_ASAP7_75t_L g7326 ( 
.A1(n_7304),
.A2(n_7269),
.B1(n_7283),
.B2(n_7302),
.Y(n_7326)
);

INVx1_ASAP7_75t_L g7327 ( 
.A(n_7299),
.Y(n_7327)
);

NOR2x1_ASAP7_75t_L g7328 ( 
.A(n_7259),
.B(n_1476),
.Y(n_7328)
);

INVx3_ASAP7_75t_L g7329 ( 
.A(n_7281),
.Y(n_7329)
);

XOR2xp5_ASAP7_75t_L g7330 ( 
.A(n_7276),
.B(n_1478),
.Y(n_7330)
);

INVx1_ASAP7_75t_L g7331 ( 
.A(n_7261),
.Y(n_7331)
);

NAND4xp75_ASAP7_75t_L g7332 ( 
.A(n_7278),
.B(n_1480),
.C(n_1478),
.D(n_1479),
.Y(n_7332)
);

OAI22xp33_ASAP7_75t_L g7333 ( 
.A1(n_7314),
.A2(n_1481),
.B1(n_1479),
.B2(n_1480),
.Y(n_7333)
);

NOR2xp33_ASAP7_75t_L g7334 ( 
.A(n_7272),
.B(n_1482),
.Y(n_7334)
);

AOI22xp33_ASAP7_75t_L g7335 ( 
.A1(n_7279),
.A2(n_1485),
.B1(n_1482),
.B2(n_1483),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_7281),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_7289),
.Y(n_7337)
);

NOR3xp33_ASAP7_75t_L g7338 ( 
.A(n_7292),
.B(n_1486),
.C(n_1487),
.Y(n_7338)
);

INVx1_ASAP7_75t_L g7339 ( 
.A(n_7277),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_7274),
.Y(n_7340)
);

INVxp67_ASAP7_75t_L g7341 ( 
.A(n_7258),
.Y(n_7341)
);

NAND2xp5_ASAP7_75t_L g7342 ( 
.A(n_7287),
.B(n_1486),
.Y(n_7342)
);

NOR2xp67_ASAP7_75t_L g7343 ( 
.A(n_7291),
.B(n_1487),
.Y(n_7343)
);

INVx2_ASAP7_75t_L g7344 ( 
.A(n_7282),
.Y(n_7344)
);

NOR3xp33_ASAP7_75t_L g7345 ( 
.A(n_7307),
.B(n_1488),
.C(n_1489),
.Y(n_7345)
);

NAND2x1p5_ASAP7_75t_L g7346 ( 
.A(n_7301),
.B(n_1488),
.Y(n_7346)
);

HB1xp67_ASAP7_75t_L g7347 ( 
.A(n_7290),
.Y(n_7347)
);

INVx1_ASAP7_75t_L g7348 ( 
.A(n_7257),
.Y(n_7348)
);

INVx2_ASAP7_75t_L g7349 ( 
.A(n_7294),
.Y(n_7349)
);

XOR2x1_ASAP7_75t_L g7350 ( 
.A(n_7313),
.B(n_1489),
.Y(n_7350)
);

INVx2_ASAP7_75t_L g7351 ( 
.A(n_7294),
.Y(n_7351)
);

NAND4xp75_ASAP7_75t_L g7352 ( 
.A(n_7255),
.B(n_1492),
.C(n_1490),
.D(n_1491),
.Y(n_7352)
);

AND3x2_ASAP7_75t_L g7353 ( 
.A(n_7262),
.B(n_1490),
.C(n_1492),
.Y(n_7353)
);

INVx2_ASAP7_75t_L g7354 ( 
.A(n_7308),
.Y(n_7354)
);

INVx1_ASAP7_75t_L g7355 ( 
.A(n_7310),
.Y(n_7355)
);

AND2x4_ASAP7_75t_L g7356 ( 
.A(n_7311),
.B(n_1493),
.Y(n_7356)
);

AO22x1_ASAP7_75t_L g7357 ( 
.A1(n_7298),
.A2(n_1496),
.B1(n_1494),
.B2(n_1495),
.Y(n_7357)
);

NOR2x1_ASAP7_75t_L g7358 ( 
.A(n_7263),
.B(n_7253),
.Y(n_7358)
);

NAND4xp75_ASAP7_75t_L g7359 ( 
.A(n_7271),
.B(n_1496),
.C(n_1494),
.D(n_1495),
.Y(n_7359)
);

OR2x2_ASAP7_75t_L g7360 ( 
.A(n_7321),
.B(n_1497),
.Y(n_7360)
);

AND2x2_ASAP7_75t_L g7361 ( 
.A(n_7322),
.B(n_1497),
.Y(n_7361)
);

NOR3xp33_ASAP7_75t_L g7362 ( 
.A(n_7275),
.B(n_1498),
.C(n_1499),
.Y(n_7362)
);

INVx1_ASAP7_75t_L g7363 ( 
.A(n_7252),
.Y(n_7363)
);

XNOR2xp5_ASAP7_75t_L g7364 ( 
.A(n_7312),
.B(n_1499),
.Y(n_7364)
);

AOI22xp5_ASAP7_75t_L g7365 ( 
.A1(n_7265),
.A2(n_1502),
.B1(n_1500),
.B2(n_1501),
.Y(n_7365)
);

INVx1_ASAP7_75t_L g7366 ( 
.A(n_7306),
.Y(n_7366)
);

NAND2xp5_ASAP7_75t_L g7367 ( 
.A(n_7270),
.B(n_1500),
.Y(n_7367)
);

NAND2xp5_ASAP7_75t_L g7368 ( 
.A(n_7319),
.B(n_1501),
.Y(n_7368)
);

INVxp67_ASAP7_75t_L g7369 ( 
.A(n_7293),
.Y(n_7369)
);

NAND2x1p5_ASAP7_75t_L g7370 ( 
.A(n_7317),
.B(n_1502),
.Y(n_7370)
);

INVx1_ASAP7_75t_L g7371 ( 
.A(n_7316),
.Y(n_7371)
);

OAI22xp5_ASAP7_75t_L g7372 ( 
.A1(n_7273),
.A2(n_7254),
.B1(n_7285),
.B2(n_7305),
.Y(n_7372)
);

XNOR2x1_ASAP7_75t_L g7373 ( 
.A(n_7323),
.B(n_1503),
.Y(n_7373)
);

NOR2x1_ASAP7_75t_L g7374 ( 
.A(n_7260),
.B(n_1503),
.Y(n_7374)
);

NOR2x1_ASAP7_75t_L g7375 ( 
.A(n_7280),
.B(n_1504),
.Y(n_7375)
);

NAND4xp75_ASAP7_75t_L g7376 ( 
.A(n_7267),
.B(n_1506),
.C(n_1504),
.D(n_1505),
.Y(n_7376)
);

INVx1_ASAP7_75t_SL g7377 ( 
.A(n_7315),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_7318),
.Y(n_7378)
);

INVx1_ASAP7_75t_L g7379 ( 
.A(n_7303),
.Y(n_7379)
);

INVxp67_ASAP7_75t_L g7380 ( 
.A(n_7320),
.Y(n_7380)
);

NOR2x1_ASAP7_75t_L g7381 ( 
.A(n_7286),
.B(n_1508),
.Y(n_7381)
);

HB1xp67_ASAP7_75t_L g7382 ( 
.A(n_7295),
.Y(n_7382)
);

AO211x2_ASAP7_75t_L g7383 ( 
.A1(n_7327),
.A2(n_7296),
.B(n_7300),
.C(n_7288),
.Y(n_7383)
);

NOR4xp25_ASAP7_75t_L g7384 ( 
.A(n_7355),
.B(n_7309),
.C(n_7297),
.D(n_7268),
.Y(n_7384)
);

NOR3xp33_ASAP7_75t_SL g7385 ( 
.A(n_7336),
.B(n_7284),
.C(n_7256),
.Y(n_7385)
);

AND2x4_ASAP7_75t_L g7386 ( 
.A(n_7329),
.B(n_7264),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_7350),
.Y(n_7387)
);

AOI21xp5_ASAP7_75t_L g7388 ( 
.A1(n_7339),
.A2(n_1509),
.B(n_1510),
.Y(n_7388)
);

NOR2xp67_ASAP7_75t_L g7389 ( 
.A(n_7360),
.B(n_1510),
.Y(n_7389)
);

NOR2x1_ASAP7_75t_L g7390 ( 
.A(n_7331),
.B(n_1511),
.Y(n_7390)
);

NOR3xp33_ASAP7_75t_L g7391 ( 
.A(n_7354),
.B(n_1511),
.C(n_1512),
.Y(n_7391)
);

O2A1O1Ixp33_ASAP7_75t_L g7392 ( 
.A1(n_7347),
.A2(n_7344),
.B(n_7341),
.C(n_7363),
.Y(n_7392)
);

A2O1A1Ixp33_ASAP7_75t_L g7393 ( 
.A1(n_7326),
.A2(n_1514),
.B(n_1512),
.C(n_1513),
.Y(n_7393)
);

AO211x2_ASAP7_75t_L g7394 ( 
.A1(n_7371),
.A2(n_7348),
.B(n_7366),
.C(n_7337),
.Y(n_7394)
);

NOR3xp33_ASAP7_75t_SL g7395 ( 
.A(n_7340),
.B(n_1514),
.C(n_1515),
.Y(n_7395)
);

OAI22xp33_ASAP7_75t_L g7396 ( 
.A1(n_7365),
.A2(n_7377),
.B1(n_7367),
.B2(n_7343),
.Y(n_7396)
);

NOR4xp25_ASAP7_75t_L g7397 ( 
.A(n_7349),
.B(n_1518),
.C(n_1516),
.D(n_1517),
.Y(n_7397)
);

NAND5xp2_ASAP7_75t_L g7398 ( 
.A(n_7370),
.B(n_1521),
.C(n_1519),
.D(n_1520),
.E(n_1522),
.Y(n_7398)
);

HB1xp67_ASAP7_75t_L g7399 ( 
.A(n_7325),
.Y(n_7399)
);

OR2x6_ASAP7_75t_L g7400 ( 
.A(n_7351),
.B(n_1520),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_7328),
.Y(n_7401)
);

AND2x2_ASAP7_75t_L g7402 ( 
.A(n_7381),
.B(n_1521),
.Y(n_7402)
);

NOR2x1_ASAP7_75t_L g7403 ( 
.A(n_7324),
.B(n_1522),
.Y(n_7403)
);

AND2x4_ASAP7_75t_L g7404 ( 
.A(n_7358),
.B(n_1810),
.Y(n_7404)
);

NOR4xp25_ASAP7_75t_L g7405 ( 
.A(n_7380),
.B(n_1525),
.C(n_1523),
.D(n_1524),
.Y(n_7405)
);

NAND4xp75_ASAP7_75t_L g7406 ( 
.A(n_7375),
.B(n_7374),
.C(n_7361),
.D(n_7379),
.Y(n_7406)
);

INVx2_ASAP7_75t_SL g7407 ( 
.A(n_7346),
.Y(n_7407)
);

NOR3xp33_ASAP7_75t_L g7408 ( 
.A(n_7369),
.B(n_1523),
.C(n_1524),
.Y(n_7408)
);

NAND3xp33_ASAP7_75t_L g7409 ( 
.A(n_7373),
.B(n_1525),
.C(n_1526),
.Y(n_7409)
);

NOR3xp33_ASAP7_75t_SL g7410 ( 
.A(n_7376),
.B(n_1526),
.C(n_1527),
.Y(n_7410)
);

XNOR2xp5_ASAP7_75t_L g7411 ( 
.A(n_7330),
.B(n_1527),
.Y(n_7411)
);

OAI211xp5_ASAP7_75t_L g7412 ( 
.A1(n_7378),
.A2(n_1530),
.B(n_1528),
.C(n_1529),
.Y(n_7412)
);

HB1xp67_ASAP7_75t_L g7413 ( 
.A(n_7356),
.Y(n_7413)
);

OAI211xp5_ASAP7_75t_SL g7414 ( 
.A1(n_7382),
.A2(n_1530),
.B(n_1528),
.C(n_1529),
.Y(n_7414)
);

INVx1_ASAP7_75t_SL g7415 ( 
.A(n_7353),
.Y(n_7415)
);

NAND3xp33_ASAP7_75t_SL g7416 ( 
.A(n_7345),
.B(n_1531),
.C(n_1532),
.Y(n_7416)
);

INVx1_ASAP7_75t_L g7417 ( 
.A(n_7356),
.Y(n_7417)
);

NOR3xp33_ASAP7_75t_SL g7418 ( 
.A(n_7352),
.B(n_1531),
.C(n_1532),
.Y(n_7418)
);

XNOR2xp5_ASAP7_75t_L g7419 ( 
.A(n_7364),
.B(n_1533),
.Y(n_7419)
);

NAND5xp2_ASAP7_75t_L g7420 ( 
.A(n_7338),
.B(n_1535),
.C(n_1533),
.D(n_1534),
.E(n_1536),
.Y(n_7420)
);

NAND4xp75_ASAP7_75t_L g7421 ( 
.A(n_7368),
.B(n_7334),
.C(n_7342),
.D(n_7332),
.Y(n_7421)
);

NAND3xp33_ASAP7_75t_SL g7422 ( 
.A(n_7362),
.B(n_1534),
.C(n_1536),
.Y(n_7422)
);

AND2x2_ASAP7_75t_L g7423 ( 
.A(n_7359),
.B(n_1537),
.Y(n_7423)
);

NAND4xp25_ASAP7_75t_L g7424 ( 
.A(n_7372),
.B(n_1540),
.C(n_1538),
.D(n_1539),
.Y(n_7424)
);

OAI211xp5_ASAP7_75t_SL g7425 ( 
.A1(n_7335),
.A2(n_1541),
.B(n_1539),
.C(n_1540),
.Y(n_7425)
);

AND5x1_ASAP7_75t_L g7426 ( 
.A(n_7357),
.B(n_1543),
.C(n_1541),
.D(n_1542),
.E(n_1544),
.Y(n_7426)
);

NAND4xp25_ASAP7_75t_L g7427 ( 
.A(n_7333),
.B(n_1544),
.C(n_1542),
.D(n_1543),
.Y(n_7427)
);

NAND4xp75_ASAP7_75t_L g7428 ( 
.A(n_7327),
.B(n_1548),
.C(n_1545),
.D(n_1546),
.Y(n_7428)
);

NAND4xp75_ASAP7_75t_L g7429 ( 
.A(n_7327),
.B(n_1550),
.C(n_1546),
.D(n_1549),
.Y(n_7429)
);

HB1xp67_ASAP7_75t_L g7430 ( 
.A(n_7389),
.Y(n_7430)
);

O2A1O1Ixp33_ASAP7_75t_L g7431 ( 
.A1(n_7399),
.A2(n_1551),
.B(n_1549),
.C(n_1550),
.Y(n_7431)
);

AND2x2_ASAP7_75t_L g7432 ( 
.A(n_7413),
.B(n_1552),
.Y(n_7432)
);

HB1xp67_ASAP7_75t_L g7433 ( 
.A(n_7400),
.Y(n_7433)
);

INVx1_ASAP7_75t_L g7434 ( 
.A(n_7390),
.Y(n_7434)
);

CKINVDCx16_ASAP7_75t_R g7435 ( 
.A(n_7387),
.Y(n_7435)
);

BUFx2_ASAP7_75t_L g7436 ( 
.A(n_7400),
.Y(n_7436)
);

CKINVDCx16_ASAP7_75t_R g7437 ( 
.A(n_7407),
.Y(n_7437)
);

INVx1_ASAP7_75t_L g7438 ( 
.A(n_7402),
.Y(n_7438)
);

CKINVDCx5p33_ASAP7_75t_R g7439 ( 
.A(n_7417),
.Y(n_7439)
);

XNOR2xp5_ASAP7_75t_L g7440 ( 
.A(n_7394),
.B(n_1553),
.Y(n_7440)
);

CKINVDCx5p33_ASAP7_75t_R g7441 ( 
.A(n_7415),
.Y(n_7441)
);

NAND2xp5_ASAP7_75t_L g7442 ( 
.A(n_7401),
.B(n_7392),
.Y(n_7442)
);

INVx1_ASAP7_75t_SL g7443 ( 
.A(n_7404),
.Y(n_7443)
);

INVx1_ASAP7_75t_L g7444 ( 
.A(n_7404),
.Y(n_7444)
);

INVx1_ASAP7_75t_L g7445 ( 
.A(n_7411),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_7406),
.Y(n_7446)
);

CKINVDCx16_ASAP7_75t_R g7447 ( 
.A(n_7386),
.Y(n_7447)
);

CKINVDCx5p33_ASAP7_75t_R g7448 ( 
.A(n_7386),
.Y(n_7448)
);

BUFx4f_ASAP7_75t_SL g7449 ( 
.A(n_7423),
.Y(n_7449)
);

HB1xp67_ASAP7_75t_L g7450 ( 
.A(n_7419),
.Y(n_7450)
);

NOR2xp67_ASAP7_75t_L g7451 ( 
.A(n_7398),
.B(n_1553),
.Y(n_7451)
);

CKINVDCx5p33_ASAP7_75t_R g7452 ( 
.A(n_7385),
.Y(n_7452)
);

INVx2_ASAP7_75t_SL g7453 ( 
.A(n_7403),
.Y(n_7453)
);

NOR2xp33_ASAP7_75t_R g7454 ( 
.A(n_7422),
.B(n_7416),
.Y(n_7454)
);

OR2x2_ASAP7_75t_L g7455 ( 
.A(n_7420),
.B(n_1554),
.Y(n_7455)
);

HB1xp67_ASAP7_75t_L g7456 ( 
.A(n_7421),
.Y(n_7456)
);

AOI22x1_ASAP7_75t_L g7457 ( 
.A1(n_7388),
.A2(n_1557),
.B1(n_1555),
.B2(n_1556),
.Y(n_7457)
);

HB1xp67_ASAP7_75t_L g7458 ( 
.A(n_7383),
.Y(n_7458)
);

OAI22xp33_ASAP7_75t_L g7459 ( 
.A1(n_7435),
.A2(n_7424),
.B1(n_7427),
.B2(n_7409),
.Y(n_7459)
);

AOI31xp33_ASAP7_75t_L g7460 ( 
.A1(n_7440),
.A2(n_7433),
.A3(n_7448),
.B(n_7443),
.Y(n_7460)
);

AOI322xp5_ASAP7_75t_L g7461 ( 
.A1(n_7447),
.A2(n_7396),
.A3(n_7418),
.B1(n_7410),
.B2(n_7395),
.C1(n_7391),
.C2(n_7408),
.Y(n_7461)
);

AOI322xp5_ASAP7_75t_L g7462 ( 
.A1(n_7458),
.A2(n_7393),
.A3(n_7426),
.B1(n_7384),
.B2(n_7425),
.C1(n_7405),
.C2(n_7397),
.Y(n_7462)
);

OAI221xp5_ASAP7_75t_L g7463 ( 
.A1(n_7442),
.A2(n_7446),
.B1(n_7452),
.B2(n_7456),
.C(n_7441),
.Y(n_7463)
);

AOI322xp5_ASAP7_75t_L g7464 ( 
.A1(n_7437),
.A2(n_7414),
.A3(n_7429),
.B1(n_7428),
.B2(n_7412),
.C1(n_1558),
.C2(n_1562),
.Y(n_7464)
);

INVx2_ASAP7_75t_L g7465 ( 
.A(n_7436),
.Y(n_7465)
);

OAI211xp5_ASAP7_75t_L g7466 ( 
.A1(n_7434),
.A2(n_1558),
.B(n_1556),
.C(n_1557),
.Y(n_7466)
);

NAND3xp33_ASAP7_75t_L g7467 ( 
.A(n_7430),
.B(n_1559),
.C(n_1560),
.Y(n_7467)
);

OAI221xp5_ASAP7_75t_L g7468 ( 
.A1(n_7453),
.A2(n_7439),
.B1(n_7451),
.B2(n_7457),
.C(n_7438),
.Y(n_7468)
);

NAND2xp5_ASAP7_75t_L g7469 ( 
.A(n_7444),
.B(n_1807),
.Y(n_7469)
);

AOI322xp5_ASAP7_75t_L g7470 ( 
.A1(n_7450),
.A2(n_1567),
.A3(n_1566),
.B1(n_1564),
.B2(n_1562),
.C1(n_1563),
.C2(n_1565),
.Y(n_7470)
);

AOI221xp5_ASAP7_75t_SL g7471 ( 
.A1(n_7445),
.A2(n_1566),
.B1(n_1563),
.B2(n_1565),
.C(n_1567),
.Y(n_7471)
);

OAI221xp5_ASAP7_75t_L g7472 ( 
.A1(n_7455),
.A2(n_1570),
.B1(n_1568),
.B2(n_1569),
.C(n_1571),
.Y(n_7472)
);

HB1xp67_ASAP7_75t_L g7473 ( 
.A(n_7432),
.Y(n_7473)
);

NOR2x1_ASAP7_75t_L g7474 ( 
.A(n_7431),
.B(n_1569),
.Y(n_7474)
);

OAI221xp5_ASAP7_75t_L g7475 ( 
.A1(n_7449),
.A2(n_1572),
.B1(n_1570),
.B2(n_1571),
.C(n_1573),
.Y(n_7475)
);

INVx1_ASAP7_75t_L g7476 ( 
.A(n_7454),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7447),
.Y(n_7477)
);

AOI322xp5_ASAP7_75t_L g7478 ( 
.A1(n_7447),
.A2(n_1580),
.A3(n_1579),
.B1(n_1577),
.B2(n_1574),
.C1(n_1576),
.C2(n_1578),
.Y(n_7478)
);

AOI22xp5_ASAP7_75t_L g7479 ( 
.A1(n_7477),
.A2(n_7465),
.B1(n_7463),
.B2(n_7476),
.Y(n_7479)
);

AOI22xp5_ASAP7_75t_L g7480 ( 
.A1(n_7473),
.A2(n_1578),
.B1(n_1576),
.B2(n_1577),
.Y(n_7480)
);

OAI22x1_ASAP7_75t_L g7481 ( 
.A1(n_7474),
.A2(n_1582),
.B1(n_1579),
.B2(n_1581),
.Y(n_7481)
);

INVx1_ASAP7_75t_L g7482 ( 
.A(n_7460),
.Y(n_7482)
);

OA22x2_ASAP7_75t_L g7483 ( 
.A1(n_7466),
.A2(n_1584),
.B1(n_1581),
.B2(n_1582),
.Y(n_7483)
);

OAI22x1_ASAP7_75t_L g7484 ( 
.A1(n_7467),
.A2(n_1587),
.B1(n_1585),
.B2(n_1586),
.Y(n_7484)
);

AOI211xp5_ASAP7_75t_SL g7485 ( 
.A1(n_7468),
.A2(n_1590),
.B(n_1585),
.C(n_1588),
.Y(n_7485)
);

OAI22x1_ASAP7_75t_L g7486 ( 
.A1(n_7469),
.A2(n_1592),
.B1(n_1590),
.B2(n_1591),
.Y(n_7486)
);

OAI22xp5_ASAP7_75t_L g7487 ( 
.A1(n_7472),
.A2(n_1594),
.B1(n_1591),
.B2(n_1593),
.Y(n_7487)
);

HB1xp67_ASAP7_75t_L g7488 ( 
.A(n_7475),
.Y(n_7488)
);

OAI22x1_ASAP7_75t_L g7489 ( 
.A1(n_7461),
.A2(n_7462),
.B1(n_7459),
.B2(n_7471),
.Y(n_7489)
);

AOI22xp5_ASAP7_75t_L g7490 ( 
.A1(n_7464),
.A2(n_1597),
.B1(n_1594),
.B2(n_1596),
.Y(n_7490)
);

NAND3xp33_ASAP7_75t_L g7491 ( 
.A(n_7479),
.B(n_7478),
.C(n_7470),
.Y(n_7491)
);

NAND4xp25_ASAP7_75t_L g7492 ( 
.A(n_7482),
.B(n_1600),
.C(n_1596),
.D(n_1599),
.Y(n_7492)
);

AOI211xp5_ASAP7_75t_L g7493 ( 
.A1(n_7488),
.A2(n_1601),
.B(n_1599),
.C(n_1600),
.Y(n_7493)
);

XOR2xp5_ASAP7_75t_L g7494 ( 
.A(n_7489),
.B(n_7490),
.Y(n_7494)
);

NOR3xp33_ASAP7_75t_SL g7495 ( 
.A(n_7487),
.B(n_1602),
.C(n_1603),
.Y(n_7495)
);

NOR3xp33_ASAP7_75t_L g7496 ( 
.A(n_7480),
.B(n_1602),
.C(n_1604),
.Y(n_7496)
);

AOI221xp5_ASAP7_75t_L g7497 ( 
.A1(n_7481),
.A2(n_1607),
.B1(n_1605),
.B2(n_1606),
.C(n_1608),
.Y(n_7497)
);

INVx3_ASAP7_75t_L g7498 ( 
.A(n_7494),
.Y(n_7498)
);

OAI22xp5_ASAP7_75t_L g7499 ( 
.A1(n_7493),
.A2(n_7483),
.B1(n_7485),
.B2(n_7484),
.Y(n_7499)
);

CKINVDCx20_ASAP7_75t_R g7500 ( 
.A(n_7491),
.Y(n_7500)
);

INVx2_ASAP7_75t_L g7501 ( 
.A(n_7495),
.Y(n_7501)
);

AOI22xp33_ASAP7_75t_L g7502 ( 
.A1(n_7496),
.A2(n_7486),
.B1(n_1607),
.B2(n_1605),
.Y(n_7502)
);

INVx2_ASAP7_75t_L g7503 ( 
.A(n_7498),
.Y(n_7503)
);

OAI22xp5_ASAP7_75t_L g7504 ( 
.A1(n_7500),
.A2(n_7497),
.B1(n_7492),
.B2(n_1610),
.Y(n_7504)
);

AOI21xp5_ASAP7_75t_L g7505 ( 
.A1(n_7501),
.A2(n_1606),
.B(n_1609),
.Y(n_7505)
);

INVxp67_ASAP7_75t_SL g7506 ( 
.A(n_7499),
.Y(n_7506)
);

OAI22xp5_ASAP7_75t_SL g7507 ( 
.A1(n_7503),
.A2(n_7502),
.B1(n_1611),
.B2(n_1609),
.Y(n_7507)
);

OAI22xp33_ASAP7_75t_L g7508 ( 
.A1(n_7506),
.A2(n_1612),
.B1(n_1610),
.B2(n_1611),
.Y(n_7508)
);

OAI21xp5_ASAP7_75t_L g7509 ( 
.A1(n_7505),
.A2(n_1613),
.B(n_1614),
.Y(n_7509)
);

OAI21xp5_ASAP7_75t_L g7510 ( 
.A1(n_7509),
.A2(n_7504),
.B(n_1613),
.Y(n_7510)
);

NAND2xp5_ASAP7_75t_L g7511 ( 
.A(n_7507),
.B(n_1614),
.Y(n_7511)
);

AOI22xp5_ASAP7_75t_L g7512 ( 
.A1(n_7511),
.A2(n_7508),
.B1(n_1617),
.B2(n_1615),
.Y(n_7512)
);

OAI21xp5_ASAP7_75t_L g7513 ( 
.A1(n_7512),
.A2(n_7510),
.B(n_1615),
.Y(n_7513)
);

AOI22xp5_ASAP7_75t_SL g7514 ( 
.A1(n_7513),
.A2(n_1621),
.B1(n_1616),
.B2(n_1620),
.Y(n_7514)
);

AOI221xp5_ASAP7_75t_L g7515 ( 
.A1(n_7514),
.A2(n_1622),
.B1(n_1616),
.B2(n_1620),
.C(n_1623),
.Y(n_7515)
);

AOI21xp5_ASAP7_75t_L g7516 ( 
.A1(n_7515),
.A2(n_1622),
.B(n_1623),
.Y(n_7516)
);

AOI211xp5_ASAP7_75t_L g7517 ( 
.A1(n_7516),
.A2(n_1626),
.B(n_1624),
.C(n_1625),
.Y(n_7517)
);


endmodule