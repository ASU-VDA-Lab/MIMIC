module fake_ariane_3041_n_2155 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2155);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2155;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_212;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_2144;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_2012;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_94),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_68),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_51),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_82),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_156),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_57),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_63),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_98),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_85),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_127),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_38),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_151),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_87),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_153),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_22),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_50),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_171),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_120),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_110),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_73),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_89),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_70),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_63),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_6),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_144),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_56),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_25),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_49),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_146),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_66),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_33),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_70),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_49),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_167),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_87),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_58),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_60),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_162),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_125),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_56),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_61),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_31),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_62),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_89),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_186),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_72),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_21),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_16),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_81),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_31),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_173),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_150),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_27),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_52),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_191),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_184),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_179),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_177),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_138),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_152),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_12),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_17),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_136),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_75),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_90),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_41),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_29),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_113),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_126),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_42),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_26),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_28),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_35),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_36),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_111),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_59),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_148),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_105),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_165),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_32),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_172),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_161),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_37),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_65),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_4),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_39),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_83),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_52),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_195),
.Y(n_303)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_166),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_44),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_160),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_142),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_96),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_79),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_72),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_2),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_164),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_88),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_77),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_149),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_28),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_180),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_115),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_88),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_73),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_145),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_51),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_60),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_155),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_39),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_108),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_130),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_104),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_83),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_68),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_75),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_64),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_76),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_66),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_57),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_78),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_188),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_169),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_13),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_178),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_62),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_45),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_42),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_189),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_24),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_45),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_54),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_14),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_124),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_23),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_194),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_106),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_118),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_35),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_78),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_196),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_141),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_32),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_64),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_119),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_100),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_69),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_34),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_4),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_91),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_80),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_117),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_183),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_27),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_1),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_46),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_114),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_95),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_17),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_12),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_157),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_103),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_55),
.Y(n_382)
);

BUFx8_ASAP7_75t_SL g383 ( 
.A(n_8),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_3),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_71),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_97),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_30),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_182),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_112),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g390 ( 
.A(n_67),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_53),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_132),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_251),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_383),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_203),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_257),
.B(n_0),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_235),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_235),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_235),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_208),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_235),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_208),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_219),
.B(n_0),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_235),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_235),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g406 ( 
.A(n_251),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_235),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_254),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_305),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_296),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_235),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_336),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_235),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_359),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_375),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_235),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_200),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_200),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_280),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_280),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_305),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_201),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_205),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_216),
.Y(n_424)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_257),
.B(n_3),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_205),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_207),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_206),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_202),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_204),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_210),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_212),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_257),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_245),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_206),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_214),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_228),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_258),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_233),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_233),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_281),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_261),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_261),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_326),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_309),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_231),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_309),
.Y(n_447)
);

INVxp33_ASAP7_75t_SL g448 ( 
.A(n_223),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_223),
.B(n_219),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_232),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_224),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_321),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_321),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_L g454 ( 
.A(n_224),
.B(n_5),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_324),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_234),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_324),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_237),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_207),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_268),
.B(n_7),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_364),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_358),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_238),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_243),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_377),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_244),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_246),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_249),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_218),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_L g473 ( 
.A(n_224),
.B(n_7),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_268),
.B(n_8),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_256),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_263),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_379),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_387),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_388),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_225),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_363),
.B(n_10),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_225),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_225),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_270),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_363),
.B(n_10),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_250),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_218),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g490 ( 
.A(n_288),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_226),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_226),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_395),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_423),
.B(n_217),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_370),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_423),
.B(n_370),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_448),
.B(n_227),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_433),
.B(n_217),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_424),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_408),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g505 ( 
.A1(n_488),
.A2(n_278),
.B(n_230),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_410),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_405),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_217),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_488),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_398),
.Y(n_510)
);

CKINVDCx8_ASAP7_75t_R g511 ( 
.A(n_394),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_398),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_R g513 ( 
.A(n_429),
.B(n_197),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_399),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_434),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_438),
.B(n_390),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_414),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_426),
.B(n_229),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_415),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_430),
.Y(n_521)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_401),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_431),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_401),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_404),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_432),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_436),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_407),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_411),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_426),
.B(n_227),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_411),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_413),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_437),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_419),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_416),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_446),
.B(n_463),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_393),
.B(n_259),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_416),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_R g543 ( 
.A(n_420),
.B(n_271),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_468),
.B(n_227),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_409),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_482),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_428),
.B(n_230),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_428),
.B(n_435),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_435),
.B(n_229),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_409),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_482),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_484),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_403),
.B(n_250),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_465),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_484),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_485),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_485),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_467),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_439),
.B(n_440),
.Y(n_560)
);

NAND2x1_ASAP7_75t_L g561 ( 
.A(n_440),
.B(n_230),
.Y(n_561)
);

NOR2x1_ASAP7_75t_L g562 ( 
.A(n_442),
.B(n_198),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_469),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_476),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_477),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_451),
.B(n_199),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_442),
.B(n_229),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_443),
.B(n_240),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_513),
.B(n_490),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_548),
.B(n_490),
.Y(n_575)
);

NAND3x1_ASAP7_75t_L g576 ( 
.A(n_497),
.B(n_483),
.C(n_403),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_529),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_548),
.B(n_451),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_501),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_529),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_529),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_494),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_531),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_493),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_548),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_525),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_541),
.B(n_393),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_531),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_534),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_497),
.A2(n_460),
.B1(n_487),
.B2(n_474),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_534),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_544),
.B(n_486),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_544),
.B(n_445),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_500),
.B(n_445),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_501),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_500),
.A2(n_406),
.B1(n_483),
.B2(n_421),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_503),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_539),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_504),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_525),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_539),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_555),
.B(n_447),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_501),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_539),
.Y(n_606)
);

AND2x6_ASAP7_75t_L g607 ( 
.A(n_570),
.B(n_278),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_546),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_513),
.B(n_421),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_540),
.B(n_450),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_546),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_L g612 ( 
.A1(n_541),
.A2(n_402),
.B1(n_400),
.B2(n_307),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_560),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_571),
.B(n_456),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_541),
.B(n_400),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_518),
.B(n_492),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_546),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_496),
.B(n_417),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_553),
.A2(n_402),
.B1(n_425),
.B2(n_396),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_546),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_545),
.B(n_458),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_546),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_568),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_571),
.B(n_412),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_555),
.B(n_447),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_553),
.A2(n_425),
.B1(n_396),
.B2(n_454),
.Y(n_626)
);

AND2x6_ASAP7_75t_L g627 ( 
.A(n_570),
.B(n_278),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_555),
.B(n_452),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_568),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_557),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_540),
.B(n_452),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_557),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_518),
.B(n_492),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_568),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_567),
.B(n_453),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_521),
.B(n_453),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_567),
.B(n_455),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_514),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_514),
.B(n_522),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_514),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_498),
.B(n_455),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_557),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_522),
.B(n_457),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_568),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_494),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_557),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_506),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_457),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_502),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_522),
.B(n_461),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_524),
.B(n_250),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_494),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_557),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_527),
.B(n_461),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_495),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_557),
.Y(n_657)
);

AND2x6_ASAP7_75t_L g658 ( 
.A(n_496),
.B(n_286),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_494),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_545),
.A2(n_307),
.B1(n_322),
.B2(n_259),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_557),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_558),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_496),
.B(n_286),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_550),
.B(n_464),
.Y(n_664)
);

AND2x6_ASAP7_75t_L g665 ( 
.A(n_496),
.B(n_286),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_558),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_495),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_560),
.B(n_464),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_558),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_537),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_525),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_550),
.A2(n_337),
.B1(n_335),
.B2(n_322),
.Y(n_673)
);

AND2x2_ASAP7_75t_SL g674 ( 
.A(n_505),
.B(n_360),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_537),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_518),
.B(n_417),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_537),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_533),
.B(n_466),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_510),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_525),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_533),
.B(n_466),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_558),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_563),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_502),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_563),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_563),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_496),
.B(n_471),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_563),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_528),
.A2(n_337),
.B1(n_335),
.B2(n_283),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_502),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_563),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_549),
.B(n_360),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_549),
.B(n_360),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_563),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_551),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_508),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_551),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_536),
.B(n_471),
.Y(n_701)
);

BUFx6f_ASAP7_75t_L g702 ( 
.A(n_494),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_525),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_525),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_552),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_549),
.B(n_418),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_503),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_525),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_572),
.B(n_418),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_494),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_552),
.Y(n_711)
);

INVx4_ASAP7_75t_SL g712 ( 
.A(n_547),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_554),
.B(n_472),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_499),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_562),
.A2(n_473),
.B1(n_454),
.B2(n_472),
.Y(n_715)
);

BUFx4f_ASAP7_75t_L g716 ( 
.A(n_547),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_R g717 ( 
.A(n_493),
.B(n_441),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_515),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_562),
.A2(n_473),
.B1(n_480),
.B2(n_475),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_556),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_569),
.B(n_475),
.Y(n_721)
);

INVx4_ASAP7_75t_SL g722 ( 
.A(n_547),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_499),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_499),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_499),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_695),
.A2(n_481),
.B1(n_480),
.B2(n_547),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_615),
.B(n_517),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_613),
.B(n_642),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_698),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_649),
.B(n_559),
.Y(n_730)
);

NAND2x1_ASAP7_75t_L g731 ( 
.A(n_695),
.B(n_510),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_594),
.B(n_564),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_698),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_596),
.B(n_593),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_700),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_700),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_591),
.B(n_565),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_705),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_601),
.B(n_561),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_705),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_625),
.B(n_566),
.Y(n_741)
);

BUFx5_ASAP7_75t_L g742 ( 
.A(n_674),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_576),
.A2(n_252),
.B1(n_308),
.B2(n_226),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_674),
.A2(n_640),
.B(n_611),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_656),
.B(n_512),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_615),
.B(n_519),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_711),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_650),
.B(n_508),
.Y(n_748)
);

AND2x2_ASAP7_75t_SL g749 ( 
.A(n_674),
.B(n_371),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_650),
.B(n_508),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_711),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_583),
.Y(n_752)
);

HB1xp67_ASAP7_75t_L g753 ( 
.A(n_599),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_695),
.A2(n_481),
.B1(n_547),
.B2(n_505),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_720),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_585),
.B(n_511),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_576),
.A2(n_543),
.B1(n_561),
.B2(n_569),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_591),
.B(n_512),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_686),
.B(n_523),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_686),
.B(n_569),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_693),
.B(n_572),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_693),
.B(n_699),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_699),
.B(n_586),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_586),
.B(n_572),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_656),
.B(n_523),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_720),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_637),
.B(n_526),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_656),
.B(n_526),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_671),
.B(n_511),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_678),
.B(n_530),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_683),
.B(n_530),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_671),
.B(n_675),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_618),
.B(n_511),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_706),
.B(n_709),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_618),
.B(n_275),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_583),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_706),
.B(n_532),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_655),
.B(n_532),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_675),
.B(n_427),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_695),
.A2(n_547),
.B1(n_505),
.B2(n_556),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_585),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_608),
.Y(n_782)
);

NAND2x1p5_ASAP7_75t_L g783 ( 
.A(n_716),
.B(n_505),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_714),
.A2(n_538),
.B(n_535),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_721),
.A2(n_538),
.B(n_542),
.C(n_535),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_575),
.A2(n_543),
.B1(n_380),
.B2(n_542),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_639),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_706),
.B(n_499),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_706),
.B(n_499),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_695),
.A2(n_547),
.B1(n_505),
.B2(n_459),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_639),
.Y(n_791)
);

OR2x6_ASAP7_75t_L g792 ( 
.A(n_677),
.B(n_427),
.Y(n_792)
);

INVx3_ASAP7_75t_L g793 ( 
.A(n_639),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_701),
.B(n_459),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_664),
.A2(n_252),
.B(n_362),
.C(n_308),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_709),
.B(n_499),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_695),
.A2(n_547),
.B1(n_489),
.B2(n_470),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_608),
.A2(n_252),
.B(n_362),
.C(n_308),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_611),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_709),
.B(n_507),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_589),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_573),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_714),
.A2(n_507),
.B(n_489),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_R g804 ( 
.A(n_677),
.B(n_516),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_713),
.B(n_470),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_618),
.B(n_575),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_617),
.A2(n_362),
.B(n_348),
.C(n_240),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_709),
.B(n_507),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_668),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_618),
.B(n_507),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_716),
.B(n_371),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_676),
.B(n_507),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_616),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_616),
.B(n_220),
.Y(n_814)
);

NOR3xp33_ASAP7_75t_L g815 ( 
.A(n_614),
.B(n_239),
.C(n_220),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_617),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_648),
.B(n_516),
.Y(n_817)
);

AND2x6_ASAP7_75t_SL g818 ( 
.A(n_624),
.B(n_239),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_634),
.B(n_241),
.Y(n_819)
);

O2A1O1Ixp33_ASAP7_75t_L g820 ( 
.A1(n_689),
.A2(n_253),
.B(n_255),
.C(n_241),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_632),
.B(n_507),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_676),
.B(n_507),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_669),
.B(n_547),
.Y(n_824)
);

NOR2xp67_ASAP7_75t_L g825 ( 
.A(n_574),
.B(n_209),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_604),
.A2(n_273),
.B(n_319),
.C(n_385),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_578),
.B(n_547),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_668),
.B(n_371),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_620),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_695),
.A2(n_696),
.B1(n_658),
.B2(n_665),
.Y(n_830)
);

AOI22xp33_ASAP7_75t_L g831 ( 
.A1(n_696),
.A2(n_289),
.B1(n_317),
.B2(n_338),
.Y(n_831)
);

AND2x6_ASAP7_75t_SL g832 ( 
.A(n_717),
.B(n_253),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_589),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_573),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_592),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_718),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_622),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_588),
.B(n_516),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_609),
.B(n_285),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_578),
.B(n_380),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_634),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_636),
.B(n_240),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_696),
.A2(n_291),
.B1(n_339),
.B2(n_255),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_621),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_622),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_668),
.B(n_264),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_579),
.B(n_287),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_696),
.A2(n_291),
.B1(n_338),
.B2(n_262),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_579),
.B(n_294),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_579),
.B(n_250),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_648),
.B(n_298),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_679),
.Y(n_852)
);

NOR2x1p5_ASAP7_75t_L g853 ( 
.A(n_588),
.B(n_348),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_598),
.A2(n_325),
.B1(n_300),
.B2(n_312),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_691),
.A2(n_479),
.B1(n_478),
.B2(n_462),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_638),
.B(n_619),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_696),
.A2(n_347),
.B1(n_272),
.B2(n_269),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_696),
.A2(n_339),
.B1(n_262),
.B2(n_273),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_623),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_592),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_679),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_623),
.A2(n_276),
.B(n_274),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_600),
.Y(n_863)
);

INVx5_ASAP7_75t_L g864 ( 
.A(n_658),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_628),
.B(n_348),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_629),
.B(n_274),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_597),
.B(n_313),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_612),
.B(n_314),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_696),
.A2(n_344),
.B1(n_276),
.B2(n_361),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_679),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_629),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_630),
.B(n_289),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_630),
.B(n_635),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_573),
.B(n_582),
.Y(n_874)
);

INVx8_ASAP7_75t_L g875 ( 
.A(n_658),
.Y(n_875)
);

NOR2xp67_ASAP7_75t_L g876 ( 
.A(n_621),
.B(n_610),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_658),
.A2(n_665),
.B1(n_663),
.B2(n_627),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_635),
.B(n_290),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_645),
.B(n_290),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_645),
.B(n_297),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_660),
.B(n_515),
.Y(n_881)
);

INVx1_ASAP7_75t_SL g882 ( 
.A(n_707),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_644),
.B(n_297),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_SL g884 ( 
.A1(n_673),
.A2(n_444),
.B1(n_626),
.B2(n_323),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_577),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_597),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_573),
.Y(n_887)
);

AOI22xp5_ASAP7_75t_L g888 ( 
.A1(n_658),
.A2(n_221),
.B1(n_222),
.B2(n_392),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_573),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_658),
.A2(n_215),
.B1(n_211),
.B2(n_389),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_597),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_651),
.B(n_605),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_605),
.B(n_299),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_605),
.B(n_641),
.Y(n_894)
);

NAND2x1_ASAP7_75t_L g895 ( 
.A(n_658),
.B(n_509),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_641),
.B(n_299),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_641),
.A2(n_332),
.B1(n_391),
.B2(n_334),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_729),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_875),
.Y(n_899)
);

BUFx4f_ASAP7_75t_L g900 ( 
.A(n_875),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_779),
.B(n_715),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_806),
.B(n_712),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_875),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_774),
.B(n_712),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_864),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_752),
.Y(n_906)
);

OR2x2_ASAP7_75t_SL g907 ( 
.A(n_730),
.B(n_302),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_752),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_802),
.Y(n_909)
);

INVx5_ASAP7_75t_L g910 ( 
.A(n_864),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_SL g911 ( 
.A(n_781),
.B(n_328),
.C(n_316),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_737),
.A2(n_665),
.B1(n_663),
.B2(n_627),
.Y(n_912)
);

BUFx2_ASAP7_75t_SL g913 ( 
.A(n_864),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_836),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_734),
.B(n_663),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_SL g916 ( 
.A(n_737),
.B(n_342),
.C(n_333),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_787),
.Y(n_917)
);

INVxp33_ASAP7_75t_SL g918 ( 
.A(n_756),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_728),
.B(n_663),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_733),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_SL g921 ( 
.A(n_756),
.B(n_346),
.C(n_345),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_735),
.Y(n_922)
);

INVxp67_ASAP7_75t_SL g923 ( 
.A(n_809),
.Y(n_923)
);

INVxp67_ASAP7_75t_SL g924 ( 
.A(n_809),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_758),
.B(n_663),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_R g926 ( 
.A(n_804),
.B(n_769),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_787),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_779),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_776),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_802),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_776),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_758),
.B(n_663),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_732),
.B(n_725),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_882),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_813),
.B(n_719),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_801),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_749),
.A2(n_708),
.B1(n_602),
.B2(n_672),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_874),
.A2(n_714),
.B(n_724),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_749),
.A2(n_665),
.B1(n_663),
.B2(n_627),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_801),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_833),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_SL g942 ( 
.A1(n_817),
.A2(n_665),
.B1(n_627),
.B2(n_607),
.Y(n_942)
);

BUFx10_ASAP7_75t_L g943 ( 
.A(n_839),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_741),
.B(n_665),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_874),
.A2(n_724),
.B(n_708),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_779),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_794),
.A2(n_805),
.B1(n_773),
.B2(n_841),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_736),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_738),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_884),
.A2(n_665),
.B1(n_627),
.B2(n_607),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_SL g951 ( 
.A(n_804),
.B(n_851),
.C(n_353),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_740),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_747),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_833),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_864),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_846),
.A2(n_580),
.B(n_577),
.Y(n_956)
);

AND2x6_ASAP7_75t_L g957 ( 
.A(n_830),
.B(n_861),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_861),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_840),
.B(n_748),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_835),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_751),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_750),
.B(n_580),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_794),
.B(n_581),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_805),
.B(n_581),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_763),
.B(n_584),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_802),
.Y(n_966)
);

BUFx2_ASAP7_75t_L g967 ( 
.A(n_792),
.Y(n_967)
);

BUFx4f_ASAP7_75t_L g968 ( 
.A(n_811),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_755),
.Y(n_969)
);

NOR2x1_ASAP7_75t_L g970 ( 
.A(n_727),
.B(n_587),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_870),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_764),
.B(n_584),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_870),
.B(n_582),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_767),
.B(n_590),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_R g975 ( 
.A(n_746),
.B(n_652),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_786),
.B(n_725),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_766),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_767),
.A2(n_778),
.B(n_759),
.C(n_757),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_742),
.B(n_852),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_739),
.B(n_712),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_835),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_885),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_778),
.B(n_590),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_742),
.B(n_582),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_860),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_760),
.B(n_595),
.Y(n_986)
);

NAND2xp33_ASAP7_75t_R g987 ( 
.A(n_838),
.B(n_661),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_782),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_844),
.B(n_587),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_860),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_792),
.B(n_595),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_761),
.B(n_606),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_799),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_816),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_863),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_759),
.B(n_606),
.Y(n_996)
);

BUFx4f_ASAP7_75t_L g997 ( 
.A(n_811),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_739),
.Y(n_998)
);

OR2x6_ASAP7_75t_SL g999 ( 
.A(n_854),
.B(n_351),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_802),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_792),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_772),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_838),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_762),
.B(n_600),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_SL g1005 ( 
.A(n_897),
.B(n_367),
.C(n_365),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_753),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_742),
.B(n_582),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_838),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_777),
.B(n_603),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_822),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_834),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_742),
.A2(n_627),
.B1(n_607),
.B2(n_672),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_863),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_895),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_834),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_886),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_829),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_834),
.Y(n_1018)
);

NAND2xp33_ASAP7_75t_SL g1019 ( 
.A(n_731),
.B(n_587),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_834),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_R g1021 ( 
.A(n_881),
.B(n_716),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_876),
.Y(n_1022)
);

INVx3_ASAP7_75t_L g1023 ( 
.A(n_886),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_887),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_837),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_832),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_742),
.B(n_725),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_887),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_814),
.B(n_603),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_812),
.B(n_607),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_845),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_823),
.B(n_607),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_852),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_742),
.B(n_582),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_818),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_770),
.B(n_607),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_859),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_771),
.B(n_607),
.Y(n_1038)
);

INVx3_ASAP7_75t_L g1039 ( 
.A(n_887),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_871),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_855),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_788),
.B(n_627),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_810),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_839),
.B(n_587),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_814),
.Y(n_1045)
);

BUFx4f_ASAP7_75t_L g1046 ( 
.A(n_739),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_789),
.B(n_708),
.Y(n_1047)
);

NOR2xp67_ASAP7_75t_L g1048 ( 
.A(n_825),
.B(n_661),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_891),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_894),
.A2(n_724),
.B(n_672),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_877),
.B(n_725),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_R g1052 ( 
.A(n_791),
.B(n_661),
.Y(n_1052)
);

AND3x1_ASAP7_75t_SL g1053 ( 
.A(n_853),
.B(n_317),
.C(n_302),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_796),
.B(n_602),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_887),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_891),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_873),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_800),
.B(n_808),
.Y(n_1058)
);

AO22x1_ASAP7_75t_L g1059 ( 
.A1(n_743),
.A2(n_319),
.B1(n_344),
.B2(n_349),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_889),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_819),
.B(n_602),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_819),
.B(n_602),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_866),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_889),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_872),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_889),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_744),
.A2(n_662),
.B(n_657),
.Y(n_1067)
);

NOR2x2_ASAP7_75t_L g1068 ( 
.A(n_815),
.B(n_631),
.Y(n_1068)
);

INVx4_ASAP7_75t_L g1069 ( 
.A(n_889),
.Y(n_1069)
);

BUFx8_ASAP7_75t_L g1070 ( 
.A(n_831),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_791),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_847),
.B(n_672),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_847),
.B(n_680),
.Y(n_1073)
);

AND2x2_ASAP7_75t_SL g1074 ( 
.A(n_877),
.B(n_250),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_793),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_775),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_793),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_827),
.Y(n_1078)
);

AND3x1_ASAP7_75t_SL g1079 ( 
.A(n_868),
.B(n_350),
.C(n_349),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_783),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_SL g1081 ( 
.A(n_797),
.B(n_725),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_849),
.B(n_680),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_824),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_849),
.B(n_680),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_783),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_797),
.B(n_712),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_878),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_883),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_867),
.B(n_682),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_892),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_831),
.A2(n_647),
.B1(n_684),
.B2(n_670),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1072),
.A2(n_850),
.B(n_784),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_959),
.B(n_1088),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_998),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_SL g1095 ( 
.A(n_918),
.B(n_1070),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_1074),
.B(n_1029),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_922),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_906),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_978),
.B(n_867),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_915),
.A2(n_919),
.B(n_1036),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_1002),
.B(n_893),
.Y(n_1101)
);

OAI21xp33_ASAP7_75t_SL g1102 ( 
.A1(n_1074),
.A2(n_848),
.B(n_843),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_906),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_908),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_910),
.B(n_745),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1073),
.A2(n_765),
.B(n_745),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1082),
.A2(n_768),
.B(n_765),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1038),
.A2(n_803),
.B(n_768),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_SL g1109 ( 
.A1(n_1017),
.A2(n_932),
.B(n_925),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_952),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_968),
.B(n_862),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_968),
.A2(n_843),
.B1(n_858),
.B2(n_848),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1057),
.B(n_858),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_956),
.A2(n_785),
.B(n_846),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_968),
.A2(n_869),
.B1(n_790),
.B2(n_857),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_956),
.A2(n_828),
.B(n_879),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1061),
.A2(n_795),
.B(n_880),
.C(n_820),
.Y(n_1117)
);

A2O1A1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_1087),
.A2(n_869),
.B(n_826),
.C(n_856),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1087),
.A2(n_896),
.B(n_821),
.C(n_726),
.Y(n_1119)
);

INVx6_ASAP7_75t_SL g1120 ( 
.A(n_980),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_961),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1084),
.A2(n_996),
.B(n_1044),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_1005),
.B(n_807),
.C(n_798),
.Y(n_1123)
);

INVx4_ASAP7_75t_SL g1124 ( 
.A(n_957),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_908),
.Y(n_1125)
);

BUFx2_ASAP7_75t_SL g1126 ( 
.A(n_934),
.Y(n_1126)
);

HB1xp67_ASAP7_75t_L g1127 ( 
.A(n_928),
.Y(n_1127)
);

NOR2x1_ASAP7_75t_SL g1128 ( 
.A(n_913),
.B(n_828),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_903),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_934),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_1006),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1067),
.A2(n_780),
.B(n_723),
.Y(n_1132)
);

AOI21xp33_ASAP7_75t_L g1133 ( 
.A1(n_1070),
.A2(n_821),
.B(n_888),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1085),
.A2(n_780),
.B(n_723),
.Y(n_1134)
);

O2A1O1Ixp5_ASAP7_75t_L g1135 ( 
.A1(n_933),
.A2(n_865),
.B(n_842),
.C(n_724),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1085),
.A2(n_710),
.A3(n_631),
.B(n_633),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_946),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_912),
.A2(n_726),
.B(n_790),
.C(n_369),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_997),
.A2(n_890),
.B1(n_754),
.B2(n_682),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1029),
.B(n_754),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1070),
.A2(n_288),
.B1(n_385),
.B2(n_361),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_944),
.A2(n_703),
.B(n_680),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_938),
.A2(n_710),
.B(n_643),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1050),
.A2(n_643),
.B(n_633),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_945),
.A2(n_654),
.B(n_647),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_974),
.A2(n_704),
.B(n_703),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_984),
.A2(n_1027),
.B(n_1007),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_997),
.A2(n_682),
.B1(n_704),
.B2(n_703),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_991),
.B(n_722),
.Y(n_1149)
);

INVx3_ASAP7_75t_SL g1150 ( 
.A(n_1076),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1030),
.A2(n_662),
.B(n_657),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_991),
.B(n_722),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_983),
.A2(n_704),
.B(n_703),
.Y(n_1153)
);

AOI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_681),
.B(n_666),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1057),
.B(n_704),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_SL g1156 ( 
.A1(n_899),
.A2(n_939),
.B(n_903),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1034),
.A2(n_667),
.B(n_654),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_1017),
.A2(n_670),
.B(n_667),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_980),
.B(n_722),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_947),
.B(n_1043),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1090),
.A2(n_692),
.B(n_684),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1090),
.A2(n_692),
.B(n_681),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1032),
.A2(n_685),
.B(n_666),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1090),
.A2(n_687),
.B(n_685),
.Y(n_1164)
);

INVx4_ASAP7_75t_SL g1165 ( 
.A(n_957),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1054),
.A2(n_688),
.B(n_687),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1058),
.A2(n_690),
.B(n_688),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_946),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1002),
.B(n_722),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1078),
.A2(n_694),
.B(n_690),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1083),
.A2(n_697),
.A3(n_694),
.B(n_369),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_979),
.A2(n_697),
.B(n_357),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1083),
.A2(n_357),
.A3(n_350),
.B(n_378),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_962),
.A2(n_653),
.B(n_646),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_972),
.A2(n_653),
.B(n_646),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_898),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1043),
.B(n_646),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_976),
.A2(n_382),
.B(n_378),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_918),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_998),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_997),
.B(n_382),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_929),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1063),
.B(n_646),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_986),
.A2(n_702),
.B(n_659),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_898),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_929),
.A2(n_315),
.B(n_213),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_SL g1187 ( 
.A(n_913),
.B(n_646),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_920),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1065),
.B(n_653),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_914),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_SL g1191 ( 
.A1(n_1069),
.A2(n_13),
.B(n_14),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1051),
.A2(n_702),
.B(n_659),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_920),
.B(n_288),
.Y(n_1193)
);

BUFx4_ASAP7_75t_SL g1194 ( 
.A(n_967),
.Y(n_1194)
);

AOI31xp67_ASAP7_75t_L g1195 ( 
.A1(n_1060),
.A2(n_702),
.A3(n_659),
.B(n_653),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_935),
.B(n_948),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_903),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_948),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_SL g1199 ( 
.A(n_910),
.B(n_653),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_949),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_SL g1201 ( 
.A1(n_1069),
.A2(n_15),
.B(n_18),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_901),
.B(n_659),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1078),
.A2(n_1047),
.B(n_1042),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_949),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_L g1205 ( 
.A1(n_975),
.A2(n_374),
.B(n_368),
.Y(n_1205)
);

AND2x6_ASAP7_75t_SL g1206 ( 
.A(n_1035),
.B(n_372),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_980),
.B(n_659),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1014),
.A2(n_702),
.B(n_520),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_935),
.B(n_702),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_953),
.B(n_373),
.Y(n_1210)
);

O2A1O1Ixp5_ASAP7_75t_L g1211 ( 
.A1(n_973),
.A2(n_250),
.B(n_282),
.C(n_284),
.Y(n_1211)
);

AO21x2_ASAP7_75t_L g1212 ( 
.A1(n_1081),
.A2(n_964),
.B(n_963),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_931),
.A2(n_520),
.A3(n_509),
.B(n_288),
.Y(n_1213)
);

BUFx2_ASAP7_75t_SL g1214 ( 
.A(n_967),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_953),
.B(n_384),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_992),
.A2(n_310),
.B(n_236),
.Y(n_1216)
);

NAND2x1_ASAP7_75t_L g1217 ( 
.A(n_899),
.B(n_509),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1048),
.A2(n_520),
.B(n_509),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_969),
.B(n_15),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_969),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1001),
.Y(n_1221)
);

BUFx4_ASAP7_75t_SL g1222 ( 
.A(n_1001),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_977),
.A2(n_198),
.B(n_311),
.C(n_266),
.Y(n_1223)
);

AO32x2_ASAP7_75t_L g1224 ( 
.A1(n_937),
.A2(n_520),
.A3(n_509),
.B1(n_366),
.B2(n_301),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1004),
.A2(n_520),
.B(n_509),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_977),
.B(n_18),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_965),
.A2(n_520),
.B(n_509),
.Y(n_1227)
);

AO22x2_ASAP7_75t_L g1228 ( 
.A1(n_901),
.A2(n_266),
.B1(n_198),
.B2(n_311),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1009),
.A2(n_306),
.B(n_386),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1086),
.B(n_266),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1045),
.B(n_19),
.Y(n_1231)
);

AOI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1076),
.A2(n_242),
.B1(n_376),
.B2(n_260),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1014),
.A2(n_520),
.B(n_304),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1014),
.A2(n_304),
.B(n_311),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_943),
.B(n_19),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_SL g1236 ( 
.A1(n_1069),
.A2(n_20),
.B(n_21),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_931),
.A2(n_304),
.B(n_264),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_943),
.B(n_20),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_916),
.B(n_366),
.C(n_282),
.Y(n_1239)
);

OR2x2_ASAP7_75t_L g1240 ( 
.A(n_1008),
.B(n_22),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_903),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_900),
.A2(n_303),
.B(n_356),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_936),
.A2(n_304),
.B(n_264),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_SL g1244 ( 
.A(n_911),
.B(n_247),
.C(n_248),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_900),
.A2(n_318),
.B(n_265),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_900),
.A2(n_320),
.B(n_267),
.Y(n_1246)
);

OA21x2_ASAP7_75t_L g1247 ( 
.A1(n_936),
.A2(n_327),
.B(n_277),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_899),
.B(n_99),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_943),
.B(n_23),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_940),
.A2(n_304),
.B(n_264),
.Y(n_1250)
);

AO21x2_ASAP7_75t_L g1251 ( 
.A1(n_1089),
.A2(n_304),
.B(n_264),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_982),
.B(n_24),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_940),
.A2(n_304),
.B(n_264),
.Y(n_1253)
);

BUFx8_ASAP7_75t_SL g1254 ( 
.A(n_1035),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_994),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_941),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_SL g1257 ( 
.A1(n_1049),
.A2(n_25),
.B(n_26),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_988),
.A2(n_279),
.B(n_292),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1112),
.A2(n_1086),
.B1(n_999),
.B2(n_907),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1228),
.A2(n_926),
.B1(n_1086),
.B2(n_1003),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_SL g1261 ( 
.A1(n_1109),
.A2(n_1012),
.B(n_982),
.Y(n_1261)
);

AOI221xp5_ASAP7_75t_L g1262 ( 
.A1(n_1102),
.A2(n_1059),
.B1(n_921),
.B2(n_951),
.C(n_1037),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1098),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1099),
.A2(n_999),
.B1(n_907),
.B2(n_989),
.Y(n_1264)
);

OA21x2_ASAP7_75t_L g1265 ( 
.A1(n_1237),
.A2(n_954),
.B(n_941),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1122),
.A2(n_970),
.B(n_1062),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1098),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1094),
.B(n_910),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1228),
.A2(n_1003),
.B1(n_1021),
.B2(n_950),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1095),
.B(n_998),
.Y(n_1270)
);

AOI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1225),
.A2(n_993),
.B(n_988),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1097),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1119),
.A2(n_990),
.A3(n_1013),
.B(n_985),
.Y(n_1273)
);

AO21x2_ASAP7_75t_L g1274 ( 
.A1(n_1227),
.A2(n_1010),
.B(n_993),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1093),
.B(n_1046),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1126),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1237),
.A2(n_960),
.B(n_954),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1130),
.B(n_1026),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1243),
.A2(n_981),
.B(n_960),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1103),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1254),
.Y(n_1281)
);

OAI21xp33_ASAP7_75t_SL g1282 ( 
.A1(n_1111),
.A2(n_1216),
.B(n_1235),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1196),
.B(n_1059),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1115),
.A2(n_1010),
.B1(n_1025),
.B2(n_1031),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1181),
.B(n_1025),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1160),
.B(n_1031),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1218),
.A2(n_1144),
.B(n_1092),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1103),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1104),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1243),
.A2(n_985),
.B(n_981),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1111),
.A2(n_1071),
.B(n_1040),
.C(n_1023),
.Y(n_1291)
);

AO222x2_ASAP7_75t_L g1292 ( 
.A1(n_1181),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.C1(n_36),
.C2(n_37),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1104),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1125),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1140),
.B(n_1040),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1138),
.A2(n_1033),
.B1(n_1046),
.B2(n_1016),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1096),
.B(n_1033),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1125),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1140),
.B(n_1046),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1096),
.B(n_1080),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1101),
.B(n_1137),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1182),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1230),
.B(n_958),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1101),
.B(n_958),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1250),
.A2(n_1013),
.B(n_995),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1207),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1119),
.A2(n_990),
.A3(n_995),
.B(n_1064),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1256),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1250),
.A2(n_1028),
.B(n_1039),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1253),
.A2(n_1049),
.B(n_1056),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1219),
.A2(n_1071),
.B(n_1023),
.C(n_971),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1106),
.A2(n_923),
.B(n_924),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1230),
.B(n_1056),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1256),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_SL g1316 ( 
.A1(n_1226),
.A2(n_1023),
.B(n_971),
.C(n_1077),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1228),
.A2(n_1022),
.B1(n_1026),
.B2(n_902),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1131),
.B(n_917),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1248),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1253),
.A2(n_1144),
.B(n_1233),
.Y(n_1320)
);

OA21x2_ASAP7_75t_L g1321 ( 
.A1(n_1114),
.A2(n_1091),
.B(n_1060),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1168),
.Y(n_1322)
);

OR3x4_ASAP7_75t_SL g1323 ( 
.A(n_1254),
.B(n_1053),
.C(n_1079),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1110),
.Y(n_1324)
);

AOI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1141),
.A2(n_366),
.B1(n_301),
.B2(n_284),
.C(n_282),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1241),
.Y(n_1326)
);

INVx1_ASAP7_75t_SL g1327 ( 
.A(n_1150),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1141),
.A2(n_902),
.B1(n_957),
.B2(n_904),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1193),
.B(n_917),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1193),
.B(n_927),
.Y(n_1330)
);

CKINVDCx8_ASAP7_75t_R g1331 ( 
.A(n_1214),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1176),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1185),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1223),
.A2(n_1066),
.A3(n_1064),
.B(n_1075),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_1202),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1202),
.A2(n_987),
.B1(n_957),
.B2(n_902),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1150),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1121),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1233),
.A2(n_1028),
.B(n_1039),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1255),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1161),
.A2(n_1028),
.B(n_1039),
.Y(n_1341)
);

OAI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1138),
.A2(n_1016),
.B1(n_1075),
.B2(n_942),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1207),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1188),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1165),
.B(n_927),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1161),
.A2(n_1055),
.B(n_1066),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1192),
.A2(n_905),
.B(n_904),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1136),
.Y(n_1348)
);

INVx6_ASAP7_75t_L g1349 ( 
.A(n_1159),
.Y(n_1349)
);

AO21x2_ASAP7_75t_L g1350 ( 
.A1(n_1223),
.A2(n_1052),
.B(n_904),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1133),
.A2(n_957),
.B1(n_1080),
.B2(n_905),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_1194),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1177),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1143),
.A2(n_1055),
.B(n_1077),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1231),
.A2(n_1068),
.B1(n_910),
.B2(n_903),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1143),
.A2(n_1145),
.B(n_1192),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1145),
.A2(n_1055),
.B(n_1077),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1234),
.A2(n_955),
.B(n_1019),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1190),
.B(n_957),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1094),
.B(n_910),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1200),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1204),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1136),
.Y(n_1364)
);

AND2x6_ASAP7_75t_SL g1365 ( 
.A(n_1238),
.B(n_1068),
.Y(n_1365)
);

NAND2x1p5_ASAP7_75t_L g1366 ( 
.A(n_1180),
.B(n_909),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1234),
.A2(n_955),
.B(n_1019),
.Y(n_1367)
);

AOI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1114),
.A2(n_1024),
.B(n_1020),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1179),
.B(n_909),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1222),
.Y(n_1370)
);

BUFx4_ASAP7_75t_SL g1371 ( 
.A(n_1206),
.Y(n_1371)
);

AOI22x1_ASAP7_75t_L g1372 ( 
.A1(n_1107),
.A2(n_1024),
.B1(n_1020),
.B2(n_1018),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1220),
.Y(n_1373)
);

OA21x2_ASAP7_75t_L g1374 ( 
.A1(n_1116),
.A2(n_352),
.B(n_293),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1179),
.B(n_1024),
.Y(n_1375)
);

AOI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1174),
.A2(n_1024),
.B(n_1020),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1116),
.A2(n_354),
.B(n_295),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1162),
.A2(n_331),
.B(n_340),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1162),
.A2(n_1157),
.B(n_1164),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1159),
.Y(n_1380)
);

INVxp67_ASAP7_75t_L g1381 ( 
.A(n_1127),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1258),
.A2(n_1024),
.B1(n_1020),
.B2(n_1018),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1118),
.A2(n_955),
.B(n_1018),
.C(n_1015),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1157),
.A2(n_1020),
.B(n_1018),
.Y(n_1384)
);

OA21x2_ASAP7_75t_L g1385 ( 
.A1(n_1134),
.A2(n_330),
.B(n_341),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1136),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1164),
.A2(n_1018),
.B(n_1015),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1180),
.B(n_909),
.Y(n_1388)
);

INVx5_ASAP7_75t_L g1389 ( 
.A(n_1159),
.Y(n_1389)
);

CKINVDCx6p67_ASAP7_75t_R g1390 ( 
.A(n_1241),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1221),
.B(n_909),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1136),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1208),
.A2(n_1015),
.B(n_1011),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1175),
.A2(n_1015),
.B(n_1011),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1248),
.Y(n_1395)
);

OA21x2_ASAP7_75t_L g1396 ( 
.A1(n_1134),
.A2(n_343),
.B(n_329),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1124),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1167),
.A2(n_1015),
.B(n_1011),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1171),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1205),
.A2(n_1011),
.B1(n_1000),
.B2(n_966),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1113),
.A2(n_1011),
.B1(n_1000),
.B2(n_966),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1165),
.B(n_909),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1252),
.Y(n_1403)
);

INVx6_ASAP7_75t_L g1404 ( 
.A(n_1207),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1171),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1208),
.A2(n_1147),
.B(n_1135),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1240),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1241),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1147),
.A2(n_1000),
.B(n_966),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1118),
.A2(n_1249),
.B(n_1239),
.C(n_1117),
.Y(n_1410)
);

BUFx12f_ASAP7_75t_L g1411 ( 
.A(n_1240),
.Y(n_1411)
);

AND2x4_ASAP7_75t_L g1412 ( 
.A(n_1165),
.B(n_930),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1248),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1232),
.B(n_930),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1124),
.B(n_1149),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1169),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1124),
.B(n_930),
.Y(n_1417)
);

CKINVDCx14_ASAP7_75t_R g1418 ( 
.A(n_1244),
.Y(n_1418)
);

CKINVDCx8_ASAP7_75t_R g1419 ( 
.A(n_1124),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1149),
.B(n_930),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1169),
.B(n_930),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1241),
.B(n_1000),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1100),
.A2(n_1178),
.B(n_1132),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1178),
.A2(n_1132),
.B(n_1184),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1210),
.B(n_1000),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1215),
.B(n_1152),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1209),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1158),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1129),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1171),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1139),
.A2(n_966),
.B1(n_366),
.B2(n_301),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1264),
.A2(n_1123),
.B1(n_1189),
.B2(n_1183),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1259),
.A2(n_1186),
.B1(n_1247),
.B2(n_1201),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1407),
.B(n_1152),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1263),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1292),
.B(n_1120),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1272),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1319),
.A2(n_1156),
.B(n_1166),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1352),
.Y(n_1439)
);

OAI221xp5_ASAP7_75t_L g1440 ( 
.A1(n_1282),
.A2(n_1229),
.B1(n_1203),
.B2(n_1108),
.C(n_1246),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1281),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1285),
.B(n_1173),
.Y(n_1442)
);

INVx2_ASAP7_75t_SL g1443 ( 
.A(n_1370),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1418),
.A2(n_282),
.B1(n_301),
.B2(n_366),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1324),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1259),
.A2(n_1247),
.B1(n_1186),
.B2(n_1191),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1307),
.B(n_1241),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1419),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1319),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1304),
.B(n_1120),
.Y(n_1450)
);

CKINVDCx16_ASAP7_75t_R g1451 ( 
.A(n_1411),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1307),
.B(n_1129),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1331),
.Y(n_1453)
);

OAI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1262),
.A2(n_1242),
.B1(n_1245),
.B2(n_1170),
.C(n_1154),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1338),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1301),
.B(n_1173),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1322),
.Y(n_1457)
);

NAND3x1_ASAP7_75t_L g1458 ( 
.A(n_1278),
.B(n_1151),
.C(n_1163),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1397),
.B(n_1156),
.Y(n_1459)
);

OR2x6_ASAP7_75t_L g1460 ( 
.A(n_1397),
.B(n_1105),
.Y(n_1460)
);

AO31x2_ASAP7_75t_L g1461 ( 
.A1(n_1348),
.A2(n_1142),
.A3(n_1128),
.B(n_1153),
.Y(n_1461)
);

OR2x6_ASAP7_75t_L g1462 ( 
.A(n_1319),
.B(n_1105),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1331),
.Y(n_1463)
);

OAI221xp5_ASAP7_75t_L g1464 ( 
.A1(n_1410),
.A2(n_1155),
.B1(n_1211),
.B2(n_1247),
.C(n_1186),
.Y(n_1464)
);

NAND3xp33_ASAP7_75t_L g1465 ( 
.A(n_1403),
.B(n_282),
.C(n_284),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1340),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1395),
.A2(n_1187),
.B(n_1199),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1395),
.A2(n_1146),
.B(n_966),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1301),
.B(n_1173),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1395),
.A2(n_1148),
.B(n_1212),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1259),
.A2(n_1120),
.B1(n_1129),
.B2(n_1197),
.Y(n_1471)
);

NAND3xp33_ASAP7_75t_SL g1472 ( 
.A(n_1327),
.B(n_1236),
.C(n_1217),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1320),
.A2(n_1172),
.B(n_1257),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1373),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1259),
.A2(n_1251),
.B1(n_1212),
.B2(n_1224),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1260),
.A2(n_1212),
.B1(n_1251),
.B2(n_282),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1269),
.A2(n_1251),
.B1(n_284),
.B2(n_366),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1322),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1284),
.A2(n_284),
.B1(n_301),
.B2(n_355),
.C(n_1224),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1263),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1343),
.B(n_1129),
.Y(n_1481)
);

CKINVDCx16_ASAP7_75t_R g1482 ( 
.A(n_1411),
.Y(n_1482)
);

NAND2x1_ASAP7_75t_L g1483 ( 
.A(n_1413),
.B(n_1197),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1332),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1295),
.B(n_1173),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1413),
.A2(n_1369),
.B1(n_1276),
.B2(n_1426),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1343),
.B(n_1197),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1325),
.A2(n_284),
.B1(n_301),
.B2(n_1197),
.Y(n_1488)
);

AOI221xp5_ASAP7_75t_L g1489 ( 
.A1(n_1431),
.A2(n_355),
.B1(n_1224),
.B2(n_1171),
.C(n_43),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1295),
.B(n_1213),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1413),
.A2(n_1172),
.B(n_1224),
.C(n_355),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1345),
.B(n_1213),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1345),
.B(n_1389),
.Y(n_1493)
);

BUFx12f_ASAP7_75t_L g1494 ( 
.A(n_1281),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1332),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1303),
.B(n_38),
.Y(n_1496)
);

NOR3xp33_ASAP7_75t_SL g1497 ( 
.A(n_1375),
.B(n_40),
.C(n_41),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1303),
.B(n_1329),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1419),
.Y(n_1499)
);

AO22x2_ASAP7_75t_L g1500 ( 
.A1(n_1399),
.A2(n_1430),
.B1(n_1405),
.B2(n_1364),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1329),
.B(n_40),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1345),
.B(n_1213),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1286),
.A2(n_355),
.B1(n_44),
.B2(n_46),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1355),
.B(n_355),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1299),
.A2(n_355),
.B1(n_304),
.B2(n_1213),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1267),
.Y(n_1506)
);

OAI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1286),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1299),
.A2(n_1283),
.B1(n_1317),
.B2(n_1328),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1267),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1389),
.B(n_1195),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1288),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1371),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1337),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1314),
.A2(n_304),
.B1(n_48),
.B2(n_50),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1330),
.A2(n_304),
.B1(n_53),
.B2(n_54),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1288),
.Y(n_1516)
);

AND2x4_ASAP7_75t_SL g1517 ( 
.A(n_1390),
.B(n_102),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1314),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_1518)
);

OAI221xp5_ASAP7_75t_L g1519 ( 
.A1(n_1275),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.C(n_69),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1298),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1381),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.C(n_77),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1297),
.B(n_74),
.Y(n_1522)
);

BUFx10_ASAP7_75t_L g1523 ( 
.A(n_1365),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1330),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1304),
.B(n_84),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1297),
.B(n_84),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1383),
.A2(n_85),
.B(n_86),
.C(n_90),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1429),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1335),
.B(n_1333),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1398),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1414),
.A2(n_1336),
.B(n_1342),
.C(n_1266),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1296),
.A2(n_1360),
.B1(n_1425),
.B2(n_1400),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1391),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1416),
.B(n_92),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1404),
.B(n_93),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1390),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1389),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1270),
.A2(n_93),
.B1(n_101),
.B2(n_109),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1356),
.A2(n_122),
.B(n_123),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1349),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1300),
.A2(n_187),
.B1(n_133),
.B2(n_134),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1391),
.A2(n_128),
.B1(n_135),
.B2(n_137),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1398),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1333),
.A2(n_139),
.B(n_140),
.C(n_143),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1344),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1344),
.A2(n_147),
.B1(n_154),
.B2(n_159),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1300),
.A2(n_185),
.B1(n_168),
.B2(n_170),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1300),
.A2(n_163),
.B1(n_174),
.B2(n_175),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1359),
.A2(n_176),
.B1(n_1363),
.B2(n_1362),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1271),
.A2(n_1430),
.B(n_1399),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1318),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1323),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1404),
.Y(n_1553)
);

NOR2x1_ASAP7_75t_SL g1554 ( 
.A(n_1300),
.B(n_1326),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1359),
.Y(n_1555)
);

OAI221xp5_ASAP7_75t_L g1556 ( 
.A1(n_1313),
.A2(n_1382),
.B1(n_1351),
.B2(n_1363),
.C(n_1362),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1356),
.A2(n_1287),
.B(n_1320),
.Y(n_1557)
);

CKINVDCx11_ASAP7_75t_R g1558 ( 
.A(n_1402),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1415),
.A2(n_1350),
.B1(n_1427),
.B2(n_1353),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1415),
.A2(n_1350),
.B1(n_1427),
.B2(n_1404),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1389),
.A2(n_1380),
.B1(n_1349),
.B2(n_1421),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1389),
.A2(n_1349),
.B1(n_1380),
.B2(n_1388),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1402),
.Y(n_1564)
);

BUFx2_ASAP7_75t_L g1565 ( 
.A(n_1402),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1380),
.B(n_1420),
.Y(n_1566)
);

BUFx3_ASAP7_75t_L g1567 ( 
.A(n_1380),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_SL g1568 ( 
.A(n_1412),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1420),
.A2(n_1412),
.B1(n_1350),
.B2(n_1417),
.Y(n_1569)
);

NOR3xp33_ASAP7_75t_SL g1570 ( 
.A(n_1422),
.B(n_1394),
.C(n_1316),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1420),
.B(n_1280),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1280),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1289),
.B(n_1306),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1412),
.Y(n_1574)
);

NAND2xp33_ASAP7_75t_SL g1575 ( 
.A(n_1326),
.B(n_1408),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1291),
.A2(n_1312),
.B(n_1372),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1374),
.A2(n_1377),
.B1(n_1396),
.B2(n_1385),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1298),
.Y(n_1578)
);

AOI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1417),
.A2(n_1401),
.B1(n_1408),
.B2(n_1398),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1308),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1366),
.A2(n_1388),
.B1(n_1361),
.B2(n_1268),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1289),
.B(n_1315),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1374),
.A2(n_1377),
.B1(n_1378),
.B2(n_1372),
.C(n_1428),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1393),
.A2(n_1261),
.B(n_1387),
.Y(n_1584)
);

BUFx4f_ASAP7_75t_SL g1585 ( 
.A(n_1428),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_L g1586 ( 
.A1(n_1374),
.A2(n_1377),
.B1(n_1378),
.B2(n_1385),
.C(n_1396),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1366),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1393),
.A2(n_1261),
.B(n_1387),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1293),
.B(n_1309),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1293),
.B(n_1315),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1294),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1366),
.A2(n_1388),
.B1(n_1268),
.B2(n_1361),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1294),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1268),
.A2(n_1361),
.B1(n_1378),
.B2(n_1374),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1306),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1309),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1302),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1378),
.A2(n_1377),
.B1(n_1321),
.B2(n_1368),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1321),
.A2(n_1368),
.B1(n_1271),
.B2(n_1396),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1385),
.A2(n_1396),
.B1(n_1364),
.B2(n_1386),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1302),
.B(n_1273),
.Y(n_1601)
);

NAND2x1p5_ASAP7_75t_L g1602 ( 
.A(n_1321),
.B(n_1341),
.Y(n_1602)
);

OAI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1436),
.A2(n_1385),
.B1(n_1392),
.B2(n_1386),
.C(n_1348),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1524),
.A2(n_1321),
.B1(n_1376),
.B2(n_1347),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1498),
.B(n_1334),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1524),
.A2(n_1376),
.B1(n_1347),
.B2(n_1392),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1484),
.B(n_1334),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1486),
.B(n_1409),
.Y(n_1608)
);

OR2x6_ASAP7_75t_L g1609 ( 
.A(n_1459),
.B(n_1423),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1436),
.A2(n_1274),
.B1(n_1423),
.B2(n_1265),
.Y(n_1610)
);

AOI221xp5_ASAP7_75t_L g1611 ( 
.A1(n_1503),
.A2(n_1274),
.B1(n_1334),
.B2(n_1308),
.C(n_1273),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1444),
.A2(n_1274),
.B1(n_1265),
.B2(n_1311),
.Y(n_1612)
);

AND2x4_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1409),
.Y(n_1613)
);

OAI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1515),
.A2(n_1507),
.B1(n_1519),
.B2(n_1503),
.Y(n_1614)
);

AOI222xp33_ASAP7_75t_L g1615 ( 
.A1(n_1507),
.A2(n_1277),
.B1(n_1279),
.B2(n_1305),
.C1(n_1290),
.C2(n_1334),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1495),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1456),
.A2(n_1469),
.B1(n_1508),
.B2(n_1477),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1545),
.B(n_1334),
.Y(n_1618)
);

AOI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1497),
.A2(n_1458),
.B1(n_1521),
.B2(n_1531),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1523),
.A2(n_1265),
.B1(n_1311),
.B2(n_1358),
.Y(n_1620)
);

NAND2x1_ASAP7_75t_L g1621 ( 
.A(n_1536),
.B(n_1311),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1435),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1518),
.A2(n_1497),
.B1(n_1514),
.B2(n_1531),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1555),
.B(n_1308),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1518),
.A2(n_1287),
.B1(n_1311),
.B2(n_1265),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1474),
.B(n_1308),
.Y(n_1626)
);

AOI221xp5_ASAP7_75t_L g1627 ( 
.A1(n_1514),
.A2(n_1533),
.B1(n_1527),
.B2(n_1440),
.C(n_1586),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1552),
.A2(n_1341),
.B1(n_1339),
.B2(n_1424),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1445),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1585),
.Y(n_1630)
);

NAND3xp33_ASAP7_75t_L g1631 ( 
.A(n_1527),
.B(n_1308),
.C(n_1273),
.Y(n_1631)
);

AO221x1_ASAP7_75t_L g1632 ( 
.A1(n_1471),
.A2(n_1367),
.B1(n_1358),
.B2(n_1406),
.C(n_1424),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1508),
.A2(n_1277),
.B1(n_1279),
.B2(n_1290),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1477),
.A2(n_1305),
.B1(n_1310),
.B2(n_1339),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1504),
.A2(n_1310),
.B1(n_1346),
.B2(n_1357),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1538),
.A2(n_1273),
.B1(n_1367),
.B2(n_1346),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1535),
.A2(n_1354),
.B1(n_1357),
.B2(n_1384),
.Y(n_1637)
);

AOI222xp33_ASAP7_75t_L g1638 ( 
.A1(n_1489),
.A2(n_1273),
.B1(n_1354),
.B2(n_1384),
.C1(n_1379),
.C2(n_1406),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1541),
.A2(n_1379),
.B1(n_1548),
.B2(n_1547),
.Y(n_1639)
);

OAI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1451),
.A2(n_1482),
.B1(n_1454),
.B2(n_1522),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1510),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1466),
.Y(n_1642)
);

OAI22xp5_ASAP7_75t_L g1643 ( 
.A1(n_1541),
.A2(n_1547),
.B1(n_1548),
.B2(n_1463),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1453),
.A2(n_1463),
.B1(n_1513),
.B2(n_1457),
.Y(n_1644)
);

CKINVDCx14_ASAP7_75t_R g1645 ( 
.A(n_1441),
.Y(n_1645)
);

AND2x4_ASAP7_75t_L g1646 ( 
.A(n_1492),
.B(n_1502),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1504),
.A2(n_1525),
.B1(n_1439),
.B2(n_1443),
.Y(n_1647)
);

INVx5_ASAP7_75t_L g1648 ( 
.A(n_1459),
.Y(n_1648)
);

NOR2x1_ASAP7_75t_L g1649 ( 
.A(n_1528),
.B(n_1453),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1485),
.A2(n_1442),
.B1(n_1476),
.B2(n_1523),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1501),
.B(n_1478),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1476),
.A2(n_1433),
.B1(n_1446),
.B2(n_1502),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1492),
.A2(n_1597),
.B1(n_1532),
.B2(n_1434),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1437),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1560),
.A2(n_1562),
.B1(n_1475),
.B2(n_1479),
.Y(n_1655)
);

AOI211xp5_ASAP7_75t_L g1656 ( 
.A1(n_1535),
.A2(n_1526),
.B(n_1544),
.C(n_1549),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1455),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1490),
.B(n_1580),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1576),
.A2(n_1438),
.B(n_1470),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1529),
.B(n_1571),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1560),
.A2(n_1562),
.B1(n_1559),
.B2(n_1496),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_SL g1662 ( 
.A1(n_1517),
.A2(n_1472),
.B(n_1544),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1596),
.B(n_1551),
.Y(n_1663)
);

INVx4_ASAP7_75t_L g1664 ( 
.A(n_1585),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1559),
.A2(n_1556),
.B1(n_1595),
.B2(n_1582),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1512),
.Y(n_1666)
);

BUFx8_ASAP7_75t_SL g1667 ( 
.A(n_1494),
.Y(n_1667)
);

AO31x2_ASAP7_75t_L g1668 ( 
.A1(n_1598),
.A2(n_1599),
.A3(n_1594),
.B(n_1491),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1582),
.B(n_1590),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1590),
.A2(n_1568),
.B1(n_1432),
.B2(n_1505),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1572),
.B(n_1591),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1568),
.A2(n_1505),
.B1(n_1464),
.B2(n_1558),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1528),
.A2(n_1499),
.B1(n_1448),
.B2(n_1542),
.Y(n_1673)
);

OAI22xp33_ASAP7_75t_L g1674 ( 
.A1(n_1448),
.A2(n_1499),
.B1(n_1546),
.B2(n_1540),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1540),
.A2(n_1567),
.B1(n_1459),
.B2(n_1449),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1554),
.B(n_1449),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1534),
.B(n_1566),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1577),
.A2(n_1583),
.B1(n_1491),
.B2(n_1600),
.C(n_1465),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1593),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1488),
.A2(n_1536),
.B1(n_1449),
.B2(n_1450),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1577),
.A2(n_1516),
.B1(n_1565),
.B2(n_1564),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1589),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1450),
.A2(n_1579),
.B1(n_1600),
.B2(n_1488),
.C(n_1570),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1566),
.B(n_1561),
.Y(n_1684)
);

AO22x1_ASAP7_75t_L g1685 ( 
.A1(n_1493),
.A2(n_1487),
.B1(n_1481),
.B2(n_1452),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1567),
.A2(n_1449),
.B1(n_1462),
.B2(n_1460),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1493),
.A2(n_1509),
.B1(n_1520),
.B2(n_1511),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1462),
.A2(n_1517),
.B1(n_1553),
.B2(n_1483),
.Y(n_1688)
);

AOI222xp33_ASAP7_75t_L g1689 ( 
.A1(n_1573),
.A2(n_1601),
.B1(n_1563),
.B2(n_1530),
.C1(n_1543),
.C2(n_1480),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1575),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1452),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1481),
.B(n_1487),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1530),
.A2(n_1543),
.B1(n_1500),
.B2(n_1550),
.C(n_1563),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1574),
.Y(n_1694)
);

OAI211xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1570),
.A2(n_1584),
.B(n_1588),
.C(n_1468),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1447),
.B(n_1574),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1602),
.A2(n_1510),
.B1(n_1587),
.B2(n_1467),
.C(n_1462),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1500),
.B(n_1587),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1473),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1460),
.A2(n_1592),
.B1(n_1581),
.B2(n_1447),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1500),
.B(n_1511),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1460),
.A2(n_1473),
.B(n_1557),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1537),
.A2(n_1473),
.B1(n_1539),
.B2(n_1506),
.Y(n_1703)
);

CKINVDCx11_ASAP7_75t_R g1704 ( 
.A(n_1537),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1537),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1578),
.Y(n_1706)
);

AOI221xp5_ASAP7_75t_L g1707 ( 
.A1(n_1461),
.A2(n_737),
.B1(n_497),
.B2(n_612),
.C(n_500),
.Y(n_1707)
);

NAND3xp33_ASAP7_75t_L g1708 ( 
.A(n_1461),
.B(n_737),
.C(n_591),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1461),
.B(n_1498),
.Y(n_1709)
);

BUFx8_ASAP7_75t_SL g1710 ( 
.A(n_1461),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_1512),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1436),
.A2(n_737),
.B1(n_497),
.B2(n_612),
.C(n_500),
.Y(n_1712)
);

OAI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1497),
.A2(n_737),
.B(n_591),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1484),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1498),
.B(n_1484),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1498),
.B(n_1484),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1498),
.B(n_1484),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1436),
.A2(n_737),
.B1(n_497),
.B2(n_612),
.C(n_500),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1524),
.A2(n_737),
.B1(n_999),
.B2(n_1436),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1524),
.A2(n_737),
.B1(n_999),
.B2(n_1436),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_L g1721 ( 
.A1(n_1436),
.A2(n_1259),
.B1(n_1070),
.B2(n_1228),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1510),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1585),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1484),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1527),
.A2(n_737),
.B(n_593),
.C(n_1264),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1498),
.B(n_1529),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1498),
.B(n_1484),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1484),
.Y(n_1728)
);

OAI222xp33_ASAP7_75t_L g1729 ( 
.A1(n_1436),
.A2(n_1264),
.B1(n_1260),
.B2(n_516),
.C1(n_1141),
.C2(n_1292),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1527),
.A2(n_737),
.B(n_593),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1436),
.A2(n_1259),
.B1(n_1070),
.B2(n_1228),
.Y(n_1731)
);

OAI22xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1436),
.A2(n_999),
.B1(n_1264),
.B2(n_881),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1524),
.A2(n_737),
.B1(n_999),
.B2(n_1436),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1569),
.B(n_1492),
.Y(n_1734)
);

OAI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1436),
.A2(n_591),
.B1(n_737),
.B2(n_598),
.C(n_1264),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1436),
.A2(n_1259),
.B1(n_1070),
.B2(n_1228),
.Y(n_1736)
);

INVx6_ASAP7_75t_L g1737 ( 
.A(n_1574),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1436),
.A2(n_1259),
.B1(n_1070),
.B2(n_1228),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1524),
.A2(n_1518),
.B(n_1515),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1512),
.Y(n_1740)
);

AOI222xp33_ASAP7_75t_L g1741 ( 
.A1(n_1436),
.A2(n_1292),
.B1(n_1259),
.B2(n_737),
.C1(n_1141),
.C2(n_1264),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_SL g1742 ( 
.A1(n_1436),
.A2(n_1259),
.B1(n_1264),
.B2(n_1228),
.Y(n_1742)
);

OAI221xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1436),
.A2(n_737),
.B1(n_591),
.B2(n_598),
.C(n_1141),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1436),
.A2(n_1259),
.B1(n_1070),
.B2(n_1228),
.Y(n_1744)
);

AOI222xp33_ASAP7_75t_L g1745 ( 
.A1(n_1436),
.A2(n_1292),
.B1(n_1259),
.B2(n_737),
.C1(n_1141),
.C2(n_1264),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1699),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1699),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1616),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1690),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1714),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1709),
.B(n_1605),
.Y(n_1751)
);

BUFx3_ASAP7_75t_L g1752 ( 
.A(n_1613),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1658),
.B(n_1709),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1605),
.B(n_1715),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1624),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1724),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1699),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1622),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1728),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1715),
.B(n_1716),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1679),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1658),
.B(n_1626),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1660),
.B(n_1726),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1671),
.B(n_1607),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1729),
.A2(n_1712),
.B1(n_1718),
.B2(n_1743),
.C(n_1719),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1671),
.B(n_1618),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1629),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1716),
.B(n_1717),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1717),
.B(n_1727),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1682),
.B(n_1727),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1613),
.B(n_1668),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1642),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1613),
.B(n_1668),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1668),
.B(n_1609),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1668),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1610),
.B(n_1708),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1654),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1625),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1609),
.B(n_1608),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1641),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1608),
.B(n_1669),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1669),
.B(n_1689),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1657),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1659),
.B(n_1611),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1632),
.B(n_1637),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1646),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1734),
.B(n_1702),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1725),
.A2(n_1623),
.B(n_1643),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1663),
.B(n_1620),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1631),
.B(n_1734),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1650),
.B(n_1665),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1701),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1621),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1619),
.B(n_1628),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1745),
.A2(n_1741),
.B1(n_1720),
.B2(n_1733),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1722),
.B(n_1638),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1703),
.Y(n_1797)
);

AO21x2_ASAP7_75t_L g1798 ( 
.A1(n_1636),
.A2(n_1604),
.B(n_1639),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1706),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1646),
.B(n_1698),
.Y(n_1800)
);

NOR2xp33_ASAP7_75t_L g1801 ( 
.A(n_1730),
.B(n_1713),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1646),
.B(n_1698),
.Y(n_1802)
);

NOR2x1_ASAP7_75t_R g1803 ( 
.A(n_1664),
.B(n_1723),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1651),
.B(n_1615),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1606),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1640),
.B(n_1678),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1603),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1695),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1710),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1633),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1635),
.B(n_1677),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1762),
.B(n_1681),
.Y(n_1812)
);

OAI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1801),
.A2(n_1735),
.B(n_1739),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1749),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1754),
.B(n_1684),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1746),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1754),
.B(n_1644),
.Y(n_1817)
);

BUFx6f_ASAP7_75t_L g1818 ( 
.A(n_1786),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1801),
.B(n_1707),
.C(n_1627),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1749),
.Y(n_1820)
);

OAI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1788),
.A2(n_1656),
.B(n_1662),
.C(n_1742),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1763),
.B(n_1645),
.Y(n_1822)
);

NAND4xp25_ASAP7_75t_L g1823 ( 
.A(n_1795),
.B(n_1744),
.C(n_1721),
.D(n_1731),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1795),
.A2(n_1765),
.B1(n_1806),
.B2(n_1794),
.C(n_1784),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1772),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1754),
.B(n_1653),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1760),
.B(n_1649),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1749),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_SL g1829 ( 
.A(n_1765),
.B(n_1738),
.C(n_1736),
.Y(n_1829)
);

OAI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1806),
.A2(n_1614),
.B1(n_1683),
.B2(n_1647),
.Y(n_1830)
);

NAND3xp33_ASAP7_75t_L g1831 ( 
.A(n_1784),
.B(n_1672),
.C(n_1670),
.Y(n_1831)
);

OAI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1794),
.A2(n_1732),
.B1(n_1661),
.B2(n_1652),
.C(n_1655),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1752),
.B(n_1648),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1758),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1772),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1808),
.A2(n_1673),
.B1(n_1723),
.B2(n_1664),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1799),
.Y(n_1837)
);

OAI322xp33_ASAP7_75t_L g1838 ( 
.A1(n_1776),
.A2(n_1645),
.A3(n_1674),
.B1(n_1630),
.B2(n_1664),
.C1(n_1723),
.C2(n_1688),
.Y(n_1838)
);

OAI33xp33_ASAP7_75t_L g1839 ( 
.A1(n_1807),
.A2(n_1680),
.A3(n_1700),
.B1(n_1675),
.B2(n_1692),
.B3(n_1686),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1808),
.A2(n_1630),
.B1(n_1617),
.B2(n_1737),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1767),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1758),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1799),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1791),
.A2(n_1691),
.B1(n_1612),
.B2(n_1685),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1808),
.B(n_1693),
.C(n_1634),
.Y(n_1845)
);

AOI33xp33_ASAP7_75t_L g1846 ( 
.A1(n_1785),
.A2(n_1687),
.A3(n_1676),
.B1(n_1667),
.B2(n_1711),
.B3(n_1740),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1791),
.A2(n_1710),
.B1(n_1648),
.B2(n_1697),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1758),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1760),
.B(n_1694),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1758),
.Y(n_1850)
);

NOR3xp33_ASAP7_75t_L g1851 ( 
.A(n_1785),
.B(n_1696),
.C(n_1705),
.Y(n_1851)
);

AOI21xp5_ASAP7_75t_L g1852 ( 
.A1(n_1798),
.A2(n_1676),
.B(n_1705),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1807),
.A2(n_1691),
.B1(n_1704),
.B2(n_1737),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1760),
.B(n_1737),
.Y(n_1854)
);

OAI221xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1771),
.A2(n_1667),
.B1(n_1704),
.B2(n_1711),
.C(n_1666),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1767),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1798),
.A2(n_1666),
.B(n_1740),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1768),
.B(n_1769),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1768),
.B(n_1769),
.Y(n_1859)
);

BUFx3_ASAP7_75t_L g1860 ( 
.A(n_1780),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1768),
.B(n_1769),
.Y(n_1861)
);

NAND2xp33_ASAP7_75t_R g1862 ( 
.A(n_1809),
.B(n_1771),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1751),
.B(n_1771),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1751),
.B(n_1773),
.Y(n_1864)
);

HB1xp67_ASAP7_75t_L g1865 ( 
.A(n_1755),
.Y(n_1865)
);

OR2x6_ASAP7_75t_L g1866 ( 
.A(n_1752),
.B(n_1773),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1767),
.Y(n_1867)
);

OAI211xp5_ASAP7_75t_SL g1868 ( 
.A1(n_1778),
.A2(n_1776),
.B(n_1805),
.C(n_1781),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_SL g1869 ( 
.A1(n_1773),
.A2(n_1809),
.B1(n_1804),
.B2(n_1774),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1748),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1798),
.A2(n_1810),
.B1(n_1804),
.B2(n_1782),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1751),
.B(n_1811),
.Y(n_1872)
);

OAI31xp33_ASAP7_75t_L g1873 ( 
.A1(n_1805),
.A2(n_1804),
.A3(n_1778),
.B(n_1775),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1837),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1863),
.B(n_1864),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1816),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1865),
.Y(n_1877)
);

INVx1_ASAP7_75t_SL g1878 ( 
.A(n_1814),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1866),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1825),
.B(n_1785),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1841),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1841),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1863),
.B(n_1798),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1864),
.B(n_1798),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1856),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1866),
.B(n_1752),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1856),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1819),
.B(n_1775),
.C(n_1797),
.Y(n_1888)
);

INVx1_ASAP7_75t_SL g1889 ( 
.A(n_1814),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1872),
.B(n_1774),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1825),
.B(n_1764),
.Y(n_1891)
);

AOI21xp33_ASAP7_75t_L g1892 ( 
.A1(n_1819),
.A2(n_1797),
.B(n_1789),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1872),
.B(n_1753),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1858),
.B(n_1779),
.Y(n_1894)
);

AND2x4_ASAP7_75t_L g1895 ( 
.A(n_1866),
.B(n_1752),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1858),
.B(n_1774),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1816),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1835),
.B(n_1764),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1867),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1866),
.B(n_1786),
.Y(n_1900)
);

BUFx3_ASAP7_75t_L g1901 ( 
.A(n_1820),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1859),
.B(n_1796),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1867),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1835),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1870),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1816),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1870),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1873),
.B(n_1766),
.Y(n_1908)
);

AND2x2_ASAP7_75t_SL g1909 ( 
.A(n_1871),
.B(n_1790),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1843),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1834),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1861),
.B(n_1753),
.Y(n_1912)
);

NOR2xp33_ASAP7_75t_L g1913 ( 
.A(n_1822),
.B(n_1763),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1859),
.B(n_1779),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1834),
.Y(n_1915)
);

INVxp33_ASAP7_75t_L g1916 ( 
.A(n_1869),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1842),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1842),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1812),
.B(n_1828),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1848),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1866),
.B(n_1779),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1873),
.B(n_1766),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1848),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1850),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1850),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1815),
.B(n_1796),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1905),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1919),
.B(n_1828),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1905),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1902),
.B(n_1875),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1880),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1907),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1876),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1907),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1876),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1881),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1881),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1919),
.B(n_1812),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1882),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1901),
.B(n_1857),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1882),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1885),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1908),
.B(n_1922),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1908),
.B(n_1820),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1879),
.Y(n_1945)
);

BUFx2_ASAP7_75t_L g1946 ( 
.A(n_1879),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1909),
.A2(n_1845),
.B1(n_1829),
.B2(n_1824),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1922),
.B(n_1817),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1902),
.B(n_1869),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1885),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1887),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1913),
.B(n_1855),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1926),
.B(n_1815),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_SL g1954 ( 
.A(n_1878),
.B(n_1838),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1886),
.B(n_1852),
.Y(n_1955)
);

NAND2x2_ASAP7_75t_L g1956 ( 
.A(n_1901),
.B(n_1860),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1902),
.B(n_1849),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1876),
.Y(n_1958)
);

INVx4_ASAP7_75t_L g1959 ( 
.A(n_1901),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_L g1960 ( 
.A(n_1878),
.B(n_1868),
.Y(n_1960)
);

NAND2x1p5_ASAP7_75t_L g1961 ( 
.A(n_1886),
.B(n_1786),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1887),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1899),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1875),
.B(n_1849),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_L g1965 ( 
.A(n_1889),
.B(n_1838),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1926),
.B(n_1845),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1880),
.B(n_1770),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1926),
.B(n_1770),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1944),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1948),
.B(n_1883),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1968),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1927),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1947),
.A2(n_1909),
.B1(n_1916),
.B2(n_1892),
.Y(n_1973)
);

NAND4xp75_ASAP7_75t_L g1974 ( 
.A(n_1965),
.B(n_1813),
.C(n_1909),
.D(n_1892),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1930),
.B(n_1883),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1948),
.B(n_1883),
.Y(n_1976)
);

INVx4_ASAP7_75t_L g1977 ( 
.A(n_1959),
.Y(n_1977)
);

NOR4xp25_ASAP7_75t_SL g1978 ( 
.A(n_1946),
.B(n_1862),
.C(n_1832),
.D(n_1809),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1943),
.B(n_1884),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1929),
.Y(n_1980)
);

OAI22xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1960),
.A2(n_1888),
.B1(n_1889),
.B2(n_1836),
.Y(n_1981)
);

INVxp67_ASAP7_75t_SL g1982 ( 
.A(n_1940),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1952),
.B(n_1943),
.Y(n_1983)
);

NOR3xp33_ASAP7_75t_L g1984 ( 
.A(n_1959),
.B(n_1821),
.C(n_1830),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1930),
.B(n_1949),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1949),
.B(n_1884),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1954),
.A2(n_1888),
.B(n_1884),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_SL g1988 ( 
.A(n_1955),
.B(n_1886),
.Y(n_1988)
);

NAND5xp2_ASAP7_75t_SL g1989 ( 
.A(n_1956),
.B(n_1851),
.C(n_1853),
.D(n_1875),
.E(n_1896),
.Y(n_1989)
);

OR2x2_ASAP7_75t_L g1990 ( 
.A(n_1938),
.B(n_1912),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1966),
.B(n_1874),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1938),
.B(n_1874),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1957),
.B(n_1896),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1944),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1968),
.B(n_1912),
.Y(n_1995)
);

NOR3xp33_ASAP7_75t_SL g1996 ( 
.A(n_1953),
.B(n_1839),
.C(n_1910),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1932),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1934),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1967),
.B(n_1891),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1957),
.B(n_1896),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1939),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1931),
.B(n_1910),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1967),
.B(n_1891),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1964),
.B(n_1877),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1939),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1964),
.B(n_1894),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1946),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1928),
.B(n_1898),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1961),
.B(n_1894),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_1928),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1941),
.Y(n_2011)
);

NOR3xp33_ASAP7_75t_L g2012 ( 
.A(n_1959),
.B(n_1831),
.C(n_1846),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_SL g2013 ( 
.A(n_1955),
.B(n_1886),
.Y(n_2013)
);

AOI22xp33_ASAP7_75t_L g2014 ( 
.A1(n_1973),
.A2(n_1831),
.B1(n_1823),
.B2(n_1810),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1977),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1983),
.B(n_1945),
.Y(n_2016)
);

OAI32xp33_ASAP7_75t_L g2017 ( 
.A1(n_1984),
.A2(n_1956),
.A3(n_1945),
.B1(n_1961),
.B2(n_1823),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_2001),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1974),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2001),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1981),
.A2(n_1961),
.B1(n_1895),
.B2(n_1900),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2005),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1974),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2005),
.Y(n_2024)
);

OAI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1981),
.A2(n_1895),
.B1(n_1900),
.B2(n_1955),
.Y(n_2025)
);

INVxp67_ASAP7_75t_L g2026 ( 
.A(n_1969),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2011),
.Y(n_2027)
);

XNOR2xp5_ASAP7_75t_L g2028 ( 
.A(n_2012),
.B(n_1840),
.Y(n_2028)
);

OAI221xp5_ASAP7_75t_L g2029 ( 
.A1(n_1987),
.A2(n_1844),
.B1(n_1789),
.B2(n_1782),
.C(n_1933),
.Y(n_2029)
);

AOI22xp33_ASAP7_75t_L g2030 ( 
.A1(n_1989),
.A2(n_1810),
.B1(n_1844),
.B2(n_1796),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1990),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1996),
.B(n_1936),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1982),
.B(n_1895),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2011),
.Y(n_2034)
);

OAI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1978),
.A2(n_1895),
.B1(n_1900),
.B2(n_1893),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1989),
.A2(n_1790),
.B1(n_1847),
.B2(n_1787),
.Y(n_2036)
);

INVx1_ASAP7_75t_SL g2037 ( 
.A(n_1994),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2007),
.B(n_1937),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2010),
.Y(n_2039)
);

AOI21xp33_ASAP7_75t_L g2040 ( 
.A1(n_1991),
.A2(n_1935),
.B(n_1933),
.Y(n_2040)
);

AOI22xp5_ASAP7_75t_L g2041 ( 
.A1(n_1986),
.A2(n_1979),
.B1(n_1976),
.B2(n_1971),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1985),
.B(n_1977),
.Y(n_2042)
);

OAI221xp5_ASAP7_75t_L g2043 ( 
.A1(n_1970),
.A2(n_1935),
.B1(n_1958),
.B2(n_1826),
.C(n_1790),
.Y(n_2043)
);

NAND2xp33_ASAP7_75t_SL g2044 ( 
.A(n_1978),
.B(n_1914),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1985),
.B(n_1914),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1972),
.Y(n_2046)
);

A2O1A1Ixp33_ASAP7_75t_L g2047 ( 
.A1(n_1970),
.A2(n_1921),
.B(n_1890),
.C(n_1787),
.Y(n_2047)
);

INVxp67_ASAP7_75t_SL g2048 ( 
.A(n_1992),
.Y(n_2048)
);

AOI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1986),
.A2(n_1971),
.B1(n_1990),
.B2(n_1811),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1993),
.B(n_1890),
.Y(n_2050)
);

AND2x2_ASAP7_75t_SL g2051 ( 
.A(n_2019),
.B(n_2023),
.Y(n_2051)
);

AOI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_2019),
.A2(n_2013),
.B1(n_1988),
.B2(n_2007),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2030),
.A2(n_1995),
.B1(n_2009),
.B2(n_2000),
.Y(n_2053)
);

OAI211xp5_ASAP7_75t_L g2054 ( 
.A1(n_2023),
.A2(n_1977),
.B(n_2002),
.C(n_2009),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2042),
.B(n_2006),
.Y(n_2055)
);

NOR2xp33_ASAP7_75t_L g2056 ( 
.A(n_2037),
.B(n_1977),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2020),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2020),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_2044),
.B(n_2008),
.Y(n_2059)
);

OAI32xp33_ASAP7_75t_L g2060 ( 
.A1(n_2044),
.A2(n_2032),
.A3(n_2025),
.B1(n_2021),
.B2(n_2029),
.Y(n_2060)
);

O2A1O1Ixp33_ASAP7_75t_L g2061 ( 
.A1(n_2017),
.A2(n_1997),
.B(n_1998),
.C(n_1980),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_2028),
.A2(n_1995),
.B1(n_1993),
.B2(n_2000),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_R g2063 ( 
.A(n_2015),
.B(n_1972),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2022),
.Y(n_2064)
);

AOI221xp5_ASAP7_75t_L g2065 ( 
.A1(n_2017),
.A2(n_2014),
.B1(n_2040),
.B2(n_2048),
.C(n_2043),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2022),
.Y(n_2066)
);

NAND2x1_ASAP7_75t_L g2067 ( 
.A(n_2042),
.B(n_2006),
.Y(n_2067)
);

OAI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_2049),
.A2(n_2008),
.B1(n_2003),
.B2(n_1999),
.Y(n_2068)
);

OAI21xp33_ASAP7_75t_L g2069 ( 
.A1(n_2028),
.A2(n_1980),
.B(n_1998),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2031),
.B(n_1975),
.Y(n_2070)
);

AOI211xp5_ASAP7_75t_SL g2071 ( 
.A1(n_2026),
.A2(n_1975),
.B(n_1997),
.C(n_2004),
.Y(n_2071)
);

OAI222xp33_ASAP7_75t_L g2072 ( 
.A1(n_2036),
.A2(n_2003),
.B1(n_1999),
.B2(n_1958),
.C1(n_1890),
.C2(n_1792),
.Y(n_2072)
);

AOI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_2016),
.A2(n_1811),
.B1(n_1787),
.B2(n_1942),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2042),
.A2(n_2039),
.B(n_2033),
.Y(n_2074)
);

INVx1_ASAP7_75t_SL g2075 ( 
.A(n_2031),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2045),
.B(n_1950),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2041),
.A2(n_1900),
.B1(n_1921),
.B2(n_1893),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2070),
.B(n_2038),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2057),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2058),
.Y(n_2080)
);

NOR2x1_ASAP7_75t_SL g2081 ( 
.A(n_2054),
.B(n_2015),
.Y(n_2081)
);

NOR4xp25_ASAP7_75t_SL g2082 ( 
.A(n_2059),
.B(n_2034),
.C(n_2024),
.D(n_2046),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_2075),
.B(n_2045),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_2069),
.B(n_2046),
.Y(n_2084)
);

INVxp67_ASAP7_75t_SL g2085 ( 
.A(n_2061),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2064),
.Y(n_2086)
);

INVx4_ASAP7_75t_L g2087 ( 
.A(n_2051),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2051),
.B(n_2050),
.Y(n_2088)
);

NOR3xp33_ASAP7_75t_L g2089 ( 
.A(n_2065),
.B(n_2024),
.C(n_2034),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2071),
.B(n_2050),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2066),
.Y(n_2091)
);

OAI21xp5_ASAP7_75t_SL g2092 ( 
.A1(n_2052),
.A2(n_2035),
.B(n_2047),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2076),
.Y(n_2093)
);

A2O1A1Ixp33_ASAP7_75t_L g2094 ( 
.A1(n_2060),
.A2(n_2027),
.B(n_2018),
.C(n_1941),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2055),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2056),
.Y(n_2096)
);

OAI211xp5_ASAP7_75t_SL g2097 ( 
.A1(n_2074),
.A2(n_1963),
.B(n_1942),
.C(n_1962),
.Y(n_2097)
);

NAND3xp33_ASAP7_75t_L g2098 ( 
.A(n_2094),
.B(n_2056),
.C(n_2062),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2083),
.Y(n_2099)
);

NAND4xp25_ASAP7_75t_L g2100 ( 
.A(n_2084),
.B(n_2053),
.C(n_2077),
.D(n_2073),
.Y(n_2100)
);

NOR4xp25_ASAP7_75t_L g2101 ( 
.A(n_2085),
.B(n_2072),
.C(n_2068),
.D(n_2063),
.Y(n_2101)
);

INVx2_ASAP7_75t_SL g2102 ( 
.A(n_2095),
.Y(n_2102)
);

NOR3xp33_ASAP7_75t_L g2103 ( 
.A(n_2087),
.B(n_2068),
.C(n_2067),
.Y(n_2103)
);

OAI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_2085),
.A2(n_2063),
.B(n_2073),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2087),
.Y(n_2105)
);

O2A1O1Ixp33_ASAP7_75t_L g2106 ( 
.A1(n_2089),
.A2(n_1963),
.B(n_1951),
.C(n_1877),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2088),
.Y(n_2107)
);

NOR3xp33_ASAP7_75t_L g2108 ( 
.A(n_2089),
.B(n_1906),
.C(n_1897),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2079),
.Y(n_2109)
);

NOR4xp25_ASAP7_75t_L g2110 ( 
.A(n_2096),
.B(n_1904),
.C(n_1903),
.D(n_1899),
.Y(n_2110)
);

OAI211xp5_ASAP7_75t_L g2111 ( 
.A1(n_2101),
.A2(n_2082),
.B(n_2092),
.C(n_2084),
.Y(n_2111)
);

AOI31xp33_ASAP7_75t_L g2112 ( 
.A1(n_2098),
.A2(n_2090),
.A3(n_2078),
.B(n_2093),
.Y(n_2112)
);

AOI321xp33_ASAP7_75t_L g2113 ( 
.A1(n_2104),
.A2(n_2091),
.A3(n_2080),
.B1(n_2086),
.B2(n_2081),
.C(n_2097),
.Y(n_2113)
);

AOI22xp33_ASAP7_75t_SL g2114 ( 
.A1(n_2107),
.A2(n_1818),
.B1(n_1781),
.B2(n_1827),
.Y(n_2114)
);

A2O1A1Ixp33_ASAP7_75t_L g2115 ( 
.A1(n_2106),
.A2(n_1897),
.B(n_1906),
.C(n_1904),
.Y(n_2115)
);

OAI211xp5_ASAP7_75t_SL g2116 ( 
.A1(n_2103),
.A2(n_1898),
.B(n_1903),
.C(n_1793),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2106),
.A2(n_2108),
.B(n_2100),
.Y(n_2117)
);

AOI221xp5_ASAP7_75t_L g2118 ( 
.A1(n_2110),
.A2(n_1897),
.B1(n_1906),
.B2(n_1748),
.C(n_1750),
.Y(n_2118)
);

AOI221xp5_ASAP7_75t_L g2119 ( 
.A1(n_2099),
.A2(n_1761),
.B1(n_1759),
.B2(n_1750),
.C(n_1756),
.Y(n_2119)
);

NAND4xp25_ASAP7_75t_L g2120 ( 
.A(n_2105),
.B(n_1860),
.C(n_1793),
.D(n_1854),
.Y(n_2120)
);

NOR4xp25_ASAP7_75t_L g2121 ( 
.A(n_2109),
.B(n_1761),
.C(n_1759),
.D(n_1756),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2112),
.B(n_2102),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2117),
.Y(n_2123)
);

AOI21x1_ASAP7_75t_L g2124 ( 
.A1(n_2111),
.A2(n_1854),
.B(n_1915),
.Y(n_2124)
);

NOR3xp33_ASAP7_75t_L g2125 ( 
.A(n_2116),
.B(n_1803),
.C(n_1917),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2121),
.B(n_1770),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_2120),
.Y(n_2127)
);

OAI211xp5_ASAP7_75t_SL g2128 ( 
.A1(n_2123),
.A2(n_2113),
.B(n_2114),
.C(n_2115),
.Y(n_2128)
);

XNOR2x1_ASAP7_75t_L g2129 ( 
.A(n_2122),
.B(n_1833),
.Y(n_2129)
);

AOI321xp33_ASAP7_75t_L g2130 ( 
.A1(n_2124),
.A2(n_2118),
.A3(n_2119),
.B1(n_1783),
.B2(n_1777),
.C(n_1911),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2127),
.B(n_1860),
.Y(n_2131)
);

XNOR2x1_ASAP7_75t_L g2132 ( 
.A(n_2126),
.B(n_1833),
.Y(n_2132)
);

NAND4xp75_ASAP7_75t_L g2133 ( 
.A(n_2125),
.B(n_1800),
.C(n_1802),
.D(n_1911),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2126),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2134),
.A2(n_1793),
.B1(n_1746),
.B2(n_1757),
.Y(n_2135)
);

BUFx8_ASAP7_75t_L g2136 ( 
.A(n_2131),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2130),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_2132),
.B(n_1924),
.Y(n_2138)
);

NAND4xp25_ASAP7_75t_L g2139 ( 
.A(n_2128),
.B(n_1803),
.C(n_1793),
.D(n_1747),
.Y(n_2139)
);

XNOR2xp5_ASAP7_75t_L g2140 ( 
.A(n_2129),
.B(n_1833),
.Y(n_2140)
);

AND2x4_ASAP7_75t_L g2141 ( 
.A(n_2137),
.B(n_2138),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2136),
.Y(n_2142)
);

CKINVDCx20_ASAP7_75t_R g2143 ( 
.A(n_2140),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2135),
.B(n_2139),
.Y(n_2144)
);

INVx4_ASAP7_75t_L g2145 ( 
.A(n_2142),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2145),
.A2(n_2141),
.B1(n_2143),
.B2(n_2144),
.Y(n_2146)
);

AND3x1_ASAP7_75t_L g2147 ( 
.A(n_2146),
.B(n_2130),
.C(n_2133),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2146),
.Y(n_2148)
);

NAND3xp33_ASAP7_75t_L g2149 ( 
.A(n_2148),
.B(n_2147),
.C(n_1924),
.Y(n_2149)
);

OAI22xp5_ASAP7_75t_L g2150 ( 
.A1(n_2147),
.A2(n_1793),
.B1(n_1924),
.B2(n_1746),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_2150),
.A2(n_1746),
.B1(n_1757),
.B2(n_1925),
.Y(n_2151)
);

AOI32xp33_ASAP7_75t_L g2152 ( 
.A1(n_2149),
.A2(n_1833),
.A3(n_1923),
.B1(n_1920),
.B2(n_1918),
.Y(n_2152)
);

AOI322xp5_ASAP7_75t_L g2153 ( 
.A1(n_2152),
.A2(n_1925),
.A3(n_1917),
.B1(n_1915),
.B2(n_1923),
.C1(n_1918),
.C2(n_1920),
.Y(n_2153)
);

AOI221xp5_ASAP7_75t_L g2154 ( 
.A1(n_2153),
.A2(n_2151),
.B1(n_1783),
.B2(n_1777),
.C(n_1818),
.Y(n_2154)
);

AOI211xp5_ASAP7_75t_L g2155 ( 
.A1(n_2154),
.A2(n_1818),
.B(n_1763),
.C(n_1757),
.Y(n_2155)
);


endmodule