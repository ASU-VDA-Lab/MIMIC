module fake_jpeg_12214_n_578 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_578);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_578;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_18),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_54),
.B(n_74),
.Y(n_127)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_60),
.Y(n_136)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_62),
.B(n_64),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_23),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_70),
.Y(n_160)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g120 ( 
.A(n_72),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_73),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_16),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_78),
.Y(n_151)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_90),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_45),
.B(n_14),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_89),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_14),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_33),
.B(n_14),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_38),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_96),
.Y(n_133)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_33),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_102),
.Y(n_179)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_20),
.Y(n_103)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_105),
.B(n_53),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_34),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_34),
.B(n_27),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_34),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_46),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_108),
.Y(n_171)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_112),
.B(n_126),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_123),
.B(n_169),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_59),
.Y(n_126)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx11_ASAP7_75t_L g195 ( 
.A(n_128),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_93),
.B(n_27),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_130),
.B(n_157),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_137),
.Y(n_180)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_143),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_71),
.B(n_26),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_155),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_110),
.B(n_26),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_63),
.B(n_31),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_70),
.A2(n_51),
.B1(n_53),
.B2(n_46),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_49),
.B1(n_52),
.B2(n_40),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_102),
.B(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_166),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_83),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_52),
.C(n_49),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_55),
.B(n_24),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_63),
.B(n_31),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_87),
.B(n_21),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_173),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_73),
.Y(n_173)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_88),
.Y(n_196)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_182),
.Y(n_251)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_183),
.Y(n_247)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_184),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_185),
.A2(n_225),
.B1(n_231),
.B2(n_122),
.Y(n_273)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_186),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_111),
.B1(n_97),
.B2(n_91),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_188),
.A2(n_205),
.B1(n_206),
.B2(n_228),
.Y(n_266)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_190),
.Y(n_250)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_191),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_194),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_214),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_124),
.B(n_41),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_198),
.B(n_201),
.Y(n_268)
);

CKINVDCx12_ASAP7_75t_R g199 ( 
.A(n_120),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_199),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_200),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_127),
.B(n_41),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_151),
.A2(n_87),
.B1(n_88),
.B2(n_39),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_203),
.A2(n_216),
.B1(n_220),
.B2(n_223),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_133),
.B(n_39),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_208),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_109),
.B1(n_77),
.B2(n_75),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_117),
.A2(n_57),
.B1(n_82),
.B2(n_86),
.Y(n_206)
);

BUFx24_ASAP7_75t_L g207 ( 
.A(n_136),
.Y(n_207)
);

BUFx8_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_118),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_148),
.B(n_44),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_210),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_44),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_131),
.B(n_100),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_221),
.Y(n_270)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_60),
.B1(n_52),
.B2(n_49),
.Y(n_213)
);

AO21x2_ASAP7_75t_SL g288 ( 
.A1(n_213),
.A2(n_143),
.B(n_140),
.Y(n_288)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_151),
.A2(n_58),
.B1(n_92),
.B2(n_43),
.Y(n_216)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_101),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_232),
.C(n_161),
.Y(n_279)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_134),
.Y(n_219)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_132),
.A2(n_43),
.B1(n_93),
.B2(n_21),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_178),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_222),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_132),
.A2(n_43),
.B1(n_48),
.B2(n_47),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_125),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_171),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_138),
.A2(n_48),
.B1(n_47),
.B2(n_42),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_227),
.A2(n_237),
.B1(n_239),
.B2(n_3),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_L g228 ( 
.A1(n_115),
.A2(n_49),
.B1(n_108),
.B2(n_51),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_113),
.A2(n_51),
.B1(n_42),
.B2(n_73),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_150),
.B(n_114),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_119),
.B(n_13),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_233),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_138),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_142),
.B(n_0),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_178),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_234),
.B(n_238),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_147),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_236),
.B(n_244),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

AOI21xp33_ASAP7_75t_L g238 ( 
.A1(n_141),
.A2(n_3),
.B(n_4),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_170),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_145),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_139),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_152),
.B(n_156),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g252 ( 
.A1(n_206),
.A2(n_176),
.B1(n_115),
.B2(n_135),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_252),
.A2(n_288),
.B1(n_189),
.B2(n_215),
.Y(n_323)
);

AOI32xp33_ASAP7_75t_L g253 ( 
.A1(n_192),
.A2(n_187),
.A3(n_202),
.B1(n_180),
.B2(n_236),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_253),
.A2(n_255),
.B(n_263),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_214),
.A2(n_160),
.B1(n_176),
.B2(n_179),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_254),
.A2(n_267),
.B1(n_289),
.B2(n_290),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_179),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_257),
.B(n_261),
.C(n_286),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_122),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_213),
.B(n_135),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_264),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_196),
.A2(n_171),
.B(n_114),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_185),
.A2(n_160),
.B1(n_113),
.B2(n_161),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_207),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_269),
.B(n_247),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_273),
.B(n_279),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_278),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_196),
.B(n_149),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_232),
.B(n_149),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_292),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_205),
.A2(n_164),
.B1(n_140),
.B2(n_139),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_229),
.A2(n_164),
.B1(n_139),
.B2(n_178),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_207),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_291),
.B(n_217),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_209),
.B(n_210),
.Y(n_292)
);

BUFx4f_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_262),
.A2(n_290),
.B1(n_279),
.B2(n_254),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_283),
.Y(n_296)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_297),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_246),
.B(n_235),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_300),
.B(n_301),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_256),
.B(n_226),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_303),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_246),
.B(n_197),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_253),
.B(n_183),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_306),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_292),
.B(n_213),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_268),
.B(n_213),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_309),
.B(n_310),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_281),
.Y(n_310)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_195),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_312),
.B(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_313),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_259),
.B(n_181),
.C(n_224),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_327),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_270),
.B(n_222),
.Y(n_315)
);

INVx4_ASAP7_75t_SL g316 ( 
.A(n_271),
.Y(n_316)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_316),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_228),
.B1(n_218),
.B2(n_212),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_317),
.A2(n_288),
.B1(n_255),
.B2(n_284),
.Y(n_359)
);

INVx13_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_272),
.B(n_182),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_321),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_323),
.A2(n_333),
.B1(n_335),
.B2(n_245),
.Y(n_349)
);

INVx13_ASAP7_75t_L g324 ( 
.A(n_271),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_282),
.Y(n_326)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_326),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_259),
.B(n_218),
.C(n_186),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_316),
.Y(n_373)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_329),
.Y(n_363)
);

BUFx8_ASAP7_75t_L g330 ( 
.A(n_269),
.Y(n_330)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_330),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_194),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_331),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_284),
.B(n_240),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_332),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_250),
.Y(n_333)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_184),
.C(n_195),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_334),
.B(n_257),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_266),
.A2(n_190),
.B1(n_237),
.B2(n_239),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_336),
.A2(n_267),
.B1(n_262),
.B2(n_245),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_285),
.B(n_241),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_264),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_340),
.A2(n_341),
.B1(n_349),
.B2(n_350),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_322),
.A2(n_266),
.B1(n_261),
.B2(n_288),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_322),
.A2(n_336),
.B1(n_323),
.B2(n_306),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_352),
.B(n_334),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_307),
.A2(n_275),
.B(n_263),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_353),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_322),
.A2(n_288),
.B1(n_287),
.B2(n_286),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_355),
.A2(n_369),
.B1(n_375),
.B2(n_295),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_325),
.A2(n_277),
.B1(n_249),
.B2(n_258),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_330),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g391 ( 
.A(n_358),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_311),
.B1(n_299),
.B2(n_308),
.Y(n_392)
);

OAI32xp33_ASAP7_75t_L g360 ( 
.A1(n_318),
.A2(n_258),
.A3(n_294),
.B1(n_241),
.B2(n_282),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_370),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g404 ( 
.A(n_361),
.B(n_299),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_309),
.A2(n_286),
.B1(n_264),
.B2(n_280),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_318),
.B(n_294),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_251),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_310),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_373),
.B(n_330),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_311),
.A2(n_250),
.B1(n_251),
.B2(n_265),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_303),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_378),
.B(n_393),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_298),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_382),
.C(n_383),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_380),
.Y(n_432)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_298),
.C(n_327),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_307),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_375),
.Y(n_438)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_347),
.Y(n_386)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_386),
.Y(n_430)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_344),
.A2(n_311),
.B1(n_314),
.B2(n_312),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_389),
.A2(n_342),
.B(n_368),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_395),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_392),
.A2(n_405),
.B1(n_369),
.B2(n_340),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_370),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_343),
.B(n_348),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_394),
.B(n_400),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_330),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_354),
.B(n_297),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_397),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_367),
.Y(n_397)
);

NOR2x1_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_300),
.Y(n_398)
);

NOR3xp33_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_373),
.C(n_362),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_355),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_338),
.B(n_329),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_347),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_346),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_402),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_341),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_344),
.A2(n_305),
.B1(n_296),
.B2(n_308),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_406),
.B(n_407),
.Y(n_416)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_366),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_274),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_410),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_365),
.A2(n_319),
.B(n_320),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_409),
.A2(n_411),
.B(n_351),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_363),
.B(n_274),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_419),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_390),
.B(n_354),
.Y(n_417)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_417),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_418),
.A2(n_424),
.B(n_438),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_353),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_420),
.B(n_426),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_382),
.B(n_383),
.C(n_399),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_429),
.C(n_415),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_350),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_398),
.B(n_358),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_428),
.B(n_433),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_372),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_396),
.B(n_362),
.Y(n_431)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_431),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_391),
.B(n_409),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_391),
.B(n_304),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_434),
.B(n_391),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_442),
.B1(n_381),
.B2(n_376),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_377),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_385),
.B(n_367),
.Y(n_441)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_392),
.A2(n_374),
.B1(n_366),
.B2(n_319),
.Y(n_442)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_411),
.B1(n_385),
.B2(n_404),
.Y(n_446)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_446),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_464),
.C(n_423),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_418),
.A2(n_395),
.B1(n_377),
.B2(n_403),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_451),
.A2(n_458),
.B1(n_468),
.B2(n_448),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_461),
.Y(n_474)
);

OAI21xp33_ASAP7_75t_L g454 ( 
.A1(n_436),
.A2(n_373),
.B(n_384),
.Y(n_454)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_454),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_455),
.A2(n_456),
.B1(n_462),
.B2(n_465),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_397),
.B1(n_386),
.B2(n_401),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_431),
.B(n_391),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_458),
.Y(n_476)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_417),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_414),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_460),
.Y(n_481)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_416),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_438),
.A2(n_397),
.B1(n_374),
.B2(n_319),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_326),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_463),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_356),
.C(n_351),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_442),
.A2(n_356),
.B1(n_333),
.B2(n_335),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_427),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_467),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_421),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_413),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_470),
.A2(n_473),
.B1(n_425),
.B2(n_422),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_313),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_471),
.Y(n_498)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_422),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_472),
.B(n_419),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_475),
.B(n_482),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_477),
.B(n_483),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_480),
.A2(n_496),
.B1(n_465),
.B2(n_456),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_420),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_449),
.B(n_426),
.C(n_412),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_429),
.C(n_424),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_490),
.C(n_495),
.Y(n_499)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g487 ( 
.A(n_451),
.B(n_413),
.Y(n_487)
);

O2A1O1Ixp33_ASAP7_75t_L g512 ( 
.A1(n_487),
.A2(n_233),
.B(n_240),
.C(n_243),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_447),
.B(n_441),
.C(n_430),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_453),
.A2(n_430),
.B(n_425),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g502 ( 
.A1(n_491),
.A2(n_457),
.B(n_459),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_469),
.A2(n_439),
.B(n_435),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_492),
.A2(n_494),
.B(n_3),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_452),
.A2(n_439),
.B(n_435),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_443),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_452),
.A2(n_333),
.B1(n_335),
.B2(n_200),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_450),
.B(n_455),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_497),
.B(n_462),
.Y(n_507)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_500),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_476),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_501),
.B(n_517),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_502),
.A2(n_503),
.B(n_512),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_489),
.A2(n_450),
.B(n_460),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_488),
.Y(n_504)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_504),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_485),
.A2(n_448),
.B1(n_473),
.B2(n_461),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_505),
.A2(n_509),
.B1(n_496),
.B2(n_480),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_507),
.B(n_497),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_493),
.A2(n_193),
.B1(n_324),
.B2(n_316),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_479),
.B(n_227),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_510),
.B(n_498),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_491),
.Y(n_530)
);

INVx13_ASAP7_75t_L g514 ( 
.A(n_494),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_516),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_487),
.A2(n_233),
.B(n_243),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_515),
.A2(n_479),
.B(n_495),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_478),
.Y(n_516)
);

FAx1_ASAP7_75t_SL g517 ( 
.A(n_490),
.B(n_3),
.CI(n_4),
.CON(n_517),
.SN(n_517)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_520),
.B(n_523),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_474),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_504),
.B(n_477),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_524),
.B(n_525),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_516),
.B(n_492),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_499),
.B(n_484),
.C(n_475),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_533),
.C(n_519),
.Y(n_538)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_527),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_513),
.A2(n_483),
.B(n_481),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_530),
.B(n_517),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_506),
.B(n_482),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_532),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_499),
.B(n_485),
.C(n_487),
.Y(n_533)
);

CKINVDCx16_ASAP7_75t_R g535 ( 
.A(n_534),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_535),
.B(n_539),
.Y(n_554)
);

AO21x1_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_508),
.B(n_503),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_536),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_518),
.A2(n_505),
.B1(n_508),
.B2(n_502),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_537),
.A2(n_548),
.B1(n_527),
.B2(n_500),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_547),
.C(n_506),
.Y(n_553)
);

BUFx24_ASAP7_75t_SL g539 ( 
.A(n_522),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_544),
.B(n_541),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g547 ( 
.A1(n_526),
.A2(n_514),
.B(n_509),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g548 ( 
.A1(n_521),
.A2(n_515),
.B1(n_514),
.B2(n_512),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_550),
.B(n_556),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_533),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_552),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_529),
.C(n_531),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_557),
.C(n_7),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_555),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_529),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_545),
.A2(n_517),
.B1(n_510),
.B2(n_530),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_532),
.C(n_511),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_558),
.A2(n_559),
.B(n_549),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_546),
.B(n_6),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_560),
.B(n_563),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_549),
.A2(n_540),
.B(n_536),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g570 ( 
.A1(n_562),
.A2(n_566),
.B(n_561),
.Y(n_570)
);

AOI322xp5_ASAP7_75t_L g563 ( 
.A1(n_554),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_558),
.C(n_552),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_567),
.B(n_569),
.Y(n_572)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_565),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_7),
.Y(n_571)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_571),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_572),
.A2(n_568),
.B(n_569),
.Y(n_574)
);

A2O1A1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_7),
.B(n_10),
.C(n_11),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_575),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_573),
.C(n_11),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_10),
.B1(n_12),
.B2(n_351),
.Y(n_578)
);


endmodule