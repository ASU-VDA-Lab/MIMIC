module fake_jpeg_3012_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_19),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_55),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_35),
.Y(n_52)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_48),
.B(n_14),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_48),
.C(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_0),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_39),
.B1(n_47),
.B2(n_45),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_63),
.B1(n_52),
.B2(n_36),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_49),
.B1(n_43),
.B2(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_1),
.Y(n_80)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_47),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_62),
.B(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_66),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_45),
.A3(n_41),
.B1(n_38),
.B2(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_44),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_57),
.B1(n_51),
.B2(n_41),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_77),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_51),
.B1(n_38),
.B2(n_3),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_78),
.A2(n_79),
.B1(n_64),
.B2(n_61),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_53),
.B1(n_17),
.B2(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_77),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_90),
.B(n_92),
.Y(n_96)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_91),
.B1(n_10),
.B2(n_11),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_8),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_25),
.C(n_26),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_93),
.A2(n_71),
.B1(n_27),
.B2(n_13),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_93),
.A2(n_30),
.B1(n_33),
.B2(n_24),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_10),
.C(n_11),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_31),
.C(n_32),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_107),
.C(n_89),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_34),
.C(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_113),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_81),
.B1(n_91),
.B2(n_101),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_107),
.C(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_95),
.A3(n_96),
.B1(n_106),
.B2(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_115),
.B(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_118),
.C(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_112),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_111),
.Y(n_124)
);


endmodule