module fake_jpeg_25819_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_13),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_31),
.Y(n_55)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_26),
.B1(n_19),
.B2(n_25),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_41),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_84)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_31),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_55),
.Y(n_71)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_26),
.B1(n_25),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_40),
.B1(n_39),
.B2(n_36),
.Y(n_76)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_55),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_72),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_40),
.B1(n_32),
.B2(n_26),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_76),
.B1(n_50),
.B2(n_42),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_28),
.B1(n_25),
.B2(n_23),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_62),
.Y(n_93)
);

OR2x2_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_28),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_16),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_20),
.B1(n_29),
.B2(n_36),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_74),
.B1(n_42),
.B2(n_30),
.Y(n_108)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_77),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_51),
.A2(n_29),
.B1(n_36),
.B2(n_40),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_47),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_80),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_37),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_23),
.B(n_35),
.C(n_15),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_49),
.B(n_35),
.Y(n_95)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_43),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_44),
.B(n_21),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_56),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_100),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_76),
.Y(n_123)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_95),
.A2(n_101),
.B(n_78),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_75),
.B1(n_84),
.B2(n_59),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_66),
.B1(n_61),
.B2(n_53),
.Y(n_139)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_0),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_110),
.Y(n_121)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_42),
.B1(n_51),
.B2(n_56),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_105),
.A2(n_81),
.B1(n_67),
.B2(n_73),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_109),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_108),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_69),
.B(n_43),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_80),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_15),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_70),
.B1(n_77),
.B2(n_62),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_117),
.B1(n_123),
.B2(n_133),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_126),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_122),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_132),
.B(n_96),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_71),
.B(n_65),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_137),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_63),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_114),
.C(n_93),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_71),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_79),
.B(n_85),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_91),
.B1(n_103),
.B2(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_87),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g138 ( 
.A(n_98),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_139),
.A2(n_141),
.B1(n_104),
.B2(n_88),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_97),
.B(n_31),
.C(n_24),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_140),
.B(n_96),
.C(n_104),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_24),
.B1(n_27),
.B2(n_18),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_96),
.A2(n_113),
.B(n_109),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_27),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_27),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_146),
.B(n_156),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_148),
.B(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_150),
.Y(n_178)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_155),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_89),
.B(n_92),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_157),
.B(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_92),
.B(n_90),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_99),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_99),
.B(n_94),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_111),
.B(n_88),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_130),
.B1(n_134),
.B2(n_17),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_87),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_24),
.C(n_18),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_119),
.C(n_140),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_18),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_167),
.A2(n_119),
.B1(n_120),
.B2(n_130),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_192),
.C(n_204),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_173),
.B(n_155),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_123),
.B1(n_120),
.B2(n_137),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_203),
.B1(n_163),
.B2(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_174),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_193),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_137),
.C(n_126),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_198),
.C(n_172),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_150),
.A2(n_123),
.B(n_141),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_205),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_151),
.B(n_15),
.C(n_16),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_146),
.C(n_154),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_134),
.C(n_130),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_209),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_157),
.C(n_148),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_213),
.C(n_214),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_210),
.A2(n_212),
.B1(n_196),
.B2(n_194),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_176),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_218),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_206),
.A2(n_169),
.B(n_165),
.C(n_175),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_164),
.C(n_158),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_185),
.B(n_147),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_221),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_144),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_165),
.C(n_173),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_229),
.C(n_230),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_182),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_197),
.B(n_156),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_226),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_225),
.Y(n_234)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_188),
.B(n_198),
.Y(n_227)
);

NAND4xp25_ASAP7_75t_SL g228 ( 
.A(n_200),
.B(n_17),
.C(n_149),
.D(n_145),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_145),
.C(n_13),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_12),
.C(n_11),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_193),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_240),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_186),
.C(n_177),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_249),
.C(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_213),
.B(n_202),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_177),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_247),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_188),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_212),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_187),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_248),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_186),
.C(n_195),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_224),
.A2(n_181),
.B1(n_196),
.B2(n_179),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_179),
.B1(n_199),
.B2(n_220),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_181),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_257),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_232),
.B(n_184),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_258),
.A2(n_250),
.B1(n_234),
.B2(n_249),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_212),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_212),
.B(n_228),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_264),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_203),
.Y(n_264)
);

AOI221xp5_ASAP7_75t_L g265 ( 
.A1(n_237),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.C(n_4),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_10),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_238),
.C(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_269),
.C(n_277),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_231),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_1),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_233),
.C(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_262),
.B(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_266),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_273),
.A2(n_261),
.B1(n_254),
.B2(n_251),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_253),
.A2(n_236),
.B1(n_239),
.B2(n_244),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_9),
.C(n_2),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_286),
.Y(n_298)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_274),
.B(n_252),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_288),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_251),
.Y(n_287)
);

AOI221xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_290),
.B1(n_270),
.B2(n_268),
.C(n_285),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_269),
.C(n_278),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_260),
.B1(n_2),
.B2(n_3),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_290),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_260),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_4),
.B(n_5),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_291),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_272),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_6),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_281),
.A2(n_270),
.B(n_277),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_299),
.A2(n_7),
.B(n_8),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_300),
.A2(n_6),
.B(n_7),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_287),
.B(n_7),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_300),
.B(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_295),
.B(n_294),
.Y(n_309)
);

OAI31xp33_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.A3(n_301),
.B(n_302),
.Y(n_310)
);

OAI31xp33_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_298),
.A3(n_307),
.B(n_9),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_9),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_312),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_8),
.Y(n_314)
);


endmodule