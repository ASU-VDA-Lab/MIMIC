module fake_jpeg_14754_n_175 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_175);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_12),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_5),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_34),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_17),
.B(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_37),
.B(n_41),
.Y(n_80)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_10),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_20),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_13),
.B(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_51),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_0),
.C(n_1),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_9),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_24),
.A2(n_28),
.B1(n_20),
.B2(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_52),
.B(n_56),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_15),
.B(n_6),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_25),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_74),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_71),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_25),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_33),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_81),
.Y(n_104)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_30),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_35),
.B(n_21),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_52),
.B(n_21),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_90),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_23),
.B1(n_18),
.B2(n_8),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_84),
.B1(n_51),
.B2(n_47),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_57),
.A2(n_23),
.B1(n_18),
.B2(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_0),
.Y(n_87)
);

CKINVDCx6p67_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_21),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_65),
.A2(n_90),
.B1(n_82),
.B2(n_89),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_59),
.B1(n_63),
.B2(n_60),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_65),
.A2(n_50),
.B1(n_49),
.B2(n_42),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_108),
.B1(n_116),
.B2(n_86),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_41),
.B(n_36),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_64),
.B(n_80),
.Y(n_117)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_102),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_106),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_76),
.A2(n_48),
.B1(n_55),
.B2(n_38),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_54),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_115),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_112),
.A2(n_64),
.B1(n_63),
.B2(n_60),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_114),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_45),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_21),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_76),
.A2(n_38),
.B1(n_45),
.B2(n_49),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_127),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_75),
.B1(n_81),
.B2(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_123),
.B1(n_125),
.B2(n_128),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_109),
.B1(n_104),
.B2(n_116),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_72),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_94),
.A2(n_71),
.B1(n_42),
.B2(n_40),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_69),
.B(n_72),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_126),
.B(n_132),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_113),
.A2(n_92),
.B1(n_93),
.B2(n_108),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_59),
.C(n_67),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_100),
.C(n_99),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_101),
.Y(n_132)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_86),
.C(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_133),
.B(n_111),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_138),
.A2(n_140),
.B1(n_150),
.B2(n_131),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_104),
.B1(n_109),
.B2(n_105),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_148),
.A3(n_136),
.B1(n_130),
.B2(n_118),
.Y(n_158)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_144),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_96),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_149),
.C(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_102),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_106),
.B1(n_91),
.B2(n_107),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_146),
.B1(n_138),
.B2(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_158),
.B1(n_147),
.B2(n_146),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_145),
.A2(n_133),
.B1(n_124),
.B2(n_125),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_152),
.A2(n_140),
.B(n_137),
.C(n_123),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_119),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_162),
.C(n_164),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_149),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_165),
.B(n_152),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_136),
.C(n_132),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_153),
.C(n_155),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_168),
.C(n_167),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_170),
.C(n_103),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_161),
.C(n_103),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_67),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_171),
.C(n_103),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);


endmodule