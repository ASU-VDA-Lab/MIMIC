module real_aes_1423_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_838, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_837, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_838;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_837;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_693;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g169 ( .A(n_0), .B(n_143), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_1), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_2), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g134 ( .A(n_3), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_4), .B(n_127), .Y(n_196) );
NAND2xp33_ASAP7_75t_SL g239 ( .A(n_5), .B(n_133), .Y(n_239) );
INVx1_ASAP7_75t_L g231 ( .A(n_6), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_7), .B(n_201), .Y(n_490) );
INVx1_ASAP7_75t_L g471 ( .A(n_8), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g830 ( .A(n_9), .Y(n_830) );
AND2x2_ASAP7_75t_L g194 ( .A(n_10), .B(n_151), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_11), .Y(n_554) );
INVx2_ASAP7_75t_L g149 ( .A(n_12), .Y(n_149) );
CKINVDCx16_ASAP7_75t_R g435 ( .A(n_13), .Y(n_435) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_13), .B(n_829), .C(n_831), .Y(n_828) );
INVx1_ASAP7_75t_L g498 ( .A(n_14), .Y(n_498) );
AOI221x1_ASAP7_75t_L g234 ( .A1(n_15), .A2(n_136), .B1(n_235), .B2(n_237), .C(n_238), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_16), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g780 ( .A(n_17), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_18), .Y(n_792) );
INVx1_ASAP7_75t_L g496 ( .A(n_19), .Y(n_496) );
INVx1_ASAP7_75t_SL g508 ( .A(n_20), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_21), .B(n_128), .Y(n_486) );
AOI221xp5_ASAP7_75t_SL g158 ( .A1(n_22), .A2(n_44), .B1(n_127), .B2(n_136), .C(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_23), .A2(n_136), .B(n_198), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_24), .B(n_143), .Y(n_199) );
AOI33xp33_ASAP7_75t_L g463 ( .A1(n_25), .A2(n_56), .A3(n_182), .B1(n_189), .B2(n_464), .B3(n_465), .Y(n_463) );
INVxp33_ASAP7_75t_L g834 ( .A(n_26), .Y(n_834) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_27), .A2(n_42), .B1(n_817), .B2(n_818), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_27), .Y(n_818) );
INVx1_ASAP7_75t_L g548 ( .A(n_28), .Y(n_548) );
OAI22xp5_ASAP7_75t_SL g108 ( .A1(n_29), .A2(n_109), .B1(n_110), .B2(n_116), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_29), .Y(n_116) );
OA21x2_ASAP7_75t_L g148 ( .A1(n_30), .A2(n_93), .B(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g152 ( .A(n_30), .B(n_93), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_31), .B(n_145), .Y(n_144) );
INVxp67_ASAP7_75t_L g233 ( .A(n_32), .Y(n_233) );
AND2x2_ASAP7_75t_L g220 ( .A(n_33), .B(n_157), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_34), .B(n_180), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_35), .A2(n_136), .B(n_168), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_36), .B(n_651), .Y(n_650) );
CKINVDCx16_ASAP7_75t_R g774 ( .A(n_36), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_37), .B(n_145), .Y(n_160) );
AND2x2_ASAP7_75t_L g133 ( .A(n_38), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g137 ( .A(n_38), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g188 ( .A(n_38), .Y(n_188) );
OR2x6_ASAP7_75t_L g778 ( .A(n_39), .B(n_779), .Y(n_778) );
INVxp67_ASAP7_75t_L g831 ( .A(n_39), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_40), .A2(n_73), .B1(n_813), .B2(n_814), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_40), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_41), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_42), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_43), .B(n_180), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_45), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_45), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_46), .A2(n_165), .B1(n_201), .B2(n_480), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_47), .A2(n_85), .B1(n_136), .B2(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_48), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_49), .B(n_128), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_50), .B(n_143), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_51), .B(n_147), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_52), .B(n_128), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_53), .Y(n_483) );
AND2x2_ASAP7_75t_L g172 ( .A(n_54), .B(n_157), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_55), .B(n_157), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_57), .B(n_128), .Y(n_454) );
INVx1_ASAP7_75t_L g130 ( .A(n_58), .Y(n_130) );
INVx1_ASAP7_75t_L g140 ( .A(n_58), .Y(n_140) );
AND2x2_ASAP7_75t_L g455 ( .A(n_59), .B(n_157), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_60), .A2(n_78), .B1(n_180), .B2(n_186), .C(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_61), .B(n_180), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_62), .B(n_127), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_63), .B(n_165), .Y(n_556) );
AOI21xp5_ASAP7_75t_SL g516 ( .A1(n_64), .A2(n_186), .B(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g211 ( .A(n_65), .B(n_157), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_66), .B(n_145), .Y(n_170) );
AND2x2_ASAP7_75t_SL g150 ( .A(n_67), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_68), .B(n_143), .Y(n_208) );
INVx1_ASAP7_75t_L g493 ( .A(n_69), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_70), .A2(n_136), .B(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g452 ( .A(n_71), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_72), .B(n_145), .Y(n_200) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_73), .B(n_147), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_73), .Y(n_813) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_74), .A2(n_186), .B(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_SL g113 ( .A1(n_75), .A2(n_97), .B1(n_114), .B2(n_115), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_75), .Y(n_114) );
INVx1_ASAP7_75t_L g132 ( .A(n_76), .Y(n_132) );
INVx1_ASAP7_75t_L g138 ( .A(n_76), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_77), .B(n_180), .Y(n_466) );
AND2x2_ASAP7_75t_L g510 ( .A(n_79), .B(n_237), .Y(n_510) );
INVx1_ASAP7_75t_L g494 ( .A(n_80), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_81), .A2(n_186), .B(n_507), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_82), .A2(n_177), .B(n_186), .C(n_485), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_83), .A2(n_88), .B1(n_127), .B2(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_84), .B(n_127), .Y(n_209) );
INVx1_ASAP7_75t_L g781 ( .A(n_86), .Y(n_781) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_87), .B(n_237), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_89), .A2(n_186), .B1(n_461), .B2(n_462), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_90), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_91), .B(n_143), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_92), .A2(n_136), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g518 ( .A(n_94), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_95), .B(n_145), .Y(n_207) );
AND2x2_ASAP7_75t_L g467 ( .A(n_96), .B(n_237), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_97), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_98), .A2(n_546), .B(n_547), .C(n_549), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_99), .B(n_127), .Y(n_171) );
INVxp67_ASAP7_75t_L g236 ( .A(n_100), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_101), .B(n_145), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_102), .A2(n_136), .B(n_141), .Y(n_135) );
BUFx2_ASAP7_75t_L g803 ( .A(n_103), .Y(n_803) );
BUFx2_ASAP7_75t_SL g823 ( .A(n_103), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_104), .B(n_128), .Y(n_519) );
AOI21xp33_ASAP7_75t_SL g105 ( .A1(n_106), .A2(n_824), .B(n_833), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_804), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_117), .B(n_776), .C(n_782), .Y(n_107) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_108), .A2(n_777), .B(n_778), .Y(n_776) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_108), .Y(n_789) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_433), .B(n_436), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx3_ASAP7_75t_SL g788 ( .A(n_119), .Y(n_788) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_325), .Y(n_119) );
NOR3xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_253), .C(n_303), .Y(n_120) );
OAI211xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_173), .B(n_221), .C(n_242), .Y(n_121) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_153), .Y(n_122) );
AND2x2_ASAP7_75t_L g252 ( .A(n_123), .B(n_154), .Y(n_252) );
INVx1_ASAP7_75t_L g383 ( .A(n_123), .Y(n_383) );
NOR2x1p5_ASAP7_75t_L g415 ( .A(n_123), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g226 ( .A(n_124), .B(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g274 ( .A(n_124), .Y(n_274) );
OR2x2_ASAP7_75t_L g278 ( .A(n_124), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_124), .B(n_156), .Y(n_290) );
OR2x2_ASAP7_75t_L g312 ( .A(n_124), .B(n_156), .Y(n_312) );
AND2x4_ASAP7_75t_L g318 ( .A(n_124), .B(n_282), .Y(n_318) );
OR2x2_ASAP7_75t_L g335 ( .A(n_124), .B(n_228), .Y(n_335) );
INVx1_ASAP7_75t_L g370 ( .A(n_124), .Y(n_370) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_124), .Y(n_392) );
OR2x2_ASAP7_75t_L g406 ( .A(n_124), .B(n_339), .Y(n_406) );
AND2x4_ASAP7_75t_SL g410 ( .A(n_124), .B(n_228), .Y(n_410) );
OR2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_150), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_135), .B(n_147), .Y(n_125) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_133), .Y(n_127) );
INVx1_ASAP7_75t_L g240 ( .A(n_128), .Y(n_240) );
AND2x4_ASAP7_75t_L g128 ( .A(n_129), .B(n_131), .Y(n_128) );
AND2x6_ASAP7_75t_L g143 ( .A(n_129), .B(n_138), .Y(n_143) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g145 ( .A(n_131), .B(n_140), .Y(n_145) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx5_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_133), .Y(n_549) );
AND2x2_ASAP7_75t_L g139 ( .A(n_134), .B(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_134), .Y(n_183) );
AND2x6_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
BUFx3_ASAP7_75t_L g184 ( .A(n_137), .Y(n_184) );
INVx2_ASAP7_75t_L g190 ( .A(n_138), .Y(n_190) );
AND2x4_ASAP7_75t_L g186 ( .A(n_139), .B(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_144), .B(n_146), .Y(n_141) );
INVxp67_ASAP7_75t_L g497 ( .A(n_143), .Y(n_497) );
INVxp67_ASAP7_75t_L g499 ( .A(n_145), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_146), .A2(n_160), .B(n_161), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_146), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_146), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_146), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_146), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_146), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g461 ( .A(n_146), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g470 ( .A1(n_146), .A2(n_453), .B(n_471), .C(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_146), .A2(n_486), .B(n_487), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_146), .B(n_201), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_146), .A2(n_453), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g517 ( .A1(n_146), .A2(n_453), .B(n_518), .C(n_519), .Y(n_517) );
INVx2_ASAP7_75t_SL g177 ( .A(n_147), .Y(n_177) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_147), .A2(n_469), .B(n_473), .Y(n_468) );
BUFx4f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx3_ASAP7_75t_L g165 ( .A(n_148), .Y(n_165) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_149), .B(n_152), .Y(n_151) );
AND2x4_ASAP7_75t_L g201 ( .A(n_149), .B(n_152), .Y(n_201) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g362 ( .A(n_154), .B(n_318), .Y(n_362) );
AND2x2_ASAP7_75t_L g409 ( .A(n_154), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_163), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
AND2x2_ASAP7_75t_L g272 ( .A(n_156), .B(n_163), .Y(n_272) );
INVx2_ASAP7_75t_L g279 ( .A(n_156), .Y(n_279) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_156), .Y(n_400) );
BUFx3_ASAP7_75t_L g416 ( .A(n_156), .Y(n_416) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_162), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_157), .Y(n_210) );
INVx2_ASAP7_75t_L g241 ( .A(n_163), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_163), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g339 ( .A(n_163), .B(n_279), .Y(n_339) );
INVx1_ASAP7_75t_L g357 ( .A(n_163), .Y(n_357) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_163), .Y(n_373) );
INVx1_ASAP7_75t_L g395 ( .A(n_163), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_163), .B(n_274), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_163), .B(n_228), .Y(n_432) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B(n_172), .Y(n_164) );
INVx4_ASAP7_75t_L g237 ( .A(n_165), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_165), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
INVx1_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_192), .Y(n_174) );
AND2x4_ASAP7_75t_L g246 ( .A(n_175), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
AND2x2_ASAP7_75t_L g262 ( .A(n_175), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g297 ( .A(n_175), .B(n_202), .Y(n_297) );
AND2x2_ASAP7_75t_L g307 ( .A(n_175), .B(n_203), .Y(n_307) );
OR2x2_ASAP7_75t_L g387 ( .A(n_175), .B(n_302), .Y(n_387) );
OAI322xp33_ASAP7_75t_L g417 ( .A1(n_175), .A2(n_330), .A3(n_369), .B1(n_402), .B2(n_418), .C1(n_419), .C2(n_420), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_175), .B(n_400), .Y(n_418) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g251 ( .A(n_176), .Y(n_251) );
AOI21x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_191), .Y(n_176) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_177), .A2(n_459), .B(n_467), .Y(n_458) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_177), .A2(n_459), .B(n_467), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_185), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_180), .A2(n_186), .B1(n_230), .B2(n_232), .Y(n_229) );
INVx1_ASAP7_75t_L g557 ( .A(n_180), .Y(n_557) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_184), .Y(n_180) );
INVx1_ASAP7_75t_L g481 ( .A(n_181), .Y(n_481) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
OR2x6_ASAP7_75t_L g453 ( .A(n_182), .B(n_190), .Y(n_453) );
INVxp33_ASAP7_75t_L g464 ( .A(n_182), .Y(n_464) );
INVx1_ASAP7_75t_L g482 ( .A(n_184), .Y(n_482) );
INVxp67_ASAP7_75t_L g555 ( .A(n_186), .Y(n_555) );
NOR2x1p5_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
INVx1_ASAP7_75t_L g465 ( .A(n_189), .Y(n_465) );
INVx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_192), .A2(n_364), .B1(n_368), .B2(n_371), .Y(n_363) );
AOI211xp5_ASAP7_75t_L g423 ( .A1(n_192), .A2(n_424), .B(n_425), .C(n_428), .Y(n_423) );
AND2x4_ASAP7_75t_SL g192 ( .A(n_193), .B(n_202), .Y(n_192) );
AND2x4_ASAP7_75t_L g245 ( .A(n_193), .B(n_213), .Y(n_245) );
HB1xp67_ASAP7_75t_L g249 ( .A(n_193), .Y(n_249) );
INVx5_ASAP7_75t_L g261 ( .A(n_193), .Y(n_261) );
INVx2_ASAP7_75t_L g270 ( .A(n_193), .Y(n_270) );
AND2x2_ASAP7_75t_L g293 ( .A(n_193), .B(n_203), .Y(n_293) );
AND2x2_ASAP7_75t_L g322 ( .A(n_193), .B(n_212), .Y(n_322) );
OR2x2_ASAP7_75t_L g331 ( .A(n_193), .B(n_251), .Y(n_331) );
OR2x2_ASAP7_75t_L g346 ( .A(n_193), .B(n_260), .Y(n_346) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_201), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_201), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_201), .B(n_233), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_201), .B(n_236), .Y(n_235) );
NOR3xp33_ASAP7_75t_L g238 ( .A(n_201), .B(n_239), .C(n_240), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_201), .A2(n_516), .B(n_520), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_202), .B(n_222), .Y(n_221) );
INVx3_ASAP7_75t_SL g330 ( .A(n_202), .Y(n_330) );
AND2x2_ASAP7_75t_L g353 ( .A(n_202), .B(n_261), .Y(n_353) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_212), .Y(n_202) );
INVx2_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
AND2x2_ASAP7_75t_L g250 ( .A(n_203), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g264 ( .A(n_203), .B(n_213), .Y(n_264) );
INVx1_ASAP7_75t_L g268 ( .A(n_203), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_203), .B(n_213), .Y(n_302) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_203), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_203), .B(n_261), .Y(n_377) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_210), .B(n_211), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_205), .B(n_209), .Y(n_204) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_210), .A2(n_214), .B(n_220), .Y(n_213) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_210), .A2(n_214), .B(n_220), .Y(n_260) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_210), .A2(n_504), .B(n_510), .Y(n_503) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_213), .Y(n_283) );
AND2x2_ASAP7_75t_L g367 ( .A(n_213), .B(n_251), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_226), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_223), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x6_ASAP7_75t_SL g431 ( .A(n_224), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_225), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_225), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g379 ( .A(n_225), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_226), .A2(n_288), .B1(n_291), .B2(n_298), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_227), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_227), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_227), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_227), .B(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
AND2x2_ASAP7_75t_L g273 ( .A(n_228), .B(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g282 ( .A(n_228), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g340 ( .A1(n_228), .A2(n_289), .B1(n_341), .B2(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g348 ( .A(n_228), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_228), .B(n_342), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_228), .B(n_272), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_228), .B(n_279), .Y(n_421) );
AND2x4_ASAP7_75t_L g228 ( .A(n_229), .B(n_234), .Y(n_228) );
INVx3_ASAP7_75t_L g447 ( .A(n_237), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_237), .A2(n_447), .B1(n_545), .B2(n_550), .Y(n_544) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_240), .A2(n_453), .B1(n_493), .B2(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_240), .B(n_548), .Y(n_547) );
OAI21xp33_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_248), .B(n_252), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_246), .Y(n_243) );
NAND4xp25_ASAP7_75t_SL g291 ( .A(n_244), .B(n_292), .C(n_294), .D(n_296), .Y(n_291) );
INVx2_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_245), .B(n_352), .Y(n_381) );
AND2x2_ASAP7_75t_L g408 ( .A(n_245), .B(n_246), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_245), .B(n_268), .Y(n_419) );
INVx1_ASAP7_75t_L g284 ( .A(n_246), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_246), .A2(n_309), .B1(n_320), .B2(n_323), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_246), .B(n_259), .C(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_246), .B(n_261), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_246), .B(n_269), .Y(n_412) );
AND2x2_ASAP7_75t_L g344 ( .A(n_247), .B(n_251), .Y(n_344) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_247), .Y(n_405) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g300 ( .A(n_249), .Y(n_300) );
INVx1_ASAP7_75t_L g390 ( .A(n_250), .Y(n_390) );
AND2x2_ASAP7_75t_L g397 ( .A(n_250), .B(n_261), .Y(n_397) );
BUFx2_ASAP7_75t_L g352 ( .A(n_251), .Y(n_352) );
NAND3xp33_ASAP7_75t_SL g253 ( .A(n_254), .B(n_275), .C(n_287), .Y(n_253) );
OAI31xp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_262), .A3(n_265), .B(n_271), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_255), .A2(n_309), .B1(n_313), .B2(n_314), .Y(n_308) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
OR2x2_ASAP7_75t_L g294 ( .A(n_257), .B(n_295), .Y(n_294) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_257), .B(n_321), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_258), .A2(n_360), .B(n_390), .C(n_391), .Y(n_389) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_259), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_260), .B(n_268), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_260), .B(n_293), .Y(n_313) );
AND2x2_ASAP7_75t_L g430 ( .A(n_263), .B(n_352), .Y(n_430) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g286 ( .A(n_264), .B(n_270), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_269), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_269), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g361 ( .A(n_269), .B(n_344), .Y(n_361) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_270), .B(n_344), .Y(n_350) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g342 ( .A(n_272), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_273), .B(n_373), .Y(n_372) );
AOI32xp33_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_283), .A3(n_284), .B1(n_285), .B2(n_837), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_276), .A2(n_361), .B1(n_397), .B2(n_398), .C(n_401), .Y(n_396) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_279), .Y(n_324) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g289 ( .A(n_281), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g394 ( .A(n_282), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_283), .B(n_305), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g327 ( .A1(n_285), .A2(n_328), .B1(n_332), .B2(n_336), .C(n_340), .Y(n_327) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
OAI211xp5_ASAP7_75t_L g303 ( .A1(n_290), .A2(n_304), .B(n_308), .C(n_319), .Y(n_303) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI322xp33_ASAP7_75t_L g401 ( .A1(n_296), .A2(n_306), .A3(n_355), .B1(n_402), .B2(n_403), .C1(n_404), .C2(n_406), .Y(n_401) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_299), .A2(n_429), .B(n_431), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_305), .A2(n_386), .B(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g427 ( .A(n_312), .B(n_393), .Y(n_427) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVxp67_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_318), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g402 ( .A(n_318), .Y(n_402) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI31xp33_ASAP7_75t_L g358 ( .A1(n_322), .A2(n_359), .A3(n_361), .B(n_362), .Y(n_358) );
NOR2x1_ASAP7_75t_L g325 ( .A(n_326), .B(n_384), .Y(n_325) );
NAND5xp2_ASAP7_75t_L g326 ( .A(n_327), .B(n_347), .C(n_358), .D(n_363), .E(n_374), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_330), .A2(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g398 ( .A(n_334), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B(n_351), .C(n_354), .Y(n_347) );
INVxp33_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
OR2x2_ASAP7_75t_L g376 ( .A(n_352), .B(n_377), .Y(n_376) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_355), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g426 ( .A(n_367), .Y(n_426) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B(n_380), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI21xp33_ASAP7_75t_L g380 ( .A1(n_376), .A2(n_381), .B(n_382), .Y(n_380) );
NAND4xp25_ASAP7_75t_L g384 ( .A(n_385), .B(n_396), .C(n_407), .D(n_423), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_394), .B(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g424 ( .A(n_406), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_411), .B2(n_413), .C(n_417), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_435), .B(n_437), .Y(n_436) );
OR2x6_ASAP7_75t_SL g786 ( .A(n_435), .B(n_787), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_435), .B(n_787), .Y(n_797) );
OR2x2_ASAP7_75t_L g801 ( .A(n_435), .B(n_778), .Y(n_801) );
INVx1_ASAP7_75t_L g777 ( .A(n_436), .Y(n_777) );
INVx2_ASAP7_75t_L g810 ( .A(n_437), .Y(n_810) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_771), .Y(n_437) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_650), .C(n_674), .D(n_740), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_439), .A2(n_674), .B1(n_774), .B2(n_838), .Y(n_775) );
NAND3x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_602), .C(n_636), .Y(n_439) );
NOR3x1_ASAP7_75t_L g440 ( .A(n_441), .B(n_561), .C(n_581), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_442), .B(n_536), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_474), .B1(n_525), .B2(n_533), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_456), .Y(n_443) );
AND2x2_ASAP7_75t_L g700 ( .A(n_444), .B(n_630), .Y(n_700) );
INVx1_ASAP7_75t_L g707 ( .A(n_444), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_444), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_444), .B(n_570), .Y(n_759) );
OR2x2_ASAP7_75t_L g769 ( .A(n_444), .B(n_770), .Y(n_769) );
INVx3_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_445), .B(n_527), .Y(n_590) );
AND2x4_ASAP7_75t_L g618 ( .A(n_445), .B(n_532), .Y(n_618) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g566 ( .A(n_446), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_446), .B(n_458), .Y(n_656) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_446), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_446), .B(n_543), .Y(n_693) );
AO21x2_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_455), .Y(n_446) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_447), .A2(n_448), .B(n_455), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g488 ( .A(n_453), .Y(n_488) );
INVxp67_ASAP7_75t_L g546 ( .A(n_453), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_456), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g764 ( .A(n_456), .B(n_601), .Y(n_764) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g754 ( .A(n_457), .B(n_693), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
INVx2_ASAP7_75t_L g532 ( .A(n_458), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_460), .B(n_466), .Y(n_459) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
INVx2_ASAP7_75t_L g542 ( .A(n_468), .Y(n_542) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_468), .Y(n_567) );
INVx1_ASAP7_75t_L g580 ( .A(n_468), .Y(n_580) );
INVxp67_ASAP7_75t_L g599 ( .A(n_468), .Y(n_599) );
AND2x4_ASAP7_75t_L g630 ( .A(n_468), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_511), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_501), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g672 ( .A(n_477), .B(n_659), .Y(n_672) );
AND2x2_ASAP7_75t_L g696 ( .A(n_477), .B(n_512), .Y(n_696) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_489), .Y(n_477) );
INVx2_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_478), .Y(n_539) );
INVx1_ASAP7_75t_L g596 ( .A(n_478), .Y(n_596) );
AND2x4_ASAP7_75t_L g605 ( .A(n_478), .B(n_523), .Y(n_605) );
AND2x2_ASAP7_75t_L g661 ( .A(n_478), .B(n_513), .Y(n_661) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_484), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .C(n_483), .Y(n_480) );
INVx3_ASAP7_75t_L g523 ( .A(n_489), .Y(n_523) );
AND2x2_ASAP7_75t_L g535 ( .A(n_489), .B(n_503), .Y(n_535) );
INVx2_ASAP7_75t_L g574 ( .A(n_489), .Y(n_574) );
NOR2x1_ASAP7_75t_SL g587 ( .A(n_489), .B(n_513), .Y(n_587) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .B(n_500), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_496), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g689 ( .A(n_501), .Y(n_689) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g612 ( .A(n_502), .Y(n_612) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_503), .Y(n_570) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_503), .Y(n_586) );
AND2x2_ASAP7_75t_L g594 ( .A(n_503), .B(n_523), .Y(n_594) );
INVx1_ASAP7_75t_L g634 ( .A(n_503), .Y(n_634) );
INVx1_ASAP7_75t_L g659 ( .A(n_503), .Y(n_659) );
OR2x2_ASAP7_75t_L g720 ( .A(n_503), .B(n_513), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
OA211x2_ASAP7_75t_L g741 ( .A1(n_511), .A2(n_742), .B(n_744), .C(n_751), .Y(n_741) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_521), .Y(n_511) );
AND2x2_ASAP7_75t_L g662 ( .A(n_512), .B(n_535), .Y(n_662) );
AND2x2_ASAP7_75t_SL g680 ( .A(n_512), .B(n_522), .Y(n_680) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g534 ( .A(n_513), .Y(n_534) );
INVx2_ASAP7_75t_L g576 ( .A(n_513), .Y(n_576) );
AND2x4_ASAP7_75t_L g639 ( .A(n_513), .B(n_596), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_513), .B(n_635), .Y(n_690) );
AND2x2_ASAP7_75t_L g733 ( .A(n_513), .B(n_574), .Y(n_733) );
OR2x6_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_522), .B(n_634), .Y(n_727) );
AND2x2_ASAP7_75t_L g747 ( .A(n_522), .B(n_570), .Y(n_747) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g635 ( .A(n_523), .Y(n_635) );
INVx1_ASAP7_75t_L g609 ( .A(n_524), .Y(n_609) );
NOR2xp67_ASAP7_75t_SL g525 ( .A(n_526), .B(n_529), .Y(n_525) );
INVx1_ASAP7_75t_L g703 ( .A(n_526), .Y(n_703) );
NOR2xp67_ASAP7_75t_L g750 ( .A(n_526), .B(n_704), .Y(n_750) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g723 ( .A(n_528), .B(n_565), .Y(n_723) );
OAI211xp5_ASAP7_75t_L g711 ( .A1(n_529), .A2(n_712), .B(n_715), .C(n_724), .Y(n_711) );
A2O1A1Ixp33_ASAP7_75t_L g755 ( .A1(n_529), .A2(n_749), .B(n_756), .C(n_760), .Y(n_755) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g640 ( .A(n_530), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g559 ( .A(n_531), .Y(n_559) );
NOR2x1_ASAP7_75t_L g579 ( .A(n_531), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g615 ( .A(n_531), .B(n_565), .Y(n_615) );
NOR2xp67_ASAP7_75t_L g725 ( .A(n_531), .B(n_565), .Y(n_725) );
AND2x2_ASAP7_75t_L g598 ( .A(n_532), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g649 ( .A(n_532), .Y(n_649) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x4_ASAP7_75t_SL g538 ( .A(n_534), .B(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g595 ( .A(n_534), .B(n_596), .Y(n_595) );
NOR2x1_ASAP7_75t_L g624 ( .A(n_534), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g643 ( .A(n_534), .B(n_644), .Y(n_643) );
NOR2xp67_ASAP7_75t_SL g726 ( .A(n_534), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_SL g537 ( .A(n_535), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_535), .B(n_608), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_540), .Y(n_536) );
INVx2_ASAP7_75t_SL g734 ( .A(n_540), .Y(n_734) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_558), .Y(n_540) );
INVx3_ASAP7_75t_L g657 ( .A(n_541), .Y(n_657) );
AND2x2_ASAP7_75t_L g678 ( .A(n_541), .B(n_669), .Y(n_678) );
AND2x2_ASAP7_75t_L g736 ( .A(n_541), .B(n_618), .Y(n_736) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx2_ASAP7_75t_L g565 ( .A(n_543), .Y(n_565) );
INVx1_ASAP7_75t_L g601 ( .A(n_543), .Y(n_601) );
INVx1_ASAP7_75t_L g621 ( .A(n_543), .Y(n_621) );
OR2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_551), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVxp67_ASAP7_75t_L g704 ( .A(n_558), .Y(n_704) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g564 ( .A(n_560), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g631 ( .A(n_560), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_568), .B1(n_571), .B2(n_577), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
AND2x2_ASAP7_75t_L g578 ( .A(n_564), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g589 ( .A(n_564), .Y(n_589) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g638 ( .A(n_569), .B(n_639), .Y(n_638) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g658 ( .A(n_573), .B(n_659), .Y(n_658) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g666 ( .A(n_574), .Y(n_666) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g714 ( .A(n_576), .B(n_605), .Y(n_714) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_578), .A2(n_672), .B(n_673), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_588), .B(n_591), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_587), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g637 ( .A(n_587), .B(n_611), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_588), .A2(n_695), .B1(n_697), .B2(n_699), .Y(n_694) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_597), .Y(n_591) );
INVxp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_SL g644 ( .A(n_594), .Y(n_644) );
AND2x2_ASAP7_75t_L g673 ( .A(n_595), .B(n_611), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_595), .B(n_633), .Y(n_705) );
AND2x2_ASAP7_75t_L g709 ( .A(n_595), .B(n_666), .Y(n_709) );
OAI21xp5_ASAP7_75t_SL g653 ( .A1(n_597), .A2(n_654), .B(n_658), .Y(n_653) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_L g614 ( .A(n_598), .B(n_615), .Y(n_614) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_598), .B(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_SL g683 ( .A(n_601), .Y(n_683) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_626), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_613), .B1(n_616), .B2(n_622), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx4_ASAP7_75t_L g625 ( .A(n_605), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_605), .B(n_611), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_605), .B(n_758), .Y(n_757) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_608), .A2(n_632), .B(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g731 ( .A(n_608), .B(n_633), .Y(n_731) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g713 ( .A(n_610), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g749 ( .A(n_611), .B(n_733), .Y(n_749) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g629 ( .A(n_615), .B(n_630), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_615), .B(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_SL g626 ( .A1(n_616), .A2(n_627), .B1(n_628), .B2(n_632), .Y(n_626) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g743 ( .A(n_620), .B(n_630), .Y(n_743) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g641 ( .A(n_621), .Y(n_641) );
AND2x2_ASAP7_75t_L g667 ( .A(n_621), .B(n_630), .Y(n_667) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_623), .B(n_764), .Y(n_763) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_624), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g718 ( .A(n_625), .Y(n_718) );
INVx1_ASAP7_75t_L g730 ( .A(n_627), .Y(n_730) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_629), .A2(n_673), .B1(n_752), .B2(n_753), .Y(n_751) );
AND2x2_ASAP7_75t_L g668 ( .A(n_630), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g739 ( .A(n_630), .B(n_692), .Y(n_739) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI211xp5_ASAP7_75t_SL g642 ( .A1(n_633), .A2(n_643), .B(n_645), .C(n_646), .Y(n_642) );
AND2x2_ASAP7_75t_SL g752 ( .A(n_633), .B(n_639), .Y(n_752) );
AND2x4_ASAP7_75t_SL g633 ( .A(n_634), .B(n_635), .Y(n_633) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_634), .Y(n_686) );
O2A1O1Ixp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_638), .B(n_640), .C(n_642), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_637), .A2(n_665), .B1(n_667), .B2(n_668), .Y(n_664) );
INVx2_ASAP7_75t_L g645 ( .A(n_639), .Y(n_645) );
AND2x2_ASAP7_75t_L g665 ( .A(n_639), .B(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_639), .Y(n_732) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVxp67_ASAP7_75t_L g773 ( .A(n_651), .Y(n_773) );
NOR2x1_ASAP7_75t_SL g651 ( .A(n_652), .B(n_663), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_660), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_654), .A2(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g684 ( .A(n_656), .Y(n_684) );
INVx1_ASAP7_75t_L g760 ( .A(n_657), .Y(n_760) );
AND2x2_ASAP7_75t_L g698 ( .A(n_661), .B(n_686), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_662), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g663 ( .A(n_664), .B(n_671), .Y(n_663) );
AND2x2_ASAP7_75t_L g765 ( .A(n_667), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
NAND2x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_710), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_694), .C(n_701), .Y(n_675) );
OAI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B1(n_681), .B2(n_685), .C1(n_687), .C2(n_691), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g737 ( .A(n_696), .Y(n_737) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .B1(n_706), .B2(n_708), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp67_ASAP7_75t_SL g710 ( .A(n_711), .B(n_728), .Y(n_710) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_721), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_718), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g770 ( .A(n_723), .Y(n_770) );
NAND2xp33_ASAP7_75t_SL g724 ( .A(n_725), .B(n_726), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_734), .B1(n_735), .B2(n_737), .C(n_738), .Y(n_728) );
NOR4xp25_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .C(n_732), .D(n_733), .Y(n_729) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OAI21xp5_ASAP7_75t_L g772 ( .A1(n_740), .A2(n_773), .B(n_774), .Y(n_772) );
NAND4xp75_ASAP7_75t_L g740 ( .A(n_741), .B(n_755), .C(n_761), .D(n_767), .Y(n_740) );
INVx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_745), .B(n_750), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVxp67_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_778), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_780), .B(n_781), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_789), .B(n_790), .Y(n_782) );
INVxp33_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND2x1_ASAP7_75t_SL g784 ( .A(n_785), .B(n_788), .Y(n_784) );
CKINVDCx11_ASAP7_75t_R g785 ( .A(n_786), .Y(n_785) );
OR3x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_798), .C(n_802), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_791), .A2(n_806), .B(n_809), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
BUFx3_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_R g808 ( .A(n_797), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
BUFx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_820), .Y(n_804) );
INVx1_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
INVx1_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
XNOR2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_815), .B1(n_816), .B2(n_819), .Y(n_811) );
INVx1_ASAP7_75t_L g819 ( .A(n_812), .Y(n_819) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
CKINVDCx11_ASAP7_75t_R g821 ( .A(n_822), .Y(n_821) );
CKINVDCx8_ASAP7_75t_R g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
INVx3_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_SL g835 ( .A(n_827), .Y(n_835) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_828), .B(n_832), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
endmodule