module fake_jpeg_8598_n_313 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_313);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_313;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_21),
.A2(n_32),
.B(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_44),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_31),
.B1(n_27),
.B2(n_32),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_51),
.B1(n_60),
.B2(n_65),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_31),
.B1(n_27),
.B2(n_23),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_56),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_37),
.A2(n_31),
.B1(n_27),
.B2(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_33),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_27),
.B1(n_24),
.B2(n_35),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_68),
.A2(n_71),
.B1(n_97),
.B2(n_34),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_39),
.B1(n_19),
.B2(n_21),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_82),
.B1(n_89),
.B2(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_39),
.B1(n_41),
.B2(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_33),
.B1(n_35),
.B2(n_23),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_85),
.B(n_100),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_25),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_41),
.Y(n_78)
);

AO22x2_ASAP7_75t_L g120 ( 
.A1(n_78),
.A2(n_59),
.B1(n_55),
.B2(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_41),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_79),
.B(n_54),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_22),
.B1(n_34),
.B2(n_26),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_81),
.B(n_84),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_20),
.B1(n_17),
.B2(n_30),
.Y(n_82)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_46),
.B(n_20),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_42),
.B(n_47),
.Y(n_104)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_58),
.A2(n_63),
.B1(n_49),
.B2(n_62),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_17),
.B1(n_28),
.B2(n_30),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_20),
.B1(n_17),
.B2(n_30),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_67),
.B1(n_34),
.B2(n_28),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_25),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_25),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_64),
.B(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_59),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_45),
.A2(n_30),
.B1(n_28),
.B2(n_64),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_64),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_100)
);

CKINVDCx6p67_ASAP7_75t_R g101 ( 
.A(n_46),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_28),
.B1(n_22),
.B2(n_26),
.Y(n_102)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_40),
.B(n_34),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_108),
.B(n_86),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_109),
.A2(n_120),
.B1(n_97),
.B2(n_77),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_110),
.B(n_40),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_0),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_0),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_117),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_122),
.C(n_89),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_94),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_71),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_128),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_55),
.C(n_40),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_126),
.B1(n_91),
.B2(n_93),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_1),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_68),
.C(n_70),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_141),
.C(n_142),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_134),
.A2(n_146),
.B1(n_153),
.B2(n_120),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_136),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_139),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_68),
.B1(n_75),
.B2(n_83),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_155),
.B(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_70),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_143),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_86),
.C(n_77),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_147),
.B(n_149),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_106),
.A2(n_83),
.B(n_98),
.Y(n_147)
);

NAND2x1p5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_78),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_104),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_150),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_99),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_78),
.B1(n_93),
.B2(n_94),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_101),
.C(n_78),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_124),
.C(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_74),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_159),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_1),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_81),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_170),
.B1(n_186),
.B2(n_190),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_168),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_153),
.A2(n_122),
.B1(n_123),
.B2(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_173),
.C(n_179),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_114),
.C(n_107),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_140),
.B1(n_158),
.B2(n_156),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_174),
.A2(n_103),
.B1(n_162),
.B2(n_25),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_107),
.B(n_125),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_175),
.A2(n_177),
.B(n_188),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_131),
.A2(n_105),
.B(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_117),
.C(n_130),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_109),
.C(n_113),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_184),
.Y(n_216)
);

OAI32xp33_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_113),
.A3(n_126),
.B1(n_22),
.B2(n_127),
.Y(n_182)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_40),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_93),
.B1(n_129),
.B2(n_115),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_40),
.B(n_94),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_129),
.B1(n_88),
.B2(n_87),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_132),
.B(n_25),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_160),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_134),
.B1(n_147),
.B2(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_136),
.A2(n_87),
.B1(n_88),
.B2(n_118),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_145),
.A2(n_118),
.B1(n_127),
.B2(n_22),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_194),
.A2(n_118),
.B1(n_152),
.B2(n_103),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_133),
.B(n_81),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_155),
.Y(n_202)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_151),
.C(n_133),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_205),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_198),
.A2(n_199),
.B(n_217),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g199 ( 
.A(n_185),
.B(n_144),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_167),
.C(n_172),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_161),
.C(n_157),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_212),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_152),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_207),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_152),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_143),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_220),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_163),
.B(n_175),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_169),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_2),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_8),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_222),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_165),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_228),
.C(n_242),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_167),
.C(n_173),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_164),
.B1(n_185),
.B2(n_170),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_234),
.B1(n_238),
.B2(n_240),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_201),
.A2(n_189),
.B1(n_169),
.B2(n_192),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_237),
.A2(n_203),
.B(n_206),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_222),
.A2(n_178),
.B1(n_182),
.B2(n_163),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_201),
.A2(n_178),
.B1(n_186),
.B2(n_180),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_171),
.C(n_184),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_172),
.B1(n_194),
.B2(n_188),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_197),
.B1(n_206),
.B2(n_200),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_202),
.C(n_218),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_199),
.C(n_209),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_257),
.B1(n_243),
.B2(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_250),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_253),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_205),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_225),
.A2(n_218),
.B(n_197),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_228),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_252),
.A2(n_261),
.B1(n_233),
.B2(n_232),
.Y(n_268)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_235),
.B(n_215),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_211),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_260),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_200),
.B1(n_199),
.B2(n_198),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_220),
.B(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_258),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_256),
.C(n_254),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_215),
.B(n_194),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_236),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_233),
.B1(n_231),
.B2(n_235),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_263),
.A2(n_268),
.B1(n_249),
.B2(n_257),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g264 ( 
.A(n_261),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_270),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_259),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_224),
.C(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_226),
.C(n_229),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_229),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_281),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_273),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_269),
.Y(n_290)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_247),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_286),
.B(n_287),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_239),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_265),
.A2(n_251),
.B1(n_245),
.B2(n_169),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_246),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.C(n_294),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_284),
.B1(n_277),
.B2(n_288),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_279),
.A2(n_274),
.B(n_275),
.Y(n_294)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_194),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_282),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_271),
.B(n_269),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_296),
.A2(n_16),
.B(n_12),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_9),
.B(n_15),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g306 ( 
.A1(n_298),
.A2(n_299),
.B(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_278),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_283),
.B(n_217),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_302),
.A2(n_303),
.A3(n_304),
.B1(n_298),
.B2(n_297),
.C1(n_10),
.C2(n_11),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_16),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_307),
.B1(n_308),
.B2(n_7),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_293),
.A3(n_290),
.B1(n_11),
.B2(n_10),
.C1(n_9),
.C2(n_2),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_308)
);

AOI321xp33_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_310),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_306),
.A2(n_2),
.B(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_5),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_6),
.Y(n_313)
);


endmodule