module fake_ariane_2499_n_1861 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1861);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1861;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_699;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_108),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_71),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_85),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_38),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_82),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_154),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_56),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_54),
.Y(n_198)
);

BUFx2_ASAP7_75t_SL g199 ( 
.A(n_39),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_55),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_52),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_24),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_3),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_6),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_49),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_43),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_23),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_77),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_52),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_120),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_92),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_147),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_37),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_56),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_2),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_13),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_157),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_133),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_12),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_14),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_70),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_105),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_19),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_149),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_113),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_75),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_8),
.Y(n_240)
);

BUFx8_ASAP7_75t_SL g241 ( 
.A(n_68),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_168),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_148),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_31),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_174),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_33),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_33),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_83),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_90),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_166),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_121),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_103),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_24),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_158),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_137),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_123),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_146),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_170),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_73),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_20),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_74),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_40),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_104),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_173),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_66),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_36),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_98),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_163),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_23),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_109),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_111),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_88),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_165),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_93),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_37),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_62),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_64),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_29),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_78),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_43),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_117),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_40),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_87),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_132),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_143),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_97),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_51),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_95),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_50),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_7),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_155),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_55),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_39),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_60),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_67),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_127),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_94),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_138),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_20),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_21),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_161),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_140),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_116),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_44),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_91),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_131),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_10),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_42),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_34),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_171),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_102),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_10),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_69),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_50),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_17),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_4),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_49),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_26),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_32),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_1),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_2),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_17),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_89),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_162),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_72),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_47),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_79),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_0),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_53),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_51),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_135),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_27),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_164),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_35),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_47),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_35),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_99),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_31),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_107),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_59),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_169),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_124),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_126),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_114),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_285),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_285),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_196),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_1),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_241),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_183),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_238),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_258),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_271),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_322),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_318),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_199),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_318),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_205),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_209),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_224),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_215),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_194),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_324),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_306),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_300),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_216),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_269),
.B(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_217),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_219),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_197),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_225),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_326),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_344),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_184),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_227),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_328),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_344),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_186),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_344),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_344),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_232),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_232),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_236),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_298),
.B(n_5),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_240),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_298),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_330),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_186),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_186),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_250),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_223),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_330),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_187),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_316),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_187),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_265),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_268),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_197),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_211),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_211),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_184),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_223),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_317),
.B(n_5),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_317),
.B(n_7),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_280),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_272),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_181),
.B(n_9),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_177),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_184),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_207),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_198),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_280),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_180),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_191),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_223),
.B(n_11),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_192),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_189),
.B(n_11),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_198),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_275),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_357),
.B(n_234),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_226),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_355),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_373),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_361),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_361),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_403),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_193),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_354),
.A2(n_204),
.B(n_203),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_356),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_356),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_380),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_417),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_234),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_359),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_370),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_190),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_417),
.B(n_206),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_210),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_234),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_377),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_377),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_362),
.Y(n_476)
);

OA21x2_ASAP7_75t_L g477 ( 
.A1(n_381),
.A2(n_218),
.B(n_214),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_419),
.B(n_221),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_382),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g481 ( 
.A1(n_382),
.A2(n_392),
.B(n_387),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_376),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_395),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_423),
.B(n_222),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_395),
.A2(n_244),
.B(n_242),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_190),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_424),
.A2(n_251),
.B(n_248),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_438),
.B(n_177),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g498 ( 
.A1(n_424),
.A2(n_264),
.B(n_255),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_429),
.B(n_274),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_438),
.B(n_245),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_404),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_436),
.B(n_319),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_397),
.A2(n_321),
.B1(n_337),
.B2(n_329),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_436),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_440),
.B(n_319),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_405),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_440),
.B(n_249),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_371),
.B(n_213),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_408),
.B(n_350),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_405),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_360),
.B(n_350),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_380),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_406),
.B(n_284),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_410),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_408),
.B(n_262),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_410),
.B(n_267),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_481),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_383),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_516),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_445),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_481),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_512),
.A2(n_386),
.B1(n_431),
.B2(n_439),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_512),
.A2(n_442),
.B1(n_427),
.B2(n_428),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_481),
.Y(n_531)
);

OR2x6_ASAP7_75t_L g532 ( 
.A(n_461),
.B(n_425),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_481),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_433),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_474),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_467),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_457),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_445),
.B(n_390),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_516),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_461),
.B(n_383),
.Y(n_541)
);

AND2x6_ASAP7_75t_L g542 ( 
.A(n_473),
.B(n_212),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_457),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_457),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_512),
.A2(n_422),
.B1(n_435),
.B2(n_331),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_445),
.B(n_364),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_516),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_463),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_467),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_467),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_467),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_514),
.B(n_374),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_448),
.B(n_378),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_516),
.B(n_379),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_512),
.A2(n_290),
.B1(n_315),
.B2(n_345),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_516),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_478),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_473),
.B(n_411),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_473),
.B(n_385),
.Y(n_561)
);

BUFx10_ASAP7_75t_L g562 ( 
.A(n_511),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_511),
.B(n_388),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_478),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_494),
.B(n_416),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_478),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_474),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_459),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_478),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_459),
.Y(n_570)
);

BUFx6f_ASAP7_75t_SL g571 ( 
.A(n_519),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_494),
.B(n_416),
.Y(n_572)
);

NOR2x1p5_ASAP7_75t_L g573 ( 
.A(n_444),
.B(n_363),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_444),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_459),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_444),
.B(n_389),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_448),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_516),
.B(n_391),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_516),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_482),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_472),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_485),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_446),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_482),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_463),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_472),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_516),
.B(n_398),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_474),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_482),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_474),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_482),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_508),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_446),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_453),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_453),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_508),
.B(n_407),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_494),
.B(n_434),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_L g600 ( 
.A(n_507),
.B(n_409),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_455),
.Y(n_601)
);

AO21x2_ASAP7_75t_L g602 ( 
.A1(n_491),
.A2(n_304),
.B(n_302),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_458),
.B(n_414),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_455),
.Y(n_604)
);

OAI21xp33_ASAP7_75t_SL g605 ( 
.A1(n_501),
.A2(n_286),
.B(n_279),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_474),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_512),
.A2(n_415),
.B1(n_401),
.B2(n_426),
.Y(n_608)
);

BUFx6f_ASAP7_75t_SL g609 ( 
.A(n_519),
.Y(n_609)
);

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_476),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_476),
.B(n_420),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_456),
.Y(n_612)
);

BUFx4f_ASAP7_75t_L g613 ( 
.A(n_454),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_485),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_493),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_446),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_454),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_508),
.B(n_421),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_474),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_508),
.B(n_430),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_519),
.A2(n_413),
.B1(n_412),
.B2(n_327),
.Y(n_621)
);

BUFx10_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_464),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_452),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_474),
.Y(n_625)
);

INVxp67_ASAP7_75t_SL g626 ( 
.A(n_452),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_493),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_490),
.B(n_443),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_490),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_458),
.B(n_365),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_454),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_460),
.B(n_207),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_474),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_504),
.B(n_367),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_490),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_469),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_504),
.B(n_368),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_519),
.B(n_176),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

NAND3xp33_ASAP7_75t_L g641 ( 
.A(n_454),
.B(n_231),
.C(n_320),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_490),
.B(n_239),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_493),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_SL g644 ( 
.A(n_506),
.B(n_200),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_493),
.Y(n_645)
);

OAI21xp33_ASAP7_75t_SL g646 ( 
.A1(n_501),
.A2(n_338),
.B(n_256),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_519),
.A2(n_230),
.B1(n_207),
.B2(n_273),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_490),
.B(n_176),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_505),
.B(n_283),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_469),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_505),
.B(n_336),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_493),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_501),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_507),
.B(n_178),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_510),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_504),
.B(n_366),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_475),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_470),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_466),
.A2(n_369),
.B1(n_393),
.B2(n_384),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_470),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_447),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_505),
.A2(n_282),
.B1(n_295),
.B2(n_288),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_504),
.B(n_466),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_465),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_454),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_460),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_480),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_460),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_505),
.B(n_178),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_446),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_480),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_460),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_460),
.B(n_200),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_483),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_624),
.B(n_505),
.Y(n_675)
);

AO221x1_ASAP7_75t_L g676 ( 
.A1(n_644),
.A2(n_212),
.B1(n_289),
.B2(n_507),
.C(n_333),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_626),
.B(n_507),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_661),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_640),
.A2(n_323),
.B1(n_343),
.B2(n_341),
.C(n_339),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_611),
.B(n_321),
.C(n_312),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_661),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_574),
.A2(n_510),
.B1(n_520),
.B2(n_507),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_546),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_596),
.Y(n_684)
);

A2O1A1Ixp33_ASAP7_75t_L g685 ( 
.A1(n_563),
.A2(n_498),
.B(n_491),
.C(n_521),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_574),
.B(n_520),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_622),
.B(n_491),
.Y(n_687)
);

AO221x1_ASAP7_75t_L g688 ( 
.A1(n_621),
.A2(n_289),
.B1(n_212),
.B2(n_352),
.C(n_349),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_546),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_596),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_526),
.B(n_520),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_599),
.B(n_520),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_597),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_561),
.B(n_468),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_597),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_594),
.B(n_520),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_599),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_622),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_601),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_594),
.B(n_521),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_622),
.B(n_498),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_601),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_630),
.B(n_521),
.Y(n_703)
);

INVxp33_ASAP7_75t_L g704 ( 
.A(n_553),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_577),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_622),
.B(n_562),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_539),
.B(n_582),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_539),
.B(n_548),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_541),
.B(n_468),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_630),
.B(n_518),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_604),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_532),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_661),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_576),
.A2(n_340),
.B1(n_182),
.B2(n_185),
.Y(n_714)
);

CKINVDCx14_ASAP7_75t_R g715 ( 
.A(n_553),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_663),
.A2(n_498),
.B(n_479),
.C(n_488),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_560),
.B(n_518),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_653),
.B(n_399),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_585),
.B(n_517),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_560),
.B(n_471),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_562),
.B(n_179),
.Y(n_721)
);

AND2x2_ASAP7_75t_SL g722 ( 
.A(n_613),
.B(n_454),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_655),
.B(n_517),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_542),
.B(n_471),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_542),
.B(n_479),
.Y(n_725)
);

NOR2x1p5_ASAP7_75t_L g726 ( 
.A(n_534),
.B(n_598),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_614),
.Y(n_727)
);

A2O1A1Ixp33_ASAP7_75t_L g728 ( 
.A1(n_552),
.A2(n_605),
.B(n_613),
.C(n_523),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_664),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_562),
.B(n_499),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_562),
.B(n_179),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_604),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_656),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_532),
.B(n_297),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_607),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_542),
.B(n_509),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_666),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_532),
.B(n_301),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_607),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_534),
.B(n_509),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_542),
.B(n_509),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_542),
.B(n_509),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_612),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_666),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_612),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_532),
.B(n_307),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_537),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_636),
.B(n_182),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_636),
.B(n_185),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_636),
.B(n_188),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_537),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_532),
.B(n_308),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_618),
.B(n_620),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_629),
.B(n_672),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_565),
.B(n_513),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_613),
.A2(n_477),
.B1(n_489),
.B2(n_515),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_666),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_L g758 ( 
.A(n_535),
.B(n_188),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_623),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_605),
.A2(n_477),
.B1(n_489),
.B2(n_513),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_565),
.B(n_572),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_623),
.Y(n_762)
);

INVx4_ASAP7_75t_SL g763 ( 
.A(n_571),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_534),
.B(n_608),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_530),
.A2(n_312),
.B1(n_323),
.B2(n_325),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_627),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_636),
.B(n_195),
.Y(n_767)
);

INVxp33_ASAP7_75t_L g768 ( 
.A(n_631),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_572),
.B(n_513),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_635),
.B(n_513),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_638),
.B(n_515),
.Y(n_771)
);

AO221x1_ASAP7_75t_L g772 ( 
.A1(n_659),
.A2(n_212),
.B1(n_289),
.B2(n_334),
.C(n_451),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_633),
.B(n_515),
.Y(n_773)
);

O2A1O1Ixp5_ASAP7_75t_L g774 ( 
.A1(n_554),
.A2(n_515),
.B(n_495),
.C(n_500),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_549),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_637),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_633),
.B(n_325),
.Y(n_777)
);

INVx2_ASAP7_75t_SL g778 ( 
.A(n_573),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_668),
.B(n_329),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_600),
.A2(n_202),
.B1(n_201),
.B2(n_195),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_535),
.B(n_201),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_617),
.A2(n_477),
.B1(n_489),
.B2(n_500),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_549),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_617),
.A2(n_477),
.B1(n_489),
.B2(n_497),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_642),
.B(n_477),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_535),
.B(n_202),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_580),
.B(n_311),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_673),
.B(n_603),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_580),
.B(n_311),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_610),
.Y(n_790)
);

AO221x1_ASAP7_75t_L g791 ( 
.A1(n_522),
.A2(n_212),
.B1(n_289),
.B2(n_647),
.C(n_567),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_649),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_673),
.B(n_545),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_538),
.A2(n_591),
.B(n_586),
.C(n_581),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_637),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_650),
.Y(n_796)
);

NOR3xp33_ASAP7_75t_L g797 ( 
.A(n_648),
.B(n_335),
.C(n_337),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_651),
.B(n_477),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_529),
.B(n_662),
.C(n_654),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_573),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_639),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_650),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_668),
.B(n_335),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_658),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_668),
.B(n_339),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_658),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_571),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_660),
.B(n_483),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_588),
.B(n_489),
.Y(n_809)
);

INVx4_ASAP7_75t_SL g810 ( 
.A(n_571),
.Y(n_810)
);

AOI22xp5_ASAP7_75t_L g811 ( 
.A1(n_609),
.A2(n_313),
.B1(n_314),
.B2(n_332),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_669),
.B(n_341),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_580),
.B(n_489),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_609),
.A2(n_313),
.B1(n_314),
.B2(n_332),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_550),
.B(n_484),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_551),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_609),
.B(n_343),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_551),
.B(n_558),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_617),
.A2(n_340),
.B1(n_346),
.B2(n_348),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_558),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_559),
.B(n_564),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_559),
.B(n_484),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_555),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_617),
.B(n_347),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_632),
.A2(n_346),
.B1(n_348),
.B2(n_351),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_660),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_564),
.B(n_486),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_632),
.B(n_347),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_566),
.B(n_486),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_667),
.A2(n_495),
.B1(n_497),
.B2(n_351),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_667),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_671),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_566),
.B(n_353),
.Y(n_833)
);

BUFx5_ASAP7_75t_L g834 ( 
.A(n_527),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_569),
.B(n_353),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_632),
.B(n_14),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_522),
.B(n_632),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_671),
.A2(n_502),
.B(n_496),
.C(n_492),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_569),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_674),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

OR2x2_ASAP7_75t_L g842 ( 
.A(n_707),
.B(n_674),
.Y(n_842)
);

NOR3xp33_ASAP7_75t_L g843 ( 
.A(n_790),
.B(n_646),
.C(n_578),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_718),
.B(n_723),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_694),
.B(n_527),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_694),
.B(n_528),
.Y(n_846)
);

NOR3xp33_ASAP7_75t_L g847 ( 
.A(n_679),
.B(n_543),
.C(n_538),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_837),
.A2(n_568),
.B(n_544),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_709),
.B(n_528),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_837),
.A2(n_522),
.B(n_531),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_687),
.A2(n_568),
.B(n_544),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_687),
.A2(n_701),
.B(n_818),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_754),
.B(n_665),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_701),
.A2(n_821),
.B(n_794),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_709),
.B(n_531),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_716),
.A2(n_522),
.B(n_533),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_754),
.B(n_665),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_809),
.A2(n_730),
.B(n_677),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_728),
.A2(n_593),
.B(n_584),
.C(n_652),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_730),
.B(n_533),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_684),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_708),
.B(n_524),
.Y(n_862)
);

AND2x4_ASAP7_75t_L g863 ( 
.A(n_763),
.B(n_524),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_813),
.A2(n_753),
.B(n_675),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_683),
.B(n_665),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_689),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_753),
.A2(n_586),
.B(n_570),
.Y(n_867)
);

O2A1O1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_765),
.A2(n_643),
.B(n_645),
.C(n_628),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_R g869 ( 
.A(n_727),
.B(n_570),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_799),
.A2(n_581),
.B1(n_591),
.B2(n_575),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_678),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_726),
.A2(n_665),
.B1(n_575),
.B2(n_641),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_700),
.A2(n_525),
.B(n_556),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_719),
.Y(n_874)
);

OAI22xp5_ASAP7_75t_L g875 ( 
.A1(n_690),
.A2(n_693),
.B1(n_699),
.B2(n_695),
.Y(n_875)
);

AOI33xp33_ASAP7_75t_L g876 ( 
.A1(n_697),
.A2(n_587),
.A3(n_590),
.B1(n_584),
.B2(n_593),
.B3(n_652),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_681),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_712),
.B(n_289),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_713),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_763),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_703),
.A2(n_525),
.B(n_557),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_710),
.A2(n_525),
.B(n_557),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_720),
.B(n_590),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_815),
.A2(n_556),
.B(n_525),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_702),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_836),
.A2(n_615),
.B(n_628),
.C(n_645),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_685),
.A2(n_641),
.B(n_643),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_779),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_755),
.A2(n_567),
.B(n_657),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_680),
.B(n_592),
.C(n_657),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_769),
.A2(n_567),
.B(n_657),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_740),
.B(n_536),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_822),
.A2(n_567),
.B(n_657),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_838),
.A2(n_589),
.B(n_634),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_827),
.A2(n_536),
.B(n_634),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_792),
.B(n_536),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_729),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_761),
.B(n_536),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_SL g899 ( 
.A(n_704),
.B(n_220),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_777),
.B(n_602),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_829),
.A2(n_606),
.B(n_634),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_773),
.A2(n_606),
.B(n_634),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_692),
.B(n_589),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_706),
.A2(n_625),
.B(n_619),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_737),
.B(n_540),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_770),
.B(n_771),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_691),
.B(n_589),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_793),
.B(n_602),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_778),
.B(n_589),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_711),
.A2(n_606),
.B1(n_625),
.B2(n_619),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_682),
.B(n_592),
.Y(n_911)
);

NOR2x1p5_ASAP7_75t_SL g912 ( 
.A(n_834),
.B(n_465),
.Y(n_912)
);

OR2x6_ASAP7_75t_L g913 ( 
.A(n_712),
.B(n_579),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_SL g914 ( 
.A1(n_706),
.A2(n_606),
.B(n_625),
.C(n_619),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_717),
.B(n_592),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_732),
.A2(n_592),
.B1(n_625),
.B2(n_619),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_836),
.A2(n_540),
.B(n_547),
.C(n_670),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_686),
.B(n_583),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_737),
.B(n_744),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_696),
.A2(n_739),
.B(n_735),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_734),
.B(n_465),
.C(n_492),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_743),
.A2(n_556),
.B(n_557),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_824),
.A2(n_540),
.B(n_547),
.C(n_670),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_779),
.B(n_823),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_745),
.A2(n_556),
.B(n_557),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_747),
.A2(n_547),
.B(n_616),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_751),
.A2(n_670),
.B(n_616),
.Y(n_927)
);

INVx4_ASAP7_75t_L g928 ( 
.A(n_763),
.Y(n_928)
);

AOI33xp33_ASAP7_75t_L g929 ( 
.A1(n_788),
.A2(n_465),
.A3(n_492),
.B1(n_496),
.B2(n_502),
.B3(n_447),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_759),
.Y(n_930)
);

NAND3xp33_ASAP7_75t_L g931 ( 
.A(n_714),
.B(n_670),
.C(n_616),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_775),
.A2(n_670),
.B(n_616),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_762),
.B(n_766),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_803),
.B(n_602),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_805),
.Y(n_935)
);

INVx2_ASAP7_75t_SL g936 ( 
.A(n_805),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_783),
.A2(n_616),
.B(n_583),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_776),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_795),
.B(n_583),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_796),
.B(n_583),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_802),
.B(n_583),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_838),
.A2(n_595),
.B(n_502),
.Y(n_942)
);

AO21x1_ASAP7_75t_L g943 ( 
.A1(n_785),
.A2(n_496),
.B(n_492),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_688),
.A2(n_579),
.B1(n_496),
.B2(n_502),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_804),
.A2(n_595),
.B(n_462),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_737),
.B(n_595),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_806),
.B(n_595),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_826),
.B(n_595),
.Y(n_948)
);

BUFx6f_ASAP7_75t_L g949 ( 
.A(n_737),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_800),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_798),
.A2(n_462),
.B(n_447),
.Y(n_951)
);

AOI22xp5_ASAP7_75t_L g952 ( 
.A1(n_721),
.A2(n_579),
.B1(n_233),
.B2(n_310),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_831),
.A2(n_595),
.B(n_462),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_744),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_810),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_744),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_832),
.B(n_447),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_721),
.A2(n_579),
.B1(n_228),
.B2(n_229),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_768),
.B(n_235),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_824),
.A2(n_462),
.B(n_487),
.C(n_475),
.Y(n_960)
);

AOI21xp33_ASAP7_75t_L g961 ( 
.A1(n_812),
.A2(n_278),
.B(n_243),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_828),
.A2(n_503),
.B(n_487),
.C(n_475),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_816),
.Y(n_963)
);

BUFx4f_ASAP7_75t_L g964 ( 
.A(n_744),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_840),
.A2(n_503),
.B(n_487),
.Y(n_965)
);

O2A1O1Ixp5_ASAP7_75t_L g966 ( 
.A1(n_731),
.A2(n_503),
.B(n_487),
.C(n_475),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_839),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_757),
.B(n_237),
.Y(n_968)
);

AOI21x1_ASAP7_75t_L g969 ( 
.A1(n_808),
.A2(n_451),
.B(n_450),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_731),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_820),
.A2(n_287),
.B(n_247),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_748),
.A2(n_291),
.B(n_252),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_810),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_757),
.B(n_246),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_757),
.B(n_253),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_757),
.B(n_254),
.Y(n_976)
);

AOI21xp33_ASAP7_75t_L g977 ( 
.A1(n_812),
.A2(n_294),
.B(n_259),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_830),
.B(n_257),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_698),
.A2(n_503),
.B1(n_487),
.B2(n_475),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_830),
.B(n_260),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_810),
.B(n_807),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_834),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_834),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_807),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_781),
.A2(n_503),
.B(n_487),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_734),
.B(n_261),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_834),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_738),
.B(n_263),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_738),
.B(n_451),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_834),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_715),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_828),
.B(n_266),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_774),
.A2(n_305),
.B(n_276),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_746),
.B(n_451),
.Y(n_994)
);

AOI21x1_ASAP7_75t_L g995 ( 
.A1(n_736),
.A2(n_451),
.B(n_450),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_722),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_781),
.A2(n_503),
.B(n_487),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_764),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_786),
.A2(n_503),
.B(n_487),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_756),
.A2(n_451),
.B(n_450),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_817),
.B(n_270),
.Y(n_1001)
);

NOR3xp33_ASAP7_75t_L g1002 ( 
.A(n_746),
.B(n_277),
.C(n_281),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_817),
.B(n_293),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_752),
.B(n_309),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_801),
.B(n_451),
.Y(n_1005)
);

NOR2xp67_ASAP7_75t_L g1006 ( 
.A(n_811),
.B(n_296),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_752),
.B(n_834),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_833),
.Y(n_1008)
);

CKINVDCx8_ASAP7_75t_R g1009 ( 
.A(n_814),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_698),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_748),
.A2(n_299),
.B(n_303),
.Y(n_1011)
);

BUFx8_ASAP7_75t_L g1012 ( 
.A(n_797),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_786),
.A2(n_787),
.B(n_789),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_787),
.A2(n_503),
.B(n_475),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_789),
.A2(n_475),
.B(n_451),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_749),
.B(n_15),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_835),
.A2(n_475),
.B(n_450),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_782),
.A2(n_450),
.B(n_449),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_750),
.B(n_18),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_750),
.A2(n_450),
.B(n_449),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_741),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_756),
.A2(n_782),
.B(n_784),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_742),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_780),
.A2(n_450),
.B(n_449),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_767),
.A2(n_450),
.B(n_449),
.Y(n_1025)
);

OAI21xp33_ASAP7_75t_L g1026 ( 
.A1(n_819),
.A2(n_449),
.B(n_446),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_767),
.B(n_19),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_861),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_888),
.B(n_722),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_1000),
.A2(n_784),
.B(n_760),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_841),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_858),
.A2(n_760),
.B(n_725),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_924),
.B(n_772),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_981),
.B(n_724),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_871),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_869),
.B(n_874),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_1009),
.B(n_825),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_885),
.Y(n_1038)
);

NAND2xp33_ASAP7_75t_SL g1039 ( 
.A(n_845),
.B(n_758),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_866),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_844),
.A2(n_998),
.B1(n_988),
.B2(n_986),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_862),
.B(n_791),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_930),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_981),
.B(n_449),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_906),
.B(n_676),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_935),
.B(n_21),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_964),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_846),
.A2(n_449),
.B(n_446),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_1004),
.B(n_22),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_1002),
.B(n_22),
.C(n_26),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_858),
.A2(n_449),
.B(n_446),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_849),
.A2(n_446),
.B(n_172),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_855),
.A2(n_159),
.B(n_151),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_877),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_847),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1055)
);

INVx3_ASAP7_75t_SL g1056 ( 
.A(n_950),
.Y(n_1056)
);

CKINVDCx8_ASAP7_75t_R g1057 ( 
.A(n_863),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_899),
.B(n_96),
.Y(n_1058)
);

AO221x2_ASAP7_75t_L g1059 ( 
.A1(n_1016),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.C(n_34),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_1007),
.B(n_30),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_964),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_880),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_978),
.A2(n_36),
.B(n_38),
.C(n_41),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_864),
.A2(n_134),
.B(n_122),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_936),
.B(n_41),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_853),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_842),
.B(n_45),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_933),
.A2(n_46),
.B1(n_48),
.B2(n_53),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_L g1069 ( 
.A1(n_943),
.A2(n_46),
.B(n_48),
.C(n_54),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_880),
.Y(n_1070)
);

OR2x6_ASAP7_75t_L g1071 ( 
.A(n_928),
.B(n_57),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_938),
.B(n_1008),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_860),
.A2(n_867),
.B(n_857),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_959),
.B(n_57),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_SL g1075 ( 
.A(n_1019),
.B(n_58),
.C(n_63),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_867),
.A2(n_58),
.B1(n_65),
.B2(n_76),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1001),
.B(n_80),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_856),
.A2(n_101),
.B(n_854),
.Y(n_1078)
);

INVx5_ASAP7_75t_L g1079 ( 
.A(n_955),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_980),
.A2(n_992),
.B(n_970),
.C(n_1027),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1003),
.B(n_984),
.Y(n_1081)
);

BUFx8_ASAP7_75t_L g1082 ( 
.A(n_949),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_866),
.B(n_865),
.Y(n_1083)
);

AO32x2_ASAP7_75t_L g1084 ( 
.A1(n_870),
.A2(n_875),
.A3(n_910),
.B1(n_916),
.B2(n_951),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_998),
.B(n_991),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_913),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_996),
.B(n_878),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_961),
.B(n_977),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_955),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_854),
.A2(n_852),
.B(n_851),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_973),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_852),
.A2(n_969),
.B(n_851),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_996),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_903),
.A2(n_859),
.B(n_883),
.C(n_886),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_920),
.A2(n_1013),
.B(n_900),
.C(n_1026),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_996),
.B(n_949),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_879),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_SL g1098 ( 
.A1(n_890),
.A2(n_993),
.B(n_894),
.C(n_1010),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_920),
.B(n_843),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_SL g1100 ( 
.A(n_972),
.B(n_1011),
.C(n_898),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_896),
.B(n_954),
.Y(n_1101)
);

NAND2x1p5_ASAP7_75t_L g1102 ( 
.A(n_973),
.B(n_863),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_917),
.A2(n_884),
.B(n_918),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_911),
.A2(n_915),
.B1(n_892),
.B2(n_872),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_954),
.B(n_956),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_908),
.B(n_1010),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_848),
.A2(n_887),
.B(n_873),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1006),
.B(n_934),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_949),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_L g1110 ( 
.A(n_1013),
.B(n_921),
.C(n_876),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_913),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_848),
.A2(n_881),
.B(n_882),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_897),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1005),
.B(n_913),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_963),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_962),
.A2(n_960),
.A3(n_923),
.B(n_1017),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_956),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_967),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_989),
.B(n_994),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_893),
.A2(n_901),
.B(n_895),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_1005),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_968),
.B(n_974),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1012),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1012),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1022),
.A2(n_931),
.B1(n_1023),
.B2(n_1021),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_907),
.B(n_929),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_957),
.Y(n_1127)
);

AND3x1_ASAP7_75t_SL g1128 ( 
.A(n_909),
.B(n_914),
.C(n_912),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_975),
.B(n_976),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_939),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_940),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_952),
.B(n_958),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_941),
.B(n_850),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_SL g1134 ( 
.A(n_971),
.B(n_904),
.C(n_889),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_919),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_946),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_893),
.A2(n_895),
.B(n_901),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_889),
.B(n_891),
.Y(n_1138)
);

OR2x6_ASAP7_75t_L g1139 ( 
.A(n_982),
.B(n_983),
.Y(n_1139)
);

NAND2x1_ASAP7_75t_L g1140 ( 
.A(n_987),
.B(n_990),
.Y(n_1140)
);

NAND2x1_ASAP7_75t_L g1141 ( 
.A(n_947),
.B(n_948),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_891),
.A2(n_902),
.B(n_904),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_868),
.B(n_1024),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_905),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_995),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_902),
.A2(n_937),
.B(n_932),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_927),
.A2(n_922),
.B(n_925),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_SL g1148 ( 
.A(n_1018),
.B(n_942),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_979),
.B(n_1025),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_965),
.B(n_945),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_922),
.B(n_925),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_945),
.A2(n_953),
.B1(n_1017),
.B2(n_999),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_966),
.A2(n_953),
.B(n_999),
.C(n_985),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_926),
.B(n_944),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_985),
.B(n_997),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_997),
.A2(n_1014),
.B1(n_1020),
.B2(n_1025),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1015),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_1020),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1015),
.Y(n_1159)
);

INVx4_ASAP7_75t_L g1160 ( 
.A(n_1014),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_869),
.B(n_733),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_844),
.B(n_526),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_924),
.B(n_709),
.Y(n_1163)
);

OAI21xp33_ASAP7_75t_L g1164 ( 
.A1(n_986),
.A2(n_563),
.B(n_988),
.Y(n_1164)
);

AOI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_874),
.A2(n_640),
.B1(n_644),
.B2(n_679),
.C(n_765),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_861),
.Y(n_1166)
);

AO22x1_ASAP7_75t_L g1167 ( 
.A1(n_986),
.A2(n_365),
.B1(n_367),
.B2(n_364),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_880),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_869),
.B(n_733),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_986),
.A2(n_728),
.B(n_1004),
.C(n_988),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_986),
.A2(n_728),
.B(n_1004),
.C(n_988),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_845),
.A2(n_846),
.B(n_849),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_888),
.B(n_733),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_871),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_924),
.B(n_709),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_845),
.A2(n_846),
.B(n_849),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_869),
.B(n_733),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_880),
.B(n_928),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_986),
.B(n_1004),
.C(n_988),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_924),
.B(n_709),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_888),
.B(n_733),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_861),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1179),
.A2(n_1164),
.B(n_1170),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1179),
.A2(n_1164),
.B(n_1171),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1051),
.A2(n_1092),
.B(n_1147),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1112),
.A2(n_1137),
.B(n_1120),
.Y(n_1186)
);

OAI21xp33_ASAP7_75t_L g1187 ( 
.A1(n_1049),
.A2(n_1074),
.B(n_1055),
.Y(n_1187)
);

AOI221x1_ASAP7_75t_L g1188 ( 
.A1(n_1076),
.A2(n_1088),
.B1(n_1078),
.B2(n_1066),
.C(n_1068),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1039),
.A2(n_1099),
.B(n_1076),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1031),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1028),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1038),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1056),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1073),
.A2(n_1176),
.B(n_1172),
.Y(n_1195)
);

AOI31xp67_ASAP7_75t_L g1196 ( 
.A1(n_1157),
.A2(n_1159),
.A3(n_1143),
.B(n_1138),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1146),
.A2(n_1142),
.B(n_1090),
.Y(n_1197)
);

AOI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1107),
.A2(n_1103),
.B(n_1155),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1180),
.B(n_1173),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1077),
.A2(n_1080),
.B(n_1037),
.C(n_1041),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1043),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1181),
.B(n_1162),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1095),
.A2(n_1156),
.A3(n_1152),
.B(n_1158),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1150),
.A2(n_1153),
.B(n_1030),
.Y(n_1205)
);

INVx8_ASAP7_75t_L g1206 ( 
.A(n_1079),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1148),
.A2(n_1149),
.B(n_1133),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1165),
.A2(n_1055),
.B1(n_1059),
.B2(n_1029),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1167),
.B(n_1081),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1040),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1148),
.A2(n_1094),
.B(n_1032),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1032),
.A2(n_1098),
.B(n_1104),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1104),
.A2(n_1141),
.B(n_1151),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1151),
.A2(n_1048),
.B(n_1052),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1126),
.A2(n_1060),
.B(n_1083),
.C(n_1132),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1145),
.A2(n_1064),
.B(n_1154),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1161),
.B(n_1169),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1177),
.B(n_1036),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1085),
.B(n_1046),
.Y(n_1219)
);

AOI221xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1068),
.A2(n_1063),
.B1(n_1045),
.B2(n_1130),
.C(n_1033),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1071),
.A2(n_1059),
.B1(n_1065),
.B2(n_1124),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1166),
.B(n_1182),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1108),
.B(n_1144),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1129),
.A2(n_1050),
.B(n_1122),
.C(n_1101),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1158),
.A2(n_1160),
.A3(n_1042),
.B(n_1106),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1082),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1071),
.A2(n_1087),
.B1(n_1034),
.B2(n_1123),
.Y(n_1227)
);

O2A1O1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1069),
.A2(n_1075),
.B(n_1110),
.C(n_1117),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1119),
.A2(n_1053),
.B(n_1110),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1140),
.A2(n_1160),
.B(n_1139),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1134),
.A2(n_1125),
.B(n_1100),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1086),
.B(n_1093),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1131),
.A2(n_1127),
.B(n_1105),
.Y(n_1233)
);

BUFx2_ASAP7_75t_R g1234 ( 
.A(n_1057),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1121),
.B(n_1047),
.Y(n_1235)
);

A2O1A1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1034),
.A2(n_1135),
.B(n_1096),
.C(n_1114),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1111),
.B(n_1082),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1044),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1079),
.Y(n_1239)
);

AOI221x1_ASAP7_75t_L g1240 ( 
.A1(n_1115),
.A2(n_1118),
.B1(n_1136),
.B2(n_1111),
.C(n_1121),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1035),
.A2(n_1174),
.B1(n_1097),
.B2(n_1054),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1044),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1136),
.A2(n_1047),
.B(n_1061),
.C(n_1089),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1084),
.A2(n_1116),
.A3(n_1128),
.B(n_1139),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1109),
.Y(n_1245)
);

AOI31xp67_ASAP7_75t_L g1246 ( 
.A1(n_1084),
.A2(n_1116),
.A3(n_1136),
.B(n_1109),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_1109),
.B(n_1178),
.Y(n_1247)
);

BUFx10_ASAP7_75t_L g1248 ( 
.A(n_1089),
.Y(n_1248)
);

INVx6_ASAP7_75t_L g1249 ( 
.A(n_1079),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1089),
.A2(n_1091),
.B(n_1168),
.C(n_1058),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1091),
.A2(n_1168),
.B(n_1116),
.C(n_1178),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1062),
.A2(n_1070),
.B(n_1168),
.C(n_1091),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1070),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1164),
.A2(n_1179),
.B(n_1049),
.C(n_1088),
.Y(n_1254)
);

AOI221x1_ASAP7_75t_L g1255 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1170),
.B2(n_1171),
.C(n_1049),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1256)
);

NOR4xp25_ASAP7_75t_L g1257 ( 
.A(n_1164),
.B(n_1179),
.C(n_1171),
.D(n_1170),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1178),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1095),
.A2(n_943),
.A3(n_951),
.B(n_1156),
.Y(n_1259)
);

AOI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1051),
.A2(n_1143),
.B(n_1147),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1164),
.A2(n_1179),
.B(n_1049),
.C(n_1088),
.Y(n_1261)
);

CKINVDCx20_ASAP7_75t_R g1262 ( 
.A(n_1031),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_1031),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_R g1264 ( 
.A(n_1031),
.B(n_727),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1171),
.B2(n_1170),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1028),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1162),
.B(n_844),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_1179),
.B(n_1079),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1113),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1051),
.A2(n_1092),
.B(n_1147),
.Y(n_1271)
);

OAI221xp5_ASAP7_75t_L g1272 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1049),
.B2(n_1074),
.C(n_1171),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1047),
.Y(n_1273)
);

BUFx12f_ASAP7_75t_L g1274 ( 
.A(n_1124),
.Y(n_1274)
);

INVxp67_ASAP7_75t_SL g1275 ( 
.A(n_1106),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1031),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1164),
.B(n_1179),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1164),
.A2(n_718),
.B1(n_369),
.B2(n_366),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1028),
.Y(n_1280)
);

INVx8_ASAP7_75t_L g1281 ( 
.A(n_1079),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1031),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1179),
.A2(n_1164),
.B(n_1170),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1074),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1120),
.A2(n_1137),
.B(n_1142),
.Y(n_1285)
);

INVx1_ASAP7_75t_SL g1286 ( 
.A(n_1093),
.Y(n_1286)
);

AOI21xp33_ASAP7_75t_L g1287 ( 
.A1(n_1164),
.A2(n_1179),
.B(n_1088),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1179),
.A2(n_1055),
.B1(n_1037),
.B2(n_1009),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1164),
.A2(n_1179),
.B1(n_1171),
.B2(n_1170),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1028),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1173),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1164),
.A2(n_1179),
.B(n_1049),
.C(n_1088),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1095),
.A2(n_943),
.A3(n_951),
.B(n_1156),
.Y(n_1294)
);

OA21x2_ASAP7_75t_L g1295 ( 
.A1(n_1120),
.A2(n_1137),
.B(n_1142),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1047),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1164),
.B(n_577),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1051),
.A2(n_1092),
.B(n_1147),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1102),
.B(n_880),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1047),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1164),
.A2(n_1179),
.B(n_1049),
.C(n_1088),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1028),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1028),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1028),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1051),
.A2(n_1092),
.B(n_1147),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1028),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1309)
);

INVx1_ASAP7_75t_SL g1310 ( 
.A(n_1093),
.Y(n_1310)
);

OA21x2_ASAP7_75t_L g1311 ( 
.A1(n_1120),
.A2(n_1137),
.B(n_1142),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1028),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1028),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1031),
.Y(n_1314)
);

NAND2x1p5_ASAP7_75t_L g1315 ( 
.A(n_1079),
.B(n_880),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_1162),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1163),
.B(n_1175),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.C(n_1179),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1164),
.A2(n_1179),
.B(n_1049),
.C(n_1088),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1056),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1047),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1170),
.A2(n_1171),
.B(n_1164),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1028),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1028),
.Y(n_1327)
);

CKINVDCx6p67_ASAP7_75t_R g1328 ( 
.A(n_1056),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1164),
.B(n_577),
.Y(n_1329)
);

BUFx2_ASAP7_75t_R g1330 ( 
.A(n_1194),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1187),
.A2(n_1221),
.B1(n_1208),
.B2(n_1288),
.Y(n_1331)
);

INVx4_ASAP7_75t_L g1332 ( 
.A(n_1191),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1187),
.A2(n_1221),
.B1(n_1208),
.B2(n_1272),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1279),
.A2(n_1329),
.B1(n_1298),
.B2(n_1287),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1192),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1262),
.Y(n_1336)
);

INVx4_ASAP7_75t_SL g1337 ( 
.A(n_1249),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1254),
.A2(n_1261),
.B1(n_1321),
.B2(n_1303),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_SL g1339 ( 
.A1(n_1265),
.A2(n_1290),
.B1(n_1184),
.B2(n_1183),
.Y(n_1339)
);

INVx3_ASAP7_75t_SL g1340 ( 
.A(n_1328),
.Y(n_1340)
);

INVx2_ASAP7_75t_SL g1341 ( 
.A(n_1264),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1276),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1263),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1322),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1283),
.A2(n_1284),
.B1(n_1209),
.B2(n_1316),
.Y(n_1345)
);

BUFx2_ASAP7_75t_SL g1346 ( 
.A(n_1282),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1274),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1284),
.A2(n_1269),
.B1(n_1319),
.B2(n_1324),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1267),
.A2(n_1277),
.B1(n_1219),
.B2(n_1223),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1275),
.B(n_1257),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1210),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1300),
.A2(n_1309),
.B1(n_1325),
.B2(n_1270),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1292),
.B(n_1317),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1202),
.B(n_1199),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1211),
.A2(n_1203),
.B1(n_1231),
.B2(n_1212),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1193),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1293),
.A2(n_1200),
.B1(n_1256),
.B2(n_1278),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1201),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1314),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1226),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1255),
.A2(n_1188),
.B(n_1227),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1218),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1266),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1190),
.A2(n_1318),
.B1(n_1289),
.B2(n_1297),
.Y(n_1364)
);

BUFx4f_ASAP7_75t_SL g1365 ( 
.A(n_1286),
.Y(n_1365)
);

BUFx8_ASAP7_75t_L g1366 ( 
.A(n_1273),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1280),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1320),
.A2(n_1195),
.B(n_1213),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1248),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1291),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1217),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1189),
.A2(n_1241),
.B1(n_1238),
.B2(n_1242),
.Y(n_1372)
);

INVx4_ASAP7_75t_L g1373 ( 
.A(n_1206),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1304),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1305),
.Y(n_1375)
);

BUFx6f_ASAP7_75t_L g1376 ( 
.A(n_1206),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1257),
.A2(n_1308),
.B1(n_1306),
.B2(n_1312),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1227),
.A2(n_1313),
.B1(n_1327),
.B2(n_1326),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1224),
.A2(n_1207),
.B1(n_1228),
.B2(n_1268),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1233),
.Y(n_1380)
);

INVx5_ASAP7_75t_L g1381 ( 
.A(n_1281),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1232),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1268),
.A2(n_1229),
.B1(n_1253),
.B2(n_1247),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1245),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1196),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1244),
.B(n_1220),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1286),
.B(n_1310),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1237),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1310),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1236),
.A2(n_1250),
.B1(n_1251),
.B2(n_1258),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1273),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1246),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1234),
.Y(n_1393)
);

AOI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1220),
.A2(n_1235),
.B1(n_1215),
.B2(n_1301),
.Y(n_1394)
);

INVx6_ASAP7_75t_L g1395 ( 
.A(n_1248),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1240),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1244),
.A2(n_1323),
.B1(n_1302),
.B2(n_1296),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1302),
.A2(n_1323),
.B1(n_1301),
.B2(n_1216),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1225),
.Y(n_1399)
);

BUFx3_ASAP7_75t_L g1400 ( 
.A(n_1315),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1239),
.Y(n_1401)
);

BUFx2_ASAP7_75t_L g1402 ( 
.A(n_1239),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1205),
.A2(n_1230),
.B(n_1214),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1243),
.A2(n_1198),
.B1(n_1285),
.B2(n_1295),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1204),
.B(n_1259),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1285),
.A2(n_1311),
.B1(n_1295),
.B2(n_1204),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1252),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1260),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1185),
.A2(n_1271),
.B1(n_1299),
.B2(n_1307),
.Y(n_1409)
);

CKINVDCx20_ASAP7_75t_R g1410 ( 
.A(n_1259),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1197),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1186),
.A2(n_1187),
.B1(n_1164),
.B2(n_1221),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1294),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1221),
.B2(n_1208),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1221),
.B2(n_1208),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1221),
.B2(n_1208),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1208),
.A2(n_1179),
.B1(n_1187),
.B2(n_1164),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1222),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1206),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1222),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1221),
.B2(n_1208),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1206),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1221),
.B2(n_1208),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1037),
.B2(n_1288),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_1322),
.Y(n_1425)
);

INVx8_ASAP7_75t_L g1426 ( 
.A(n_1206),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1221),
.B2(n_1208),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1322),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1037),
.B2(n_1288),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1208),
.A2(n_1179),
.B1(n_1272),
.B2(n_1288),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1222),
.Y(n_1431)
);

CKINVDCx6p67_ASAP7_75t_R g1432 ( 
.A(n_1322),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1276),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1187),
.A2(n_1164),
.B1(n_1037),
.B2(n_1288),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1194),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1322),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1322),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1222),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1286),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1322),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1275),
.B(n_1257),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1276),
.Y(n_1442)
);

CKINVDCx14_ASAP7_75t_R g1443 ( 
.A(n_1264),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_SL g1444 ( 
.A1(n_1208),
.A2(n_1272),
.B1(n_1209),
.B2(n_1049),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1386),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1368),
.A2(n_1403),
.B(n_1404),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1386),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1350),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1392),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1364),
.B(n_1339),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1403),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1335),
.B(n_1363),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1368),
.A2(n_1404),
.B(n_1409),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1408),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1385),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1424),
.A2(n_1434),
.B(n_1429),
.Y(n_1456)
);

INVx1_ASAP7_75t_SL g1457 ( 
.A(n_1389),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1367),
.B(n_1370),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1350),
.Y(n_1459)
);

AO21x2_ASAP7_75t_L g1460 ( 
.A1(n_1405),
.A2(n_1441),
.B(n_1399),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1441),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1374),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1375),
.B(n_1339),
.Y(n_1463)
);

OR2x2_ASAP7_75t_L g1464 ( 
.A(n_1405),
.B(n_1413),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1354),
.B(n_1357),
.Y(n_1465)
);

NOR2x1_ASAP7_75t_SL g1466 ( 
.A(n_1379),
.B(n_1390),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1387),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1411),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1356),
.B(n_1358),
.Y(n_1469)
);

AND2x6_ASAP7_75t_L g1470 ( 
.A(n_1394),
.B(n_1380),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1407),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1411),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1355),
.B(n_1348),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1383),
.A2(n_1352),
.B(n_1379),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1410),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1383),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1396),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1373),
.Y(n_1478)
);

BUFx2_ASAP7_75t_R g1479 ( 
.A(n_1393),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1417),
.A2(n_1338),
.B(n_1430),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1361),
.B(n_1390),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1412),
.A2(n_1338),
.B(n_1372),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1384),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1402),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1389),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1355),
.B(n_1348),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1381),
.Y(n_1487)
);

BUFx4f_ASAP7_75t_SL g1488 ( 
.A(n_1425),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1342),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1357),
.B(n_1418),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1377),
.B(n_1345),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1420),
.Y(n_1492)
);

OAI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1417),
.A2(n_1444),
.B(n_1333),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1439),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1407),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1433),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1414),
.A2(n_1416),
.B1(n_1423),
.B2(n_1427),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1439),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1337),
.B(n_1376),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1377),
.B(n_1345),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1382),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1431),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1442),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1371),
.A2(n_1362),
.B1(n_1331),
.B2(n_1378),
.Y(n_1504)
);

OR2x2_ASAP7_75t_L g1505 ( 
.A(n_1438),
.B(n_1415),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1397),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1443),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1397),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1407),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1353),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1406),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1406),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1421),
.B(n_1349),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1359),
.B(n_1334),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1378),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1398),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1398),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1401),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1391),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1426),
.A2(n_1419),
.B(n_1422),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1388),
.A2(n_1435),
.B(n_1343),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1346),
.B(n_1422),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1497),
.A2(n_1360),
.B1(n_1365),
.B2(n_1341),
.Y(n_1523)
);

AO21x2_ASAP7_75t_L g1524 ( 
.A1(n_1477),
.A2(n_1456),
.B(n_1480),
.Y(n_1524)
);

OAI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1480),
.A2(n_1332),
.B(n_1400),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1448),
.B(n_1366),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1467),
.B(n_1336),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1497),
.A2(n_1351),
.B1(n_1347),
.B2(n_1366),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1488),
.Y(n_1529)
);

OAI211xp5_ASAP7_75t_L g1530 ( 
.A1(n_1493),
.A2(n_1437),
.B(n_1344),
.C(n_1332),
.Y(n_1530)
);

AND2x4_ASAP7_75t_SL g1531 ( 
.A(n_1499),
.B(n_1432),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1456),
.A2(n_1493),
.B(n_1450),
.C(n_1491),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1467),
.B(n_1340),
.Y(n_1533)
);

BUFx12f_ASAP7_75t_L g1534 ( 
.A(n_1507),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1510),
.B(n_1340),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1448),
.B(n_1395),
.Y(n_1536)
);

OR2x6_ASAP7_75t_L g1537 ( 
.A(n_1481),
.B(n_1426),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1504),
.A2(n_1428),
.B1(n_1369),
.B2(n_1436),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1450),
.A2(n_1440),
.B1(n_1330),
.B2(n_1395),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1503),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1501),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1503),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_L g1543 ( 
.A1(n_1473),
.A2(n_1330),
.B1(n_1395),
.B2(n_1426),
.C(n_1486),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1473),
.A2(n_1486),
.B(n_1474),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1457),
.B(n_1485),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1466),
.A2(n_1476),
.B(n_1446),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1494),
.B(n_1498),
.Y(n_1547)
);

NOR2xp67_ASAP7_75t_L g1548 ( 
.A(n_1471),
.B(n_1459),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1481),
.A2(n_1465),
.B1(n_1491),
.B2(n_1500),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1462),
.B(n_1521),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1459),
.B(n_1461),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1521),
.B(n_1484),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1500),
.A2(n_1476),
.B(n_1482),
.C(n_1474),
.Y(n_1553)
);

OAI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1481),
.A2(n_1513),
.B1(n_1490),
.B2(n_1505),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1521),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1462),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1452),
.B(n_1458),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1483),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1452),
.B(n_1458),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1466),
.A2(n_1446),
.B(n_1451),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1478),
.Y(n_1561)
);

A2O1A1Ixp33_ASAP7_75t_L g1562 ( 
.A1(n_1482),
.A2(n_1513),
.B(n_1463),
.C(n_1515),
.Y(n_1562)
);

OAI21xp5_ASAP7_75t_L g1563 ( 
.A1(n_1481),
.A2(n_1515),
.B(n_1470),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1489),
.B(n_1496),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1495),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1505),
.A2(n_1463),
.B1(n_1514),
.B2(n_1495),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1522),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1518),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1483),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1477),
.A2(n_1512),
.B(n_1511),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1461),
.B(n_1445),
.Y(n_1571)
);

NAND2x1_ASAP7_75t_L g1572 ( 
.A(n_1470),
.B(n_1487),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1509),
.A2(n_1451),
.B1(n_1517),
.B2(n_1516),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1519),
.B(n_1522),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1449),
.B(n_1445),
.C(n_1447),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1447),
.B(n_1492),
.Y(n_1577)
);

CKINVDCx10_ASAP7_75t_R g1578 ( 
.A(n_1479),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1516),
.A2(n_1517),
.B(n_1506),
.C(n_1508),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1550),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1552),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1556),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1549),
.A2(n_1470),
.B1(n_1508),
.B2(n_1506),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1449),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1558),
.Y(n_1587)
);

NAND2x1p5_ASAP7_75t_L g1588 ( 
.A(n_1572),
.B(n_1453),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1569),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1544),
.B(n_1472),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1577),
.Y(n_1591)
);

BUFx2_ASAP7_75t_SL g1592 ( 
.A(n_1548),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1549),
.A2(n_1470),
.B1(n_1475),
.B2(n_1464),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1554),
.A2(n_1470),
.B1(n_1475),
.B2(n_1464),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1555),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1560),
.B(n_1468),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1524),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1560),
.B(n_1468),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1571),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1547),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1546),
.B(n_1455),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1576),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1537),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1554),
.A2(n_1470),
.B1(n_1475),
.B2(n_1492),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1536),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1541),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1524),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1545),
.B(n_1454),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1553),
.B(n_1540),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1575),
.B(n_1454),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1553),
.B(n_1502),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1608),
.A2(n_1562),
.B(n_1532),
.Y(n_1613)
);

OAI211xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1603),
.A2(n_1530),
.B(n_1532),
.C(n_1523),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1584),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1583),
.B(n_1581),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1594),
.B(n_1563),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1594),
.B(n_1565),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_R g1619 ( 
.A(n_1604),
.B(n_1578),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1603),
.B(n_1530),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1597),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1584),
.Y(n_1622)
);

OAI31xp33_ASAP7_75t_L g1623 ( 
.A1(n_1585),
.A2(n_1562),
.A3(n_1539),
.B(n_1580),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1574),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1581),
.B(n_1568),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1587),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1579),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_SL g1628 ( 
.A1(n_1585),
.A2(n_1539),
.B1(n_1537),
.B2(n_1538),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1596),
.Y(n_1629)
);

AOI33xp33_ASAP7_75t_L g1630 ( 
.A1(n_1596),
.A2(n_1542),
.A3(n_1564),
.B1(n_1528),
.B2(n_1543),
.B3(n_1535),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1602),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1597),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1610),
.Y(n_1633)
);

AND2x2_ASAP7_75t_SL g1634 ( 
.A(n_1593),
.B(n_1543),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1582),
.B(n_1566),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1607),
.B(n_1533),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1588),
.Y(n_1637)
);

NOR3xp33_ASAP7_75t_L g1638 ( 
.A(n_1610),
.B(n_1526),
.C(n_1525),
.Y(n_1638)
);

OAI31xp33_ASAP7_75t_L g1639 ( 
.A1(n_1605),
.A2(n_1580),
.A3(n_1566),
.B(n_1573),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1586),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1527),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1599),
.B(n_1570),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1600),
.B(n_1460),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1589),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1640),
.B(n_1586),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1629),
.B(n_1642),
.Y(n_1647)
);

NAND2x1_ASAP7_75t_SL g1648 ( 
.A(n_1643),
.B(n_1590),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1640),
.B(n_1600),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1645),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1632),
.B(n_1591),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1622),
.Y(n_1655)
);

NOR4xp25_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1630),
.C(n_1620),
.D(n_1633),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1632),
.B(n_1591),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1619),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_SL g1660 ( 
.A(n_1620),
.B(n_1590),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1616),
.B(n_1609),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1642),
.B(n_1595),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1619),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1635),
.B(n_1586),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1622),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1616),
.B(n_1609),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1616),
.B(n_1609),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1631),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1642),
.B(n_1595),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1631),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1627),
.B(n_1592),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1626),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1627),
.B(n_1592),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1635),
.B(n_1606),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1627),
.B(n_1592),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1614),
.B(n_1526),
.C(n_1525),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1636),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1624),
.B(n_1611),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1626),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1636),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1630),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1650),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1680),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_L g1686 ( 
.A(n_1663),
.B(n_1617),
.Y(n_1686)
);

OAI32xp33_ASAP7_75t_L g1687 ( 
.A1(n_1656),
.A2(n_1638),
.A3(n_1618),
.B1(n_1617),
.B2(n_1643),
.Y(n_1687)
);

INVx2_ASAP7_75t_SL g1688 ( 
.A(n_1659),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1651),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1648),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1648),
.Y(n_1691)
);

INVxp67_ASAP7_75t_SL g1692 ( 
.A(n_1659),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1669),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1647),
.B(n_1642),
.Y(n_1694)
);

INVx2_ASAP7_75t_SL g1695 ( 
.A(n_1663),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1651),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1652),
.B(n_1624),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1654),
.Y(n_1698)
);

NAND2x1_ASAP7_75t_L g1699 ( 
.A(n_1647),
.B(n_1625),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1678),
.B(n_1534),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1654),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1664),
.B(n_1644),
.Y(n_1702)
);

NAND3xp33_ASAP7_75t_SL g1703 ( 
.A(n_1677),
.B(n_1623),
.C(n_1639),
.Y(n_1703)
);

NAND2x1p5_ASAP7_75t_SL g1704 ( 
.A(n_1660),
.B(n_1618),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1669),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1681),
.Y(n_1706)
);

INVxp33_ASAP7_75t_L g1707 ( 
.A(n_1652),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1655),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1658),
.B(n_1624),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1682),
.B(n_1638),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1681),
.B(n_1529),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1658),
.B(n_1679),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1669),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1664),
.B(n_1644),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1679),
.B(n_1641),
.Y(n_1715)
);

INVxp67_ASAP7_75t_SL g1716 ( 
.A(n_1647),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1668),
.B(n_1567),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1655),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1647),
.B(n_1637),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1665),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1641),
.Y(n_1721)
);

BUFx12f_ASAP7_75t_L g1722 ( 
.A(n_1662),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1671),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1671),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1665),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1697),
.B(n_1709),
.Y(n_1726)
);

OAI31xp33_ASAP7_75t_L g1727 ( 
.A1(n_1683),
.A2(n_1623),
.A3(n_1639),
.B(n_1628),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1697),
.B(n_1672),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1709),
.B(n_1672),
.Y(n_1729)
);

CKINVDCx16_ASAP7_75t_R g1730 ( 
.A(n_1703),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1712),
.B(n_1674),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1712),
.B(n_1674),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1687),
.B(n_1675),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1689),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1689),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1696),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1695),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1695),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1692),
.Y(n_1739)
);

AND2x4_ASAP7_75t_SL g1740 ( 
.A(n_1694),
.B(n_1662),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1696),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1687),
.B(n_1675),
.Y(n_1742)
);

AOI21xp5_ASAP7_75t_L g1743 ( 
.A1(n_1686),
.A2(n_1628),
.B(n_1634),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1686),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1710),
.B(n_1661),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1686),
.B(n_1661),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1698),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1704),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1715),
.B(n_1676),
.Y(n_1749)
);

INVxp67_ASAP7_75t_SL g1750 ( 
.A(n_1688),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1722),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1698),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1716),
.B(n_1662),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1699),
.B(n_1662),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1715),
.B(n_1676),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1704),
.B(n_1646),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1688),
.B(n_1646),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1706),
.B(n_1649),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1759)
);

NAND4xp25_ASAP7_75t_L g1760 ( 
.A(n_1711),
.B(n_1670),
.C(n_1605),
.D(n_1593),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1684),
.B(n_1649),
.Y(n_1761)
);

OAI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1748),
.A2(n_1690),
.B1(n_1691),
.B2(n_1707),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1734),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1739),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1756),
.B(n_1745),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1726),
.B(n_1694),
.Y(n_1766)
);

NOR4xp25_ASAP7_75t_L g1767 ( 
.A(n_1748),
.B(n_1684),
.C(n_1685),
.D(n_1691),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1748),
.A2(n_1634),
.B(n_1690),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1739),
.B(n_1721),
.Y(n_1769)
);

NOR2xp67_ASAP7_75t_SL g1770 ( 
.A(n_1730),
.B(n_1722),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1740),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1734),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1737),
.B(n_1685),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1756),
.B(n_1702),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1717),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1738),
.B(n_1666),
.Y(n_1776)
);

NAND2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1746),
.B(n_1699),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1730),
.A2(n_1634),
.B1(n_1613),
.B2(n_1643),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1733),
.B(n_1700),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1727),
.B(n_1667),
.Y(n_1780)
);

AOI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1727),
.A2(n_1634),
.B1(n_1613),
.B2(n_1608),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1735),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1733),
.B(n_1702),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1753),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1735),
.Y(n_1786)
);

OAI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1742),
.A2(n_1612),
.B1(n_1537),
.B2(n_1573),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1763),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1772),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1750),
.Y(n_1790)
);

OAI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1778),
.A2(n_1743),
.B1(n_1744),
.B2(n_1760),
.C(n_1751),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1782),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1786),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1773),
.Y(n_1794)
);

AOI21xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1767),
.A2(n_1762),
.B(n_1780),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1781),
.A2(n_1744),
.B(n_1757),
.Y(n_1796)
);

AOI21xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1762),
.A2(n_1751),
.B(n_1753),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1781),
.A2(n_1744),
.B1(n_1613),
.B2(n_1760),
.Y(n_1798)
);

OAI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1768),
.A2(n_1758),
.B1(n_1761),
.B2(n_1741),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1774),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1766),
.B(n_1726),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1783),
.A2(n_1758),
.B1(n_1761),
.B2(n_1754),
.C(n_1723),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1787),
.B(n_1754),
.Y(n_1803)
);

NAND2x1p5_ASAP7_75t_L g1804 ( 
.A(n_1770),
.B(n_1753),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1769),
.B(n_1731),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1779),
.B(n_1753),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1765),
.B(n_1731),
.Y(n_1807)
);

OAI31xp33_ASAP7_75t_L g1808 ( 
.A1(n_1791),
.A2(n_1785),
.A3(n_1787),
.B(n_1779),
.Y(n_1808)
);

XNOR2x1_ASAP7_75t_L g1809 ( 
.A(n_1804),
.B(n_1775),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1795),
.B(n_1736),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1800),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1801),
.B(n_1784),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1790),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1788),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1799),
.A2(n_1777),
.B1(n_1736),
.B2(n_1752),
.C(n_1741),
.Y(n_1815)
);

OAI21xp33_ASAP7_75t_L g1816 ( 
.A1(n_1803),
.A2(n_1771),
.B(n_1776),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1804),
.B(n_1740),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1789),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1792),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_L g1820 ( 
.A(n_1810),
.B(n_1806),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1812),
.B(n_1807),
.Y(n_1821)
);

NOR4xp75_ASAP7_75t_SL g1822 ( 
.A(n_1810),
.B(n_1805),
.C(n_1797),
.D(n_1806),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1809),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1811),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1813),
.B(n_1799),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1814),
.B(n_1794),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1818),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1819),
.B(n_1816),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1817),
.B(n_1793),
.Y(n_1829)
);

AOI221xp5_ASAP7_75t_L g1830 ( 
.A1(n_1825),
.A2(n_1798),
.B1(n_1796),
.B2(n_1802),
.C(n_1808),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1823),
.A2(n_1798),
.B1(n_1815),
.B2(n_1828),
.C(n_1824),
.Y(n_1831)
);

NAND4xp25_ASAP7_75t_L g1832 ( 
.A(n_1820),
.B(n_1821),
.C(n_1829),
.D(n_1826),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1827),
.A2(n_1613),
.B1(n_1693),
.B2(n_1705),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1822),
.A2(n_1740),
.B1(n_1719),
.B2(n_1752),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1830),
.A2(n_1747),
.B1(n_1732),
.B2(n_1729),
.Y(n_1835)
);

NAND3xp33_ASAP7_75t_SL g1836 ( 
.A(n_1831),
.B(n_1747),
.C(n_1732),
.Y(n_1836)
);

AOI31xp33_ASAP7_75t_L g1837 ( 
.A1(n_1834),
.A2(n_1759),
.A3(n_1729),
.B(n_1728),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1832),
.B(n_1759),
.Y(n_1838)
);

OAI321xp33_ASAP7_75t_L g1839 ( 
.A1(n_1833),
.A2(n_1714),
.A3(n_1728),
.B1(n_1713),
.B2(n_1693),
.C(n_1723),
.Y(n_1839)
);

NOR2xp67_ASAP7_75t_L g1840 ( 
.A(n_1832),
.B(n_1749),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1838),
.Y(n_1841)
);

XNOR2xp5_ASAP7_75t_L g1842 ( 
.A(n_1835),
.B(n_1531),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_L g1843 ( 
.A(n_1836),
.B(n_1840),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1837),
.B(n_1749),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1839),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_L g1846 ( 
.A(n_1843),
.B(n_1719),
.C(n_1713),
.Y(n_1846)
);

NOR3xp33_ASAP7_75t_SL g1847 ( 
.A(n_1844),
.B(n_1708),
.C(n_1701),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1841),
.B(n_1755),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1849),
.Y(n_1850)
);

INVxp67_ASAP7_75t_SL g1851 ( 
.A(n_1850),
.Y(n_1851)
);

INVx3_ASAP7_75t_SL g1852 ( 
.A(n_1850),
.Y(n_1852)
);

OAI22x1_ASAP7_75t_L g1853 ( 
.A1(n_1852),
.A2(n_1842),
.B1(n_1846),
.B2(n_1845),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1851),
.A2(n_1847),
.B1(n_1755),
.B2(n_1705),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1853),
.A2(n_1725),
.B1(n_1701),
.B2(n_1720),
.Y(n_1855)
);

OAI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1854),
.A2(n_1724),
.B(n_1718),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1855),
.B(n_1856),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1857),
.A2(n_1724),
.B1(n_1725),
.B2(n_1720),
.C(n_1718),
.Y(n_1858)
);

AOI22x1_ASAP7_75t_L g1859 ( 
.A1(n_1858),
.A2(n_1708),
.B1(n_1670),
.B2(n_1673),
.Y(n_1859)
);

AOI221xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1653),
.B1(n_1657),
.B2(n_1621),
.C(n_1671),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1657),
.B(n_1653),
.C(n_1520),
.Y(n_1861)
);


endmodule