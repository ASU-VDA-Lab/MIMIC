module real_aes_6495_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_666;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_175;
wire n_168;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g542 ( .A1(n_0), .A2(n_190), .B(n_543), .C(n_546), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_1), .B(n_531), .Y(n_547) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_3), .A2(n_752), .B1(n_755), .B2(n_756), .Y(n_751) );
INVx1_ASAP7_75t_L g756 ( .A(n_3), .Y(n_756) );
INVx1_ASAP7_75t_L g208 ( .A(n_4), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_5), .B(n_179), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_6), .A2(n_446), .B(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_7), .A2(n_103), .B1(n_117), .B2(n_763), .Y(n_102) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_8), .A2(n_155), .B(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_9), .A2(n_37), .B1(n_135), .B2(n_144), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_10), .B(n_155), .Y(n_219) );
AND2x6_ASAP7_75t_L g153 ( .A(n_11), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g505 ( .A1(n_12), .A2(n_153), .B(n_449), .C(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g109 ( .A(n_13), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_13), .B(n_38), .Y(n_435) );
INVx1_ASAP7_75t_L g151 ( .A(n_14), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_15), .B(n_142), .Y(n_162) );
INVx1_ASAP7_75t_L g200 ( .A(n_16), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_17), .B(n_179), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_18), .B(n_156), .Y(n_224) );
AO32x2_ASAP7_75t_L g187 ( .A1(n_19), .A2(n_152), .A3(n_155), .B1(n_188), .B2(n_192), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_20), .B(n_144), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_21), .B(n_156), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_22), .A2(n_53), .B1(n_135), .B2(n_144), .Y(n_191) );
AOI22xp33_ASAP7_75t_SL g141 ( .A1(n_23), .A2(n_82), .B1(n_142), .B2(n_144), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_24), .B(n_144), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_25), .A2(n_152), .B(n_449), .C(n_451), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_26), .A2(n_152), .B(n_449), .C(n_496), .Y(n_495) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_28), .B(n_147), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_29), .A2(n_446), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_30), .B(n_147), .Y(n_185) );
INVx2_ASAP7_75t_L g137 ( .A(n_31), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_32), .A2(n_470), .B(n_479), .C(n_481), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_33), .B(n_144), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_34), .B(n_147), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g119 ( .A1(n_35), .A2(n_74), .B1(n_120), .B2(n_121), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_35), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_36), .B(n_164), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_38), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_39), .B(n_445), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_40), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_41), .B(n_179), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_42), .B(n_446), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_43), .A2(n_470), .B(n_479), .C(n_516), .Y(n_515) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_44), .A2(n_125), .B1(n_429), .B2(n_430), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_44), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_44), .A2(n_80), .B1(n_429), .B2(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_45), .B(n_144), .Y(n_214) );
INVx1_ASAP7_75t_L g544 ( .A(n_46), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_47), .A2(n_90), .B1(n_135), .B2(n_138), .Y(n_134) );
INVx1_ASAP7_75t_L g517 ( .A(n_48), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_49), .B(n_144), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_50), .B(n_144), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_51), .B(n_446), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_52), .B(n_206), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g228 ( .A1(n_54), .A2(n_59), .B1(n_142), .B2(n_144), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_55), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_56), .B(n_144), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_57), .B(n_144), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_58), .Y(n_760) );
INVx1_ASAP7_75t_L g154 ( .A(n_60), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_61), .B(n_446), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_62), .B(n_531), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_63), .A2(n_203), .B(n_206), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_64), .B(n_144), .Y(n_209) );
INVx1_ASAP7_75t_L g150 ( .A(n_65), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_66), .Y(n_747) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_67), .B(n_179), .Y(n_483) );
AO32x2_ASAP7_75t_L g132 ( .A1(n_68), .A2(n_133), .A3(n_146), .B1(n_152), .B2(n_155), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_69), .B(n_145), .Y(n_507) );
INVx1_ASAP7_75t_L g242 ( .A(n_70), .Y(n_242) );
INVx1_ASAP7_75t_L g177 ( .A(n_71), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_72), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_73), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g121 ( .A(n_74), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_75), .A2(n_449), .B(n_466), .C(n_470), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_76), .B(n_142), .Y(n_178) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_77), .Y(n_526) );
INVx1_ASAP7_75t_L g116 ( .A(n_78), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_79), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_80), .Y(n_754) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_81), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_83), .B(n_135), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_84), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_85), .B(n_142), .Y(n_182) );
INVx2_ASAP7_75t_L g148 ( .A(n_86), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_87), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_88), .B(n_139), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_89), .B(n_142), .Y(n_215) );
INVx2_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
OR2x2_ASAP7_75t_L g433 ( .A(n_91), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g750 ( .A(n_91), .B(n_744), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_92), .A2(n_101), .B1(n_142), .B2(n_143), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_93), .B(n_446), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_94), .Y(n_482) );
INVxp67_ASAP7_75t_L g529 ( .A(n_95), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_96), .B(n_142), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_97), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g467 ( .A(n_98), .Y(n_467) );
INVx1_ASAP7_75t_L g503 ( .A(n_99), .Y(n_503) );
AND2x2_ASAP7_75t_L g519 ( .A(n_100), .B(n_147), .Y(n_519) );
BUFx4f_ASAP7_75t_SL g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g765 ( .A(n_106), .Y(n_765) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_112), .B(n_113), .C(n_114), .Y(n_111) );
AND2x2_ASAP7_75t_L g434 ( .A(n_112), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g731 ( .A(n_113), .B(n_434), .Y(n_731) );
NOR2x2_ASAP7_75t_L g743 ( .A(n_113), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
AO221x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_745), .B1(n_748), .B2(n_757), .C(n_759), .Y(n_117) );
OAI222xp33_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_122), .B1(n_732), .B2(n_733), .C1(n_739), .C2(n_740), .Y(n_118) );
INVx1_ASAP7_75t_L g732 ( .A(n_119), .Y(n_732) );
INVxp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_124), .A2(n_431), .B1(n_436), .B2(n_729), .Y(n_123) );
INVx1_ASAP7_75t_L g735 ( .A(n_124), .Y(n_735) );
INVx2_ASAP7_75t_L g430 ( .A(n_125), .Y(n_430) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
XOR2x2_ASAP7_75t_L g752 ( .A(n_126), .B(n_753), .Y(n_752) );
AND3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_349), .C(n_397), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_277), .C(n_322), .D(n_336), .Y(n_127) );
OAI311xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_193), .A3(n_220), .B1(n_230), .C1(n_245), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_130), .B(n_157), .Y(n_129) );
OAI21xp33_ASAP7_75t_L g230 ( .A1(n_130), .A2(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g338 ( .A(n_130), .B(n_265), .Y(n_338) );
AND2x2_ASAP7_75t_L g395 ( .A(n_130), .B(n_281), .Y(n_395) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g288 ( .A(n_131), .B(n_186), .Y(n_288) );
AND2x2_ASAP7_75t_L g345 ( .A(n_131), .B(n_293), .Y(n_345) );
INVx1_ASAP7_75t_L g386 ( .A(n_131), .Y(n_386) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_132), .Y(n_254) );
AND2x2_ASAP7_75t_L g295 ( .A(n_132), .B(n_186), .Y(n_295) );
AND2x2_ASAP7_75t_L g299 ( .A(n_132), .B(n_187), .Y(n_299) );
INVx1_ASAP7_75t_L g311 ( .A(n_132), .Y(n_311) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_134), .A2(n_139), .B1(n_141), .B2(n_145), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g138 ( .A(n_136), .Y(n_138) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
AND2x6_ASAP7_75t_L g449 ( .A(n_136), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
INVx1_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_138), .Y(n_484) );
INVx2_ASAP7_75t_L g546 ( .A(n_138), .Y(n_546) );
INVx2_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_139), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_139), .A2(n_190), .B1(n_227), .B2(n_228), .Y(n_226) );
INVx4_ASAP7_75t_L g545 ( .A(n_139), .Y(n_545) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
INVx1_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
AND2x2_ASAP7_75t_L g447 ( .A(n_140), .B(n_207), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_140), .Y(n_450) );
INVx2_ASAP7_75t_L g201 ( .A(n_142), .Y(n_201) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx3_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_144), .Y(n_469) );
INVx5_ASAP7_75t_L g179 ( .A(n_145), .Y(n_179) );
INVx1_ASAP7_75t_L g456 ( .A(n_146), .Y(n_456) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_147), .A2(n_159), .B(n_169), .Y(n_158) );
OA21x2_ASAP7_75t_L g173 ( .A1(n_147), .A2(n_174), .B(n_185), .Y(n_173) );
INVx1_ASAP7_75t_L g459 ( .A(n_147), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_147), .A2(n_477), .B(n_478), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_147), .A2(n_514), .B(n_515), .Y(n_513) );
AND2x2_ASAP7_75t_SL g147 ( .A(n_148), .B(n_149), .Y(n_147) );
AND2x2_ASAP7_75t_L g156 ( .A(n_148), .B(n_149), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
NAND3xp33_ASAP7_75t_L g225 ( .A(n_152), .B(n_226), .C(n_229), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g237 ( .A1(n_152), .A2(n_238), .B(n_241), .Y(n_237) );
BUFx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_153), .A2(n_160), .B(n_165), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g174 ( .A1(n_153), .A2(n_175), .B(n_180), .Y(n_174) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_153), .A2(n_199), .B(n_204), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_153), .A2(n_213), .B(n_216), .Y(n_212) );
AND2x4_ASAP7_75t_L g446 ( .A(n_153), .B(n_447), .Y(n_446) );
INVx4_ASAP7_75t_SL g471 ( .A(n_153), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g504 ( .A(n_153), .B(n_447), .Y(n_504) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_155), .A2(n_212), .B(n_219), .Y(n_211) );
INVx4_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_155), .A2(n_494), .B(n_495), .Y(n_493) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_155), .Y(n_523) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g192 ( .A(n_156), .Y(n_192) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_170), .Y(n_157) );
AND2x2_ASAP7_75t_L g232 ( .A(n_158), .B(n_186), .Y(n_232) );
INVx2_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
AND2x2_ASAP7_75t_L g281 ( .A(n_158), .B(n_187), .Y(n_281) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_158), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_158), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g301 ( .A(n_158), .B(n_264), .Y(n_301) );
INVx1_ASAP7_75t_L g313 ( .A(n_158), .Y(n_313) );
INVx1_ASAP7_75t_L g354 ( .A(n_158), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_158), .B(n_254), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_L g241 ( .A1(n_168), .A2(n_205), .B(n_242), .C(n_243), .Y(n_241) );
NOR2xp67_ASAP7_75t_L g170 ( .A(n_171), .B(n_186), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g231 ( .A(n_172), .B(n_232), .Y(n_231) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_172), .Y(n_259) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_172), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g316 ( .A(n_172), .B(n_186), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_172), .B(n_311), .Y(n_374) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g264 ( .A(n_173), .Y(n_264) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_173), .Y(n_280) );
OR2x2_ASAP7_75t_L g353 ( .A(n_173), .B(n_354), .Y(n_353) );
O2A1O1Ixp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B(n_178), .C(n_179), .Y(n_175) );
INVx2_ASAP7_75t_L g190 ( .A(n_179), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_179), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_179), .A2(n_239), .B(n_240), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_179), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_183), .Y(n_180) );
INVx1_ASAP7_75t_L g203 ( .A(n_183), .Y(n_203) );
INVx4_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g453 ( .A(n_184), .Y(n_453) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g260 ( .A(n_187), .Y(n_260) );
AND2x2_ASAP7_75t_L g265 ( .A(n_187), .B(n_266), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_190), .A2(n_205), .B(n_208), .C(n_209), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_190), .A2(n_217), .B(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g197 ( .A(n_192), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_192), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_193), .B(n_248), .Y(n_411) );
INVx1_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_L g381 ( .A(n_194), .B(n_222), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_195), .B(n_211), .Y(n_194) );
AND2x2_ASAP7_75t_L g257 ( .A(n_195), .B(n_248), .Y(n_257) );
INVx2_ASAP7_75t_L g269 ( .A(n_195), .Y(n_269) );
AND2x2_ASAP7_75t_L g303 ( .A(n_195), .B(n_251), .Y(n_303) );
AND2x2_ASAP7_75t_L g370 ( .A(n_195), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_196), .B(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g250 ( .A(n_196), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g290 ( .A(n_196), .B(n_211), .Y(n_290) );
AND2x2_ASAP7_75t_L g307 ( .A(n_196), .B(n_308), .Y(n_307) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_210), .Y(n_196) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_197), .A2(n_237), .B(n_244), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_201), .B(n_202), .C(n_203), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_201), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_201), .A2(n_507), .B(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_203), .A2(n_467), .B(n_468), .C(n_469), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_205), .A2(n_452), .B(n_454), .Y(n_451) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g233 ( .A(n_211), .B(n_234), .Y(n_233) );
INVx3_ASAP7_75t_L g251 ( .A(n_211), .Y(n_251) );
AND2x2_ASAP7_75t_L g256 ( .A(n_211), .B(n_236), .Y(n_256) );
AND2x2_ASAP7_75t_L g329 ( .A(n_211), .B(n_308), .Y(n_329) );
AND2x2_ASAP7_75t_L g394 ( .A(n_211), .B(n_384), .Y(n_394) );
OAI311xp33_ASAP7_75t_L g277 ( .A1(n_220), .A2(n_278), .A3(n_282), .B1(n_284), .C1(n_304), .Y(n_277) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g289 ( .A(n_221), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g348 ( .A(n_221), .B(n_256), .Y(n_348) );
AND2x2_ASAP7_75t_L g422 ( .A(n_221), .B(n_303), .Y(n_422) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_222), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g357 ( .A(n_222), .Y(n_357) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx3_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
NOR2x1_ASAP7_75t_L g320 ( .A(n_223), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g377 ( .A(n_223), .B(n_251), .Y(n_377) );
AND2x4_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
INVx1_ASAP7_75t_L g274 ( .A(n_224), .Y(n_274) );
AO21x1_ASAP7_75t_L g273 ( .A1(n_226), .A2(n_229), .B(n_274), .Y(n_273) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_229), .A2(n_464), .B(n_473), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_229), .B(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_229), .B(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g501 ( .A1(n_229), .A2(n_502), .B(n_509), .Y(n_501) );
INVx3_ASAP7_75t_L g531 ( .A(n_229), .Y(n_531) );
AND2x2_ASAP7_75t_L g252 ( .A(n_232), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g305 ( .A(n_232), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g385 ( .A(n_232), .B(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_233), .A2(n_265), .B1(n_285), .B2(n_289), .C(n_291), .Y(n_284) );
INVx1_ASAP7_75t_L g409 ( .A(n_234), .Y(n_409) );
OR2x2_ASAP7_75t_L g375 ( .A(n_235), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g270 ( .A(n_236), .B(n_251), .Y(n_270) );
OR2x2_ASAP7_75t_L g272 ( .A(n_236), .B(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g297 ( .A(n_236), .Y(n_297) );
INVx2_ASAP7_75t_L g308 ( .A(n_236), .Y(n_308) );
AND2x2_ASAP7_75t_L g335 ( .A(n_236), .B(n_273), .Y(n_335) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_236), .Y(n_364) );
AOI221xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_252), .B1(n_255), .B2(n_258), .C(n_261), .Y(n_245) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
OR2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
AND2x2_ASAP7_75t_L g346 ( .A(n_248), .B(n_256), .Y(n_346) );
AND2x2_ASAP7_75t_L g396 ( .A(n_248), .B(n_250), .Y(n_396) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g283 ( .A(n_250), .B(n_254), .Y(n_283) );
AND2x2_ASAP7_75t_L g362 ( .A(n_250), .B(n_335), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_251), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g321 ( .A(n_251), .Y(n_321) );
OAI21xp33_ASAP7_75t_L g331 ( .A1(n_252), .A2(n_332), .B(n_334), .Y(n_331) );
OR2x2_ASAP7_75t_L g275 ( .A(n_253), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g341 ( .A(n_253), .B(n_301), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_253), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g318 ( .A(n_254), .B(n_287), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_254), .B(n_401), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_255), .B(n_281), .Y(n_391) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g314 ( .A(n_256), .B(n_269), .Y(n_314) );
INVx1_ASAP7_75t_L g330 ( .A(n_257), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_267), .B1(n_271), .B2(n_275), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx2_ASAP7_75t_L g293 ( .A(n_264), .Y(n_293) );
INVx1_ASAP7_75t_L g306 ( .A(n_264), .Y(n_306) );
INVx1_ASAP7_75t_L g276 ( .A(n_265), .Y(n_276) );
AND2x2_ASAP7_75t_L g347 ( .A(n_265), .B(n_293), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_265), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
OR2x2_ASAP7_75t_L g271 ( .A(n_268), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_268), .B(n_384), .Y(n_383) );
NOR2xp67_ASAP7_75t_L g415 ( .A(n_268), .B(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g418 ( .A(n_270), .B(n_370), .Y(n_418) );
INVx1_ASAP7_75t_SL g384 ( .A(n_272), .Y(n_384) );
AND2x2_ASAP7_75t_L g324 ( .A(n_273), .B(n_308), .Y(n_324) );
INVx1_ASAP7_75t_L g371 ( .A(n_273), .Y(n_371) );
OAI222xp33_ASAP7_75t_L g412 ( .A1(n_278), .A2(n_368), .B1(n_413), .B2(n_414), .C1(n_417), .C2(n_419), .Y(n_412) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_L g333 ( .A(n_280), .Y(n_333) );
AND2x2_ASAP7_75t_L g344 ( .A(n_281), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_281), .B(n_386), .Y(n_413) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_283), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g388 ( .A(n_285), .Y(n_388) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_SL g326 ( .A(n_288), .Y(n_326) );
AND2x2_ASAP7_75t_L g405 ( .A(n_288), .B(n_366), .Y(n_405) );
AND2x2_ASAP7_75t_L g428 ( .A(n_288), .B(n_312), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_290), .B(n_324), .Y(n_323) );
OAI32xp33_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_294), .A3(n_296), .B1(n_298), .B2(n_302), .Y(n_291) );
BUFx2_ASAP7_75t_L g366 ( .A(n_293), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_294), .B(n_312), .Y(n_393) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g332 ( .A(n_295), .B(n_333), .Y(n_332) );
AND2x4_ASAP7_75t_L g400 ( .A(n_295), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g389 ( .A(n_296), .B(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x2_ASAP7_75t_L g360 ( .A(n_299), .B(n_333), .Y(n_360) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
OAI221xp5_ASAP7_75t_SL g322 ( .A1(n_301), .A2(n_323), .B1(n_325), .B2(n_327), .C(n_331), .Y(n_322) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g334 ( .A(n_303), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g340 ( .A(n_303), .B(n_324), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_307), .B1(n_309), .B2(n_314), .C(n_315), .Y(n_304) );
INVx1_ASAP7_75t_L g423 ( .A(n_305), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_306), .B(n_400), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_307), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_312), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g378 ( .A(n_312), .Y(n_378) );
BUFx3_ASAP7_75t_L g401 ( .A(n_313), .Y(n_401) );
INVx1_ASAP7_75t_SL g342 ( .A(n_314), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_314), .B(n_356), .Y(n_355) );
AOI21xp33_ASAP7_75t_SL g315 ( .A1(n_316), .A2(n_317), .B(n_319), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_316), .A2(n_417), .B1(n_421), .B2(n_423), .C(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g363 ( .A(n_321), .B(n_324), .Y(n_363) );
INVx1_ASAP7_75t_L g427 ( .A(n_321), .Y(n_427) );
INVx2_ASAP7_75t_L g416 ( .A(n_324), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_324), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_370), .Y(n_369) );
OAI221xp5_ASAP7_75t_SL g336 ( .A1(n_337), .A2(n_339), .B1(n_341), .B2(n_342), .C(n_343), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g339 ( .A(n_340), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_346), .B1(n_347), .B2(n_348), .Y(n_343) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_345), .A2(n_407), .B1(n_408), .B2(n_410), .Y(n_406) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_348), .A2(n_425), .B(n_428), .Y(n_424) );
NOR4xp25_ASAP7_75t_SL g349 ( .A(n_350), .B(n_358), .C(n_367), .D(n_387), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .B1(n_364), .B2(n_365), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_372), .B1(n_375), .B2(n_378), .C(n_379), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g390 ( .A(n_370), .Y(n_390) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI21xp5_ASAP7_75t_SL g379 ( .A1(n_380), .A2(n_382), .B(n_385), .Y(n_379) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_391), .C(n_392), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_395), .B2(n_396), .Y(n_392) );
CKINVDCx14_ASAP7_75t_R g402 ( .A(n_396), .Y(n_402) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_412), .C(n_420), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B1(n_403), .B2(n_404), .C(n_406), .Y(n_398) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g736 ( .A(n_432), .Y(n_736) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g744 ( .A(n_434), .Y(n_744) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g737 ( .A(n_437), .Y(n_737) );
AND3x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_633), .C(n_690), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_578), .C(n_614), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_487), .B(n_533), .C(n_565), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_460), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g536 ( .A(n_442), .B(n_537), .Y(n_536) );
INVx5_ASAP7_75t_L g564 ( .A(n_442), .Y(n_564) );
AND2x2_ASAP7_75t_L g637 ( .A(n_442), .B(n_553), .Y(n_637) );
AND2x2_ASAP7_75t_L g675 ( .A(n_442), .B(n_581), .Y(n_675) );
AND2x2_ASAP7_75t_L g695 ( .A(n_442), .B(n_538), .Y(n_695) );
OR2x6_ASAP7_75t_L g442 ( .A(n_443), .B(n_457), .Y(n_442) );
AOI21xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_448), .B(n_456), .Y(n_443) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx5_ASAP7_75t_L g480 ( .A(n_449), .Y(n_480) );
INVx2_ASAP7_75t_L g455 ( .A(n_453), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_455), .A2(n_482), .B(n_483), .C(n_484), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_455), .A2(n_484), .B(n_517), .C(n_518), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_460), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_475), .Y(n_460) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_461), .Y(n_576) );
AND2x2_ASAP7_75t_L g590 ( .A(n_461), .B(n_537), .Y(n_590) );
INVx1_ASAP7_75t_L g613 ( .A(n_461), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_461), .B(n_564), .Y(n_652) );
OR2x2_ASAP7_75t_L g689 ( .A(n_461), .B(n_535), .Y(n_689) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_462), .Y(n_625) );
AND2x2_ASAP7_75t_L g632 ( .A(n_462), .B(n_538), .Y(n_632) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g553 ( .A(n_463), .B(n_538), .Y(n_553) );
BUFx2_ASAP7_75t_L g581 ( .A(n_463), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_472), .Y(n_464) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g525 ( .A1(n_471), .A2(n_480), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_SL g540 ( .A1(n_471), .A2(n_480), .B(n_541), .C(n_542), .Y(n_540) );
INVx5_ASAP7_75t_L g535 ( .A(n_475), .Y(n_535) );
BUFx2_ASAP7_75t_L g557 ( .A(n_475), .Y(n_557) );
AND2x2_ASAP7_75t_L g714 ( .A(n_475), .B(n_568), .Y(n_714) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_520), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_489), .A2(n_615), .B1(n_622), .B2(n_623), .C(n_626), .Y(n_614) );
OR2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
AND2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_490), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g549 ( .A(n_491), .B(n_500), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_491), .B(n_501), .Y(n_559) );
OR2x2_ASAP7_75t_L g570 ( .A(n_491), .B(n_522), .Y(n_570) );
AND2x2_ASAP7_75t_L g573 ( .A(n_491), .B(n_561), .Y(n_573) );
AND2x2_ASAP7_75t_L g589 ( .A(n_491), .B(n_511), .Y(n_589) );
OR2x2_ASAP7_75t_L g605 ( .A(n_491), .B(n_501), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_491), .B(n_522), .Y(n_667) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_492), .B(n_511), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_492), .B(n_501), .Y(n_662) );
OR2x2_ASAP7_75t_L g583 ( .A(n_499), .B(n_570), .Y(n_583) );
INVx2_ASAP7_75t_L g609 ( .A(n_499), .Y(n_609) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
AND2x2_ASAP7_75t_L g532 ( .A(n_500), .B(n_512), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_500), .B(n_522), .Y(n_588) );
OR2x2_ASAP7_75t_L g599 ( .A(n_500), .B(n_512), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_500), .B(n_561), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_500), .A2(n_692), .B1(n_694), .B2(n_696), .C(n_699), .Y(n_691) );
INVx5_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_501), .B(n_522), .Y(n_630) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_505), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_511), .B(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_511), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g577 ( .A(n_511), .B(n_549), .Y(n_577) );
OR2x2_ASAP7_75t_L g621 ( .A(n_511), .B(n_522), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_511), .B(n_573), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_511), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g686 ( .A(n_511), .B(n_687), .Y(n_686) );
INVx5_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_SL g550 ( .A(n_512), .B(n_521), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_SL g554 ( .A1(n_512), .A2(n_555), .B(n_558), .C(n_562), .Y(n_554) );
OR2x2_ASAP7_75t_L g592 ( .A(n_512), .B(n_588), .Y(n_592) );
OR2x2_ASAP7_75t_L g628 ( .A(n_512), .B(n_570), .Y(n_628) );
OAI311xp33_ASAP7_75t_L g634 ( .A1(n_512), .A2(n_573), .A3(n_635), .B1(n_638), .C1(n_645), .Y(n_634) );
AND2x2_ASAP7_75t_L g685 ( .A(n_512), .B(n_522), .Y(n_685) );
AND2x2_ASAP7_75t_L g693 ( .A(n_512), .B(n_548), .Y(n_693) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_512), .Y(n_711) );
AND2x2_ASAP7_75t_L g728 ( .A(n_512), .B(n_549), .Y(n_728) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_532), .Y(n_520) );
AND2x2_ASAP7_75t_L g556 ( .A(n_521), .B(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g712 ( .A(n_521), .Y(n_712) );
AND2x2_ASAP7_75t_L g548 ( .A(n_522), .B(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g561 ( .A(n_522), .Y(n_561) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_522), .Y(n_604) );
INVxp67_ASAP7_75t_L g643 ( .A(n_522), .Y(n_643) );
OA21x2_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_530), .Y(n_522) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_531), .A2(n_539), .B(n_547), .Y(n_538) );
AND2x2_ASAP7_75t_L g721 ( .A(n_532), .B(n_569), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_548), .B1(n_550), .B2(n_551), .C(n_554), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_535), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g574 ( .A(n_535), .B(n_564), .Y(n_574) );
AND2x2_ASAP7_75t_L g582 ( .A(n_535), .B(n_537), .Y(n_582) );
OR2x2_ASAP7_75t_L g594 ( .A(n_535), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g612 ( .A(n_535), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g636 ( .A(n_535), .B(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_535), .Y(n_656) );
AND2x2_ASAP7_75t_L g708 ( .A(n_535), .B(n_632), .Y(n_708) );
OAI31xp33_ASAP7_75t_L g716 ( .A1(n_535), .A2(n_585), .A3(n_684), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_536), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g680 ( .A(n_536), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_536), .B(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_L g568 ( .A(n_537), .B(n_564), .Y(n_568) );
INVx1_ASAP7_75t_L g655 ( .A(n_537), .Y(n_655) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g705 ( .A(n_538), .B(n_564), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_SL g715 ( .A(n_548), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_549), .B(n_620), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_550), .A2(n_662), .B1(n_700), .B2(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g563 ( .A(n_553), .B(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g622 ( .A(n_553), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_553), .B(n_574), .Y(n_727) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g697 ( .A(n_556), .B(n_698), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_557), .A2(n_616), .B(n_618), .Y(n_615) );
OR2x2_ASAP7_75t_L g623 ( .A(n_557), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g644 ( .A(n_557), .B(n_632), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_557), .B(n_655), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_557), .B(n_695), .Y(n_694) );
OAI221xp5_ASAP7_75t_SL g671 ( .A1(n_558), .A2(n_672), .B1(n_677), .B2(n_680), .C(n_681), .Y(n_671) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
OR2x2_ASAP7_75t_L g648 ( .A(n_559), .B(n_621), .Y(n_648) );
INVx1_ASAP7_75t_L g687 ( .A(n_559), .Y(n_687) );
INVx2_ASAP7_75t_L g663 ( .A(n_560), .Y(n_663) );
INVx1_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g602 ( .A(n_564), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_564), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g631 ( .A(n_564), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g719 ( .A(n_564), .B(n_689), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_569), .B1(n_571), .B2(n_574), .C1(n_575), .C2(n_577), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g575 ( .A(n_568), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_568), .A2(n_618), .B1(n_646), .B2(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_568), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_577), .A2(n_607), .B(n_610), .Y(n_606) );
OAI211xp5_ASAP7_75t_SL g578 ( .A1(n_579), .A2(n_583), .B(n_584), .C(n_606), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_582), .A2(n_585), .B1(n_590), .B2(n_591), .C(n_593), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_582), .B(n_670), .Y(n_669) );
INVxp67_ASAP7_75t_L g676 ( .A(n_582), .Y(n_676) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
AND2x2_ASAP7_75t_L g678 ( .A(n_587), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g595 ( .A(n_590), .Y(n_595) );
AND2x2_ASAP7_75t_L g601 ( .A(n_590), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B1(n_600), .B2(n_603), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_597), .B(n_609), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_598), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g698 ( .A(n_602), .Y(n_698) );
AND2x2_ASAP7_75t_L g717 ( .A(n_602), .B(n_632), .Y(n_717) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_609), .B(n_666), .Y(n_725) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_612), .B(n_680), .Y(n_723) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g646 ( .A(n_624), .Y(n_646) );
BUFx2_ASAP7_75t_L g670 ( .A(n_625), .Y(n_670) );
OAI21xp5_ASAP7_75t_SL g626 ( .A1(n_627), .A2(n_629), .B(n_631), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NOR3xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_649), .C(n_671), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B(n_644), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_653), .B(n_657), .C(n_660), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_650), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp67_ASAP7_75t_SL g654 ( .A(n_655), .B(n_656), .Y(n_654) );
OR2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_SL g679 ( .A(n_659), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_664), .B(n_668), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g684 ( .A(n_662), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_684), .B1(n_686), .B2(n_688), .Y(n_681) );
INVx2_ASAP7_75t_SL g702 ( .A(n_689), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_691), .B(n_706), .C(n_718), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_702), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B1(n_713), .B2(n_715), .C(n_716), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_707), .A2(n_719), .B(n_720), .C(n_722), .Y(n_718) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVxp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B1(n_726), .B2(n_728), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g738 ( .A(n_730), .Y(n_738) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI22xp5_ASAP7_75t_SL g734 ( .A1(n_735), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_734) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
BUFx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g758 ( .A(n_746), .Y(n_758) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g762 ( .A(n_750), .Y(n_762) );
INVx1_ASAP7_75t_L g755 ( .A(n_752), .Y(n_755) );
BUFx3_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
endmodule