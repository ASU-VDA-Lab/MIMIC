module fake_aes_7248_n_887 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_887);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_887;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_638;
wire n_540;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_529;
wire n_455;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx8_ASAP7_75t_SL g110 ( .A(n_38), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_76), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_82), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_89), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_33), .Y(n_114) );
BUFx10_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_9), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_65), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_49), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_54), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_95), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_39), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_106), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_3), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_88), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_9), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_96), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_45), .Y(n_128) );
INVx1_ASAP7_75t_SL g129 ( .A(n_66), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_108), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_5), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_57), .Y(n_134) );
OR2x2_ASAP7_75t_L g135 ( .A(n_85), .B(n_23), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_75), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_7), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_27), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_15), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_55), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_78), .Y(n_141) );
INVx1_ASAP7_75t_SL g142 ( .A(n_37), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_105), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_21), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_101), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_35), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_109), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_17), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_15), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_137), .Y(n_151) );
OAI22x1_ASAP7_75t_R g152 ( .A1(n_126), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_144), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_144), .B(n_19), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_110), .Y(n_155) );
INVx5_ASAP7_75t_L g156 ( .A(n_125), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_115), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
BUFx12f_ASAP7_75t_L g159 ( .A(n_115), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
OAI22x1_ASAP7_75t_SL g161 ( .A1(n_137), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_130), .A2(n_52), .B(n_103), .Y(n_163) );
INVx5_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_127), .Y(n_166) );
HB1xp67_ASAP7_75t_L g167 ( .A(n_148), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_132), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_123), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_115), .B(n_3), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_135), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_155), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_159), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_159), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_151), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g182 ( .A1(n_152), .A2(n_148), .B1(n_114), .B2(n_124), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_167), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_153), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_164), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_164), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_164), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
NAND2xp33_ASAP7_75t_R g189 ( .A(n_174), .B(n_116), .Y(n_189) );
NOR2xp67_ASAP7_75t_L g190 ( .A(n_157), .B(n_149), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_164), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_164), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_157), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_176), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_150), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_174), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_152), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_161), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_161), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_165), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_165), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_176), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_176), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_153), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_176), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_176), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_153), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_176), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_166), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_175), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_166), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_175), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_154), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_169), .Y(n_218) );
INVx3_ASAP7_75t_L g219 ( .A(n_171), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_154), .Y(n_220) );
AND2x6_ASAP7_75t_L g221 ( .A(n_169), .B(n_129), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_170), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_170), .Y(n_223) );
INVxp67_ASAP7_75t_L g224 ( .A(n_169), .Y(n_224) );
BUFx10_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_160), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_170), .B(n_111), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_160), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_173), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_171), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g231 ( .A(n_216), .B(n_154), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_222), .B(n_111), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_223), .B(n_112), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_225), .Y(n_234) );
BUFx8_ASAP7_75t_L g235 ( .A(n_221), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_212), .B(n_113), .Y(n_236) );
INVxp67_ASAP7_75t_L g237 ( .A(n_227), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_214), .B(n_113), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_227), .B(n_136), .Y(n_239) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_215), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_229), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_188), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_202), .B(n_136), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_203), .B(n_118), .Y(n_244) );
BUFx6f_ASAP7_75t_SL g245 ( .A(n_221), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_194), .B(n_162), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_190), .B(n_162), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_213), .B(n_154), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_181), .B(n_168), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_196), .Y(n_250) );
INVxp67_ASAP7_75t_SL g251 ( .A(n_220), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_183), .B(n_168), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_220), .B(n_154), .Y(n_253) );
INVxp67_ASAP7_75t_L g254 ( .A(n_189), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_225), .B(n_120), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_198), .A2(n_154), .B1(n_173), .B2(n_171), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_224), .B(n_121), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_205), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_195), .B(n_142), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_208), .B(n_171), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_178), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_211), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
NOR3xp33_ASAP7_75t_L g265 ( .A(n_182), .B(n_163), .C(n_128), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_198), .A2(n_172), .B1(n_171), .B2(n_145), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_204), .Y(n_267) );
NOR2xp33_ASAP7_75t_SL g268 ( .A(n_179), .B(n_122), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_206), .B(n_131), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_184), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_209), .B(n_134), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_185), .B(n_140), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_186), .B(n_141), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_187), .B(n_143), .Y(n_274) );
INVx1_ASAP7_75t_SL g275 ( .A(n_180), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_192), .B(n_147), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_230), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_184), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_189), .A2(n_172), .B1(n_158), .B2(n_156), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_193), .B(n_172), .Y(n_280) );
AO221x1_ASAP7_75t_L g281 ( .A1(n_199), .A2(n_172), .B1(n_160), .B2(n_163), .C(n_7), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_177), .B(n_172), .Y(n_282) );
NOR3xp33_ASAP7_75t_L g283 ( .A(n_200), .B(n_4), .C(n_5), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_221), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_221), .B(n_201), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_221), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_217), .B(n_156), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_217), .B(n_156), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_191), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_235), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_240), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_240), .B(n_199), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_231), .B(n_177), .Y(n_293) );
NOR2x2_ASAP7_75t_L g294 ( .A(n_262), .B(n_268), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_260), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_241), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_250), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_237), .B(n_156), .Y(n_300) );
NAND2xp33_ASAP7_75t_L g301 ( .A(n_234), .B(n_177), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_237), .B(n_156), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_265), .A2(n_172), .B1(n_158), .B2(n_156), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_252), .B(n_158), .Y(n_304) );
BUFx3_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_246), .B(n_158), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_263), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_249), .B(n_158), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_265), .A2(n_160), .B(n_197), .C(n_191), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_254), .A2(n_232), .B1(n_233), .B2(n_236), .Y(n_310) );
NOR2x1p5_ASAP7_75t_L g311 ( .A(n_285), .B(n_160), .Y(n_311) );
AND2x2_ASAP7_75t_SL g312 ( .A(n_253), .B(n_160), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_238), .B(n_158), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_239), .B(n_197), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_254), .B(n_6), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_253), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_275), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_234), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_234), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_234), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_256), .B(n_177), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_264), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_244), .B(n_6), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_281), .A2(n_219), .B1(n_210), .B2(n_207), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_270), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_264), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_266), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_283), .B(n_8), .Y(n_329) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_248), .A2(n_210), .B(n_207), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_264), .B(n_219), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_264), .B(n_226), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_267), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_278), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g336 ( .A1(n_291), .A2(n_283), .B1(n_247), .B2(n_279), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_316), .B(n_284), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g338 ( .A1(n_309), .A2(n_251), .B(n_286), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_322), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_317), .B(n_269), .Y(n_340) );
OR2x6_ASAP7_75t_SL g341 ( .A(n_294), .B(n_245), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_322), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_322), .B(n_257), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_325), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_297), .B(n_247), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_322), .B(n_280), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_325), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_298), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_334), .Y(n_349) );
BUFx12f_ASAP7_75t_L g350 ( .A(n_290), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_322), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_326), .B(n_271), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_310), .B(n_273), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_296), .B(n_277), .Y(n_354) );
NOR3xp33_ASAP7_75t_SL g355 ( .A(n_292), .B(n_274), .C(n_276), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_316), .B(n_272), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_290), .Y(n_357) );
O2A1O1Ixp5_ASAP7_75t_L g358 ( .A1(n_293), .A2(n_255), .B(n_259), .C(n_261), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_315), .A2(n_245), .B1(n_259), .B2(n_251), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_312), .B(n_287), .Y(n_360) );
CKINVDCx11_ASAP7_75t_R g361 ( .A(n_305), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_305), .B(n_288), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_344), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_361), .Y(n_365) );
BUFx8_ASAP7_75t_L g366 ( .A(n_350), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_342), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_335), .B(n_299), .Y(n_369) );
AND2x4_ASAP7_75t_L g370 ( .A(n_351), .B(n_333), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_335), .Y(n_371) );
BUFx12f_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_351), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_339), .B(n_319), .Y(n_374) );
OAI21x1_ASAP7_75t_SL g375 ( .A1(n_338), .A2(n_324), .B(n_349), .Y(n_375) );
OAI21x1_ASAP7_75t_L g376 ( .A1(n_358), .A2(n_293), .B(n_321), .Y(n_376) );
OAI21x1_ASAP7_75t_SL g377 ( .A1(n_344), .A2(n_303), .B(n_333), .Y(n_377) );
OR2x6_ASAP7_75t_L g378 ( .A(n_339), .B(n_315), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
INVxp67_ASAP7_75t_SL g380 ( .A(n_363), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_348), .B(n_315), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_347), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_357), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_353), .A2(n_306), .B(n_321), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_347), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_362), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_336), .B(n_329), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_354), .Y(n_390) );
INVx1_ASAP7_75t_SL g391 ( .A(n_363), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_354), .Y(n_392) );
INVx5_ASAP7_75t_L g393 ( .A(n_357), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_343), .A2(n_330), .B(n_332), .Y(n_394) );
OAI21x1_ASAP7_75t_L g395 ( .A1(n_346), .A2(n_332), .B(n_318), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_362), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_393), .Y(n_397) );
BUFx3_ASAP7_75t_L g398 ( .A(n_366), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
CKINVDCx11_ASAP7_75t_R g400 ( .A(n_372), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_392), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_388), .A2(n_336), .B1(n_323), .B2(n_345), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_393), .A2(n_323), .B1(n_294), .B2(n_341), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_371), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_379), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_379), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_386), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_390), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_393), .Y(n_414) );
OAI21x1_ASAP7_75t_L g415 ( .A1(n_376), .A2(n_318), .B(n_346), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_378), .A2(n_341), .B1(n_359), .B2(n_323), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_392), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_383), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_378), .A2(n_328), .B1(n_308), .B2(n_309), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_378), .A2(n_352), .B1(n_311), .B2(n_340), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_390), .B(n_345), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
BUFx12f_ASAP7_75t_L g424 ( .A(n_366), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_369), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_386), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_389), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_383), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_394), .Y(n_429) );
OAI22x1_ASAP7_75t_L g430 ( .A1(n_393), .A2(n_362), .B1(n_346), .B2(n_356), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_385), .A2(n_304), .B(n_300), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
BUFx4f_ASAP7_75t_L g433 ( .A(n_378), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
INVx5_ASAP7_75t_L g435 ( .A(n_393), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_370), .A2(n_304), .B1(n_355), .B2(n_362), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_381), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_387), .B(n_337), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_375), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_375), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_387), .A2(n_337), .B1(n_360), .B2(n_302), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_396), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_366), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_387), .A2(n_337), .B1(n_313), .B2(n_307), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_370), .B(n_337), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g447 ( .A1(n_380), .A2(n_337), .B1(n_307), .B2(n_327), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_435), .B(n_368), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_406), .B(n_391), .C(n_365), .Y(n_450) );
BUFx10_ASAP7_75t_L g451 ( .A(n_424), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_427), .B(n_391), .Y(n_452) );
OR2x6_ASAP7_75t_L g453 ( .A(n_424), .B(n_372), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_402), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_444), .Y(n_455) );
NOR2xp33_ASAP7_75t_R g456 ( .A(n_444), .B(n_366), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_413), .B(n_368), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_398), .B(n_370), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_435), .Y(n_459) );
NAND2xp33_ASAP7_75t_R g460 ( .A(n_400), .B(n_393), .Y(n_460) );
BUFx12f_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_398), .Y(n_462) );
AND3x2_ASAP7_75t_L g463 ( .A(n_435), .B(n_372), .C(n_370), .Y(n_463) );
XOR2xp5_ASAP7_75t_L g464 ( .A(n_416), .B(n_384), .Y(n_464) );
NAND2xp33_ASAP7_75t_R g465 ( .A(n_435), .B(n_367), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_425), .B(n_368), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_419), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_433), .A2(n_377), .B1(n_373), .B2(n_382), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_407), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_408), .B(n_367), .Y(n_471) );
CKINVDCx9p33_ASAP7_75t_R g472 ( .A(n_422), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_401), .B(n_373), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_411), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_404), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_409), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_433), .A2(n_382), .B1(n_367), .B2(n_384), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_433), .A2(n_382), .B1(n_367), .B2(n_377), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g479 ( .A1(n_405), .A2(n_318), .B(n_319), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_417), .B(n_8), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_411), .B(n_10), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_404), .Y(n_482) );
NOR3xp33_ASAP7_75t_SL g483 ( .A(n_421), .B(n_282), .C(n_314), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_410), .Y(n_484) );
NAND2xp33_ASAP7_75t_R g485 ( .A(n_399), .B(n_10), .Y(n_485) );
NOR2x1_ASAP7_75t_SL g486 ( .A(n_414), .B(n_319), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_397), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_431), .A2(n_376), .B(n_261), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_432), .B(n_11), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_399), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_430), .Y(n_491) );
INVxp33_ASAP7_75t_L g492 ( .A(n_446), .Y(n_492) );
AND3x2_ASAP7_75t_L g493 ( .A(n_446), .B(n_11), .C(n_12), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_432), .B(n_12), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_438), .B(n_334), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_426), .B(n_13), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_410), .Y(n_497) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_439), .Y(n_499) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_439), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_399), .B(n_319), .Y(n_501) );
BUFx3_ASAP7_75t_L g502 ( .A(n_403), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_403), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_443), .B(n_13), .Y(n_504) );
NAND3xp33_ASAP7_75t_SL g505 ( .A(n_436), .B(n_14), .C(n_16), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_420), .A2(n_327), .B1(n_320), .B2(n_301), .Y(n_506) );
CKINVDCx12_ASAP7_75t_R g507 ( .A(n_412), .Y(n_507) );
AO31x2_ASAP7_75t_L g508 ( .A1(n_429), .A2(n_228), .A3(n_226), .B(n_289), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_443), .B(n_14), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_430), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_412), .B(n_16), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_403), .B(n_17), .Y(n_512) );
AND2x6_ASAP7_75t_SL g513 ( .A(n_440), .B(n_18), .Y(n_513) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_447), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g515 ( .A1(n_442), .A2(n_327), .B1(n_320), .B2(n_331), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_423), .A2(n_327), .B1(n_320), .B2(n_301), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_418), .A2(n_331), .B(n_320), .Y(n_517) );
NOR2xp33_ASAP7_75t_R g518 ( .A(n_423), .B(n_18), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_418), .B(n_20), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_423), .Y(n_520) );
NAND2x1_ASAP7_75t_L g521 ( .A(n_428), .B(n_228), .Y(n_521) );
NOR2xp33_ASAP7_75t_R g522 ( .A(n_428), .B(n_22), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_440), .B(n_24), .Y(n_523) );
BUFx2_ASAP7_75t_L g524 ( .A(n_415), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_441), .B(n_25), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_441), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_415), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_445), .Y(n_528) );
BUFx3_ASAP7_75t_L g529 ( .A(n_437), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_437), .B(n_26), .Y(n_530) );
NAND2xp33_ASAP7_75t_R g531 ( .A(n_448), .B(n_28), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_467), .B(n_434), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_499), .B(n_434), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_482), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_454), .B(n_429), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_485), .A2(n_29), .B1(n_30), .B2(n_31), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_498), .B(n_32), .Y(n_537) );
INVx3_ASAP7_75t_L g538 ( .A(n_459), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_492), .B(n_34), .Y(n_539) );
NOR4xp25_ASAP7_75t_SL g540 ( .A(n_460), .B(n_36), .C(n_40), .D(n_41), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_468), .B(n_42), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_497), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_452), .B(n_43), .Y(n_543) );
INVx4_ASAP7_75t_L g544 ( .A(n_463), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_473), .B(n_44), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_474), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_458), .B(n_46), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_457), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_462), .B(n_47), .Y(n_549) );
INVx5_ASAP7_75t_L g550 ( .A(n_453), .Y(n_550) );
AND2x4_ASAP7_75t_SL g551 ( .A(n_453), .B(n_48), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_471), .B(n_50), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_466), .B(n_51), .Y(n_553) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_453), .B(n_450), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_475), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_484), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_498), .B(n_53), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_498), .B(n_56), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_459), .B(n_58), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_470), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_471), .B(n_59), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_476), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_526), .B(n_60), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_489), .B(n_61), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_529), .Y(n_566) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_449), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_496), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_494), .B(n_62), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_481), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_500), .B(n_63), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_527), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_495), .Y(n_576) );
BUFx2_ASAP7_75t_L g577 ( .A(n_472), .Y(n_577) );
CKINVDCx14_ASAP7_75t_R g578 ( .A(n_456), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_500), .B(n_64), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_487), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_500), .B(n_449), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_524), .Y(n_582) );
OAI211xp5_ASAP7_75t_SL g583 ( .A1(n_483), .A2(n_67), .B(n_68), .C(n_69), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_495), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_509), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_480), .B(n_70), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_514), .B(n_71), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_464), .Y(n_588) );
INVx3_ASAP7_75t_L g589 ( .A(n_523), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_508), .Y(n_590) );
NAND4xp25_ASAP7_75t_L g591 ( .A(n_450), .B(n_72), .C(n_73), .D(n_74), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_502), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_503), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_525), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_491), .B(n_77), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_455), .B(n_79), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_490), .B(n_80), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_510), .B(n_83), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_451), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_490), .B(n_84), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_512), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_520), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_528), .B(n_86), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_477), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_479), .B(n_87), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_518), .B(n_90), .Y(n_607) );
INVx2_ASAP7_75t_SL g608 ( .A(n_451), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_501), .B(n_91), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_477), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_508), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_501), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_508), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_486), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_530), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_479), .B(n_92), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_478), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_478), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_519), .B(n_93), .Y(n_619) );
INVx4_ASAP7_75t_L g620 ( .A(n_461), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_521), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_515), .B(n_94), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_515), .B(n_97), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_483), .B(n_98), .Y(n_624) );
INVx3_ASAP7_75t_L g625 ( .A(n_513), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_469), .B(n_99), .Y(n_626) );
BUFx3_ASAP7_75t_L g627 ( .A(n_465), .Y(n_627) );
NAND2x1_ASAP7_75t_L g628 ( .A(n_531), .B(n_100), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_469), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_505), .Y(n_630) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_517), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_506), .B(n_104), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_522), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_505), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_506), .B(n_493), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_488), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_517), .B(n_488), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_516), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_516), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_467), .B(n_499), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_548), .B(n_640), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_542), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_548), .B(n_581), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_532), .B(n_542), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_576), .B(n_584), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_534), .B(n_546), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_629), .B(n_561), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_566), .B(n_561), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_533), .B(n_566), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_577), .B(n_554), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_633), .B(n_550), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_567), .B(n_571), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_555), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_636), .B(n_563), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_568), .B(n_570), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_567), .B(n_603), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_605), .B(n_610), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_556), .B(n_572), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_535), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_593), .B(n_574), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_585), .B(n_558), .Y(n_661) );
BUFx3_ASAP7_75t_L g662 ( .A(n_550), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_617), .B(n_618), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_627), .B(n_550), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_558), .B(n_612), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_535), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_575), .Y(n_667) );
AND2x4_ASAP7_75t_SL g668 ( .A(n_544), .B(n_589), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_639), .B(n_575), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_638), .B(n_630), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_611), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_612), .B(n_588), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_592), .B(n_589), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_594), .B(n_538), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_594), .B(n_538), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_627), .B(n_550), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_614), .Y(n_677) );
INVx1_ASAP7_75t_SL g678 ( .A(n_600), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_625), .A2(n_602), .B1(n_634), .B2(n_578), .C(n_635), .Y(n_679) );
NAND2x1_ASAP7_75t_SL g680 ( .A(n_544), .B(n_625), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_580), .B(n_615), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_564), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_582), .B(n_631), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_613), .Y(n_684) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_608), .B(n_591), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_578), .B(n_595), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_582), .B(n_631), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_637), .B(n_635), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_580), .B(n_543), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_587), .B(n_596), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_637), .B(n_600), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_637), .B(n_545), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_541), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_549), .B(n_539), .Y(n_694) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_591), .A2(n_628), .B1(n_536), .B2(n_587), .C(n_606), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_590), .B(n_624), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_604), .B(n_596), .C(n_599), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_552), .Y(n_698) );
AND2x2_ASAP7_75t_L g699 ( .A(n_547), .B(n_553), .Y(n_699) );
AND2x4_ASAP7_75t_L g700 ( .A(n_551), .B(n_621), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_606), .B(n_616), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_562), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_586), .B(n_573), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_597), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_559), .B(n_599), .Y(n_705) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_616), .B(n_626), .C(n_583), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g707 ( .A(n_626), .B(n_583), .C(n_632), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_609), .B(n_620), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_620), .B(n_607), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_622), .B(n_623), .Y(n_710) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_560), .Y(n_711) );
NAND3xp33_ASAP7_75t_L g712 ( .A(n_632), .B(n_569), .C(n_565), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_537), .B(n_557), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_598), .Y(n_714) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_601), .Y(n_715) );
INVxp67_ASAP7_75t_L g716 ( .A(n_565), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_537), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_579), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_569), .B(n_557), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_619), .Y(n_720) );
OR2x2_ASAP7_75t_L g721 ( .A(n_540), .B(n_548), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_540), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_548), .B(n_640), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_548), .B(n_542), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_548), .B(n_640), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_548), .B(n_542), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_627), .B(n_566), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_548), .B(n_640), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_542), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_548), .B(n_640), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_576), .B(n_584), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_548), .B(n_542), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_548), .B(n_640), .Y(n_733) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_668), .B(n_727), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_670), .B(n_647), .Y(n_735) );
BUFx2_ASAP7_75t_L g736 ( .A(n_678), .Y(n_736) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_642), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_643), .B(n_644), .Y(n_738) );
AND2x4_ASAP7_75t_SL g739 ( .A(n_700), .B(n_727), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_665), .B(n_649), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_657), .B(n_688), .Y(n_741) );
OR2x6_ASAP7_75t_L g742 ( .A(n_650), .B(n_685), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_670), .B(n_647), .Y(n_743) );
BUFx2_ASAP7_75t_L g744 ( .A(n_642), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_657), .B(n_663), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_724), .B(n_726), .Y(n_746) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_667), .Y(n_747) );
AND2x2_ASAP7_75t_L g748 ( .A(n_688), .B(n_663), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_673), .B(n_660), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_659), .B(n_666), .Y(n_750) );
AND2x4_ASAP7_75t_L g751 ( .A(n_691), .B(n_674), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_675), .B(n_672), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_732), .B(n_646), .Y(n_753) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_667), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_652), .B(n_696), .Y(n_755) );
AND2x2_ASAP7_75t_L g756 ( .A(n_696), .B(n_661), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_641), .B(n_723), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_725), .B(n_728), .Y(n_758) );
AND2x2_ASAP7_75t_L g759 ( .A(n_730), .B(n_733), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_669), .B(n_653), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_650), .B(n_679), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_669), .B(n_729), .Y(n_762) );
BUFx3_ASAP7_75t_L g763 ( .A(n_700), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_686), .Y(n_764) );
OR2x2_ASAP7_75t_L g765 ( .A(n_658), .B(n_648), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g766 ( .A(n_679), .B(n_697), .C(n_690), .D(n_695), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_655), .B(n_645), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_716), .B(n_654), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_654), .Y(n_769) );
AND2x2_ASAP7_75t_L g770 ( .A(n_692), .B(n_677), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_690), .B(n_716), .Y(n_771) );
INVx4_ASAP7_75t_L g772 ( .A(n_662), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_706), .A2(n_707), .B1(n_701), .B2(n_712), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_656), .Y(n_774) );
INVx1_ASAP7_75t_SL g775 ( .A(n_708), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_683), .B(n_687), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_645), .B(n_731), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_683), .B(n_687), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_681), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_651), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_671), .B(n_684), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_671), .B(n_720), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_682), .B(n_693), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_715), .B(n_704), .Y(n_784) );
INVx4_ASAP7_75t_L g785 ( .A(n_662), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_715), .B(n_714), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_698), .B(n_702), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_651), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_751), .B(n_689), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_777), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_751), .B(n_709), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_744), .Y(n_792) );
O2A1O1Ixp5_ASAP7_75t_R g793 ( .A1(n_783), .A2(n_701), .B(n_719), .C(n_680), .Y(n_793) );
NOR2x1p5_ASAP7_75t_L g794 ( .A(n_766), .B(n_711), .Y(n_794) );
NOR2x1p5_ASAP7_75t_SL g795 ( .A(n_780), .B(n_721), .Y(n_795) );
OAI22xp33_ASAP7_75t_L g796 ( .A1(n_742), .A2(n_695), .B1(n_711), .B2(n_710), .Y(n_796) );
OR2x2_ASAP7_75t_L g797 ( .A(n_765), .B(n_718), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_769), .Y(n_798) );
INVx1_ASAP7_75t_SL g799 ( .A(n_736), .Y(n_799) );
AND2x2_ASAP7_75t_L g800 ( .A(n_751), .B(n_668), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_767), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_781), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_760), .Y(n_803) );
INVx2_ASAP7_75t_SL g804 ( .A(n_739), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_739), .B(n_664), .Y(n_805) );
NOR3xp33_ASAP7_75t_SL g806 ( .A(n_761), .B(n_722), .C(n_719), .Y(n_806) );
INVx1_ASAP7_75t_SL g807 ( .A(n_734), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_760), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_750), .Y(n_809) );
INVx1_ASAP7_75t_SL g810 ( .A(n_734), .Y(n_810) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_764), .B(n_775), .Y(n_811) );
NOR2x1p5_ASAP7_75t_L g812 ( .A(n_763), .B(n_664), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_761), .A2(n_676), .B1(n_699), .B2(n_705), .Y(n_813) );
OAI322xp33_ASAP7_75t_L g814 ( .A1(n_771), .A2(n_676), .A3(n_694), .B1(n_703), .B2(n_713), .C1(n_717), .C2(n_735), .Y(n_814) );
NAND4xp75_ASAP7_75t_SL g815 ( .A(n_742), .B(n_771), .C(n_773), .D(n_778), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_776), .B(n_778), .Y(n_816) );
AND2x4_ASAP7_75t_L g817 ( .A(n_763), .B(n_742), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_741), .A2(n_748), .B1(n_773), .B2(n_742), .Y(n_818) );
OAI22xp33_ASAP7_75t_L g819 ( .A1(n_772), .A2(n_785), .B1(n_788), .B2(n_774), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_750), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_741), .B(n_748), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_782), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_755), .B(n_756), .Y(n_823) );
INVx1_ASAP7_75t_SL g824 ( .A(n_784), .Y(n_824) );
NOR2x1p5_ASAP7_75t_L g825 ( .A(n_772), .B(n_785), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_776), .B(n_745), .Y(n_826) );
AND2x4_ASAP7_75t_SL g827 ( .A(n_749), .B(n_785), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_821), .B(n_743), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_807), .A2(n_772), .B1(n_753), .B2(n_749), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_798), .Y(n_830) );
OAI21xp33_ASAP7_75t_L g831 ( .A1(n_818), .A2(n_768), .B(n_762), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_825), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_801), .Y(n_833) );
INVx1_ASAP7_75t_SL g834 ( .A(n_799), .Y(n_834) );
INVxp67_ASAP7_75t_L g835 ( .A(n_799), .Y(n_835) );
AOI211xp5_ASAP7_75t_L g836 ( .A1(n_796), .A2(n_786), .B(n_737), .C(n_787), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_807), .A2(n_810), .B1(n_794), .B2(n_813), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_790), .Y(n_838) );
XOR2x2_ASAP7_75t_L g839 ( .A(n_811), .B(n_759), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_806), .A2(n_754), .B(n_747), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_809), .Y(n_841) );
NOR2x1_ASAP7_75t_L g842 ( .A(n_815), .B(n_779), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_820), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_816), .Y(n_844) );
OAI31xp33_ASAP7_75t_L g845 ( .A1(n_813), .A2(n_756), .A3(n_746), .B(n_755), .Y(n_845) );
INVxp67_ASAP7_75t_L g846 ( .A(n_824), .Y(n_846) );
OAI21xp33_ASAP7_75t_SL g847 ( .A1(n_815), .A2(n_759), .B(n_757), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_816), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_803), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_832), .B(n_810), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_844), .B(n_823), .Y(n_851) );
INVxp67_ASAP7_75t_L g852 ( .A(n_834), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_835), .Y(n_853) );
NAND2xp33_ASAP7_75t_SL g854 ( .A(n_837), .B(n_806), .Y(n_854) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_835), .Y(n_855) );
NAND3xp33_ASAP7_75t_L g856 ( .A(n_847), .B(n_793), .C(n_819), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_846), .Y(n_857) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_839), .A2(n_817), .B1(n_824), .B2(n_804), .Y(n_858) );
OAI32xp33_ASAP7_75t_L g859 ( .A1(n_832), .A2(n_800), .A3(n_792), .B1(n_791), .B2(n_826), .Y(n_859) );
NOR2xp67_ASAP7_75t_L g860 ( .A(n_829), .B(n_817), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_848), .B(n_826), .Y(n_861) );
O2A1O1Ixp33_ASAP7_75t_L g862 ( .A1(n_852), .A2(n_846), .B(n_845), .C(n_836), .Y(n_862) );
NOR2xp33_ASAP7_75t_L g863 ( .A(n_858), .B(n_831), .Y(n_863) );
OR2x2_ASAP7_75t_L g864 ( .A(n_853), .B(n_849), .Y(n_864) );
OR2x2_ASAP7_75t_L g865 ( .A(n_857), .B(n_828), .Y(n_865) );
OR2x2_ASAP7_75t_L g866 ( .A(n_855), .B(n_838), .Y(n_866) );
NOR3xp33_ASAP7_75t_L g867 ( .A(n_854), .B(n_842), .C(n_840), .Y(n_867) );
AOI21xp5_ASAP7_75t_L g868 ( .A1(n_862), .A2(n_852), .B(n_856), .Y(n_868) );
AOI22x1_ASAP7_75t_SL g869 ( .A1(n_867), .A2(n_860), .B1(n_859), .B2(n_833), .Y(n_869) );
NOR3x1_ASAP7_75t_L g870 ( .A(n_865), .B(n_861), .C(n_851), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g871 ( .A1(n_863), .A2(n_850), .B(n_827), .Y(n_871) );
INVx2_ASAP7_75t_L g872 ( .A(n_870), .Y(n_872) );
AOI221x1_ASAP7_75t_L g873 ( .A1(n_868), .A2(n_830), .B1(n_843), .B2(n_841), .C(n_805), .Y(n_873) );
NAND2xp33_ASAP7_75t_R g874 ( .A(n_869), .B(n_866), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_872), .B(n_871), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_873), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g877 ( .A(n_875), .B(n_874), .C(n_864), .D(n_805), .Y(n_877) );
O2A1O1Ixp33_ASAP7_75t_L g878 ( .A1(n_876), .A2(n_814), .B(n_789), .C(n_812), .Y(n_878) );
INVx1_ASAP7_75t_SL g879 ( .A(n_877), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_879), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_880), .A2(n_878), .B1(n_757), .B2(n_758), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_881), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g883 ( .A1(n_882), .A2(n_758), .B1(n_787), .B2(n_808), .Y(n_883) );
NAND3xp33_ASAP7_75t_L g884 ( .A(n_883), .B(n_797), .C(n_822), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_884), .A2(n_738), .B1(n_752), .B2(n_740), .Y(n_885) );
OR2x6_ASAP7_75t_L g886 ( .A(n_885), .B(n_795), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_886), .A2(n_752), .B1(n_770), .B2(n_802), .Y(n_887) );
endmodule