module real_jpeg_30823_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_0),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_1),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_1),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_1),
.B(n_124),
.Y(n_316)
);

OAI32xp33_ASAP7_75t_L g342 ( 
.A1(n_1),
.A2(n_343),
.A3(n_348),
.B1(n_350),
.B2(n_355),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_1),
.A2(n_281),
.B1(n_374),
.B2(n_377),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_1),
.A2(n_223),
.B(n_410),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_108),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_2),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_2),
.A2(n_112),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_2),
.A2(n_112),
.B1(n_286),
.B2(n_290),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_2),
.A2(n_112),
.B1(n_333),
.B2(n_337),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_3),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_4),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_4),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_4),
.A2(n_119),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_4),
.A2(n_119),
.B1(n_359),
.B2(n_362),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_4),
.A2(n_119),
.B1(n_310),
.B2(n_455),
.Y(n_454)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_7),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_7),
.A2(n_157),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_7),
.A2(n_157),
.B1(n_366),
.B2(n_370),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_7),
.A2(n_157),
.B1(n_402),
.B2(n_406),
.Y(n_401)
);

AOI22x1_ASAP7_75t_L g204 ( 
.A1(n_8),
.A2(n_205),
.B1(n_210),
.B2(n_211),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_8),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_8),
.A2(n_210),
.B1(n_230),
.B2(n_233),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_8),
.A2(n_210),
.B1(n_310),
.B2(n_312),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_9),
.A2(n_214),
.B1(n_217),
.B2(n_219),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_9),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_9),
.A2(n_219),
.B1(n_370),
.B2(n_509),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_10),
.A2(n_184),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_10),
.Y(n_257)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_11),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_12),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_12),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_12),
.A2(n_40),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_12),
.A2(n_40),
.B1(n_521),
.B2(n_525),
.Y(n_520)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_14),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_14),
.Y(n_200)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_14),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_15),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_15),
.A2(n_49),
.B1(n_247),
.B2(n_250),
.Y(n_246)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_16),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_491),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_317),
.B(n_485),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_260),
.B(n_295),
.Y(n_20)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_21),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_167),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_22),
.B(n_242),
.C(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_86),
.C(n_125),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_23),
.A2(n_24),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp67_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_57),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_25),
.B(n_57),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_45),
.B2(n_48),
.Y(n_25)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_26),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_26),
.B(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_26),
.A2(n_470),
.B1(n_471),
.B2(n_472),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_28),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_29),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_29),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_29),
.Y(n_216)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_29),
.Y(n_458)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_32),
.Y(n_259)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_32),
.Y(n_412)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_34),
.A2(n_223),
.B1(n_309),
.B2(n_314),
.Y(n_308)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_39),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_39),
.Y(n_336)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_43),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_44),
.Y(n_340)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_44),
.Y(n_409)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_48),
.Y(n_222)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_53),
.Y(n_313)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_56),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_64),
.B1(n_73),
.B2(n_78),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_63),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_66),
.Y(n_91)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_72),
.Y(n_240)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_73),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_86),
.A2(n_87),
.B1(n_125),
.B2(n_126),
.Y(n_264)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_117),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_107),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_89),
.A2(n_118),
.B1(n_124),
.B2(n_236),
.Y(n_235)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_89),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_89),
.B(n_236),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_100),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_94),
.Y(n_347)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_94),
.Y(n_524)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_97),
.Y(n_379)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_99),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_SL g123 ( 
.A(n_104),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_107),
.B(n_124),
.Y(n_277)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_114),
.Y(n_237)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_116),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_153),
.B(n_160),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_127),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_127),
.A2(n_160),
.B(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_128),
.A2(n_269),
.B1(n_274),
.B2(n_275),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_SL g307 ( 
.A(n_128),
.B(n_162),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_128),
.A2(n_161),
.B1(n_229),
.B2(n_520),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_134),
.B1(n_137),
.B2(n_139),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_137),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_138),
.Y(n_193)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_138),
.Y(n_512)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B(n_149),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_145),
.Y(n_232)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_148),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_156),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_161),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g226 ( 
.A(n_162),
.Y(n_226)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_166),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_241),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_168),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_224),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_170),
.B(n_235),
.C(n_498),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_212),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_171),
.B(n_212),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_185),
.B1(n_194),
.B2(n_204),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_172),
.A2(n_185),
.B1(n_194),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_172),
.A2(n_194),
.B1(n_358),
.B2(n_365),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_172),
.B(n_281),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_172),
.A2(n_194),
.B1(n_246),
.B2(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_173),
.A2(n_284),
.B1(n_285),
.B2(n_292),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_173),
.B(n_285),
.Y(n_383)
);

AO22x2_ASAP7_75t_SL g397 ( 
.A1(n_173),
.A2(n_285),
.B1(n_292),
.B2(n_398),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_195),
.Y(n_194)
);

OAI22x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_178),
.B1(n_180),
.B2(n_183),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_175),
.A2(n_196),
.B1(n_199),
.B2(n_201),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_177),
.Y(n_437)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_193),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_194),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_SL g382 ( 
.A1(n_194),
.A2(n_365),
.B(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_197),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_198),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_203),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_203),
.Y(n_429)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_209),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_213),
.A2(n_223),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_220),
.Y(n_471)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_SL g314 ( 
.A(n_221),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_223),
.A2(n_401),
.B(n_410),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_223),
.A2(n_255),
.B(n_504),
.Y(n_503)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_225),
.Y(n_498)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_227),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_SL g305 ( 
.A1(n_227),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g399 ( 
.A(n_227),
.B(n_281),
.Y(n_399)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx4f_ASAP7_75t_SL g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_253),
.B2(n_254),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_245),
.B(n_254),
.Y(n_515)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_250),
.Y(n_441)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_252),
.Y(n_369)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_261),
.B(n_487),
.C(n_490),
.Y(n_486)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.C(n_293),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_262),
.A2(n_263),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_266),
.A2(n_267),
.B1(n_293),
.B2(n_294),
.Y(n_297)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_276),
.C(n_283),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_268),
.B(n_283),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx4f_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_301),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_277),
.B(n_518),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_281),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_281),
.B(n_429),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_281),
.B(n_428),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_281),
.B(n_467),
.Y(n_466)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI211xp5_ASAP7_75t_L g439 ( 
.A1(n_292),
.A2(n_440),
.B(n_441),
.C(n_442),
.Y(n_439)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_296),
.Y(n_489)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_299),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_303),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_300),
.B(n_481),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_302),
.Y(n_482)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.C(n_315),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_305),
.B(n_388),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_308),
.A2(n_315),
.B1(n_316),
.B2(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI21x1_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_476),
.B(n_483),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_390),
.B(n_475),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_380),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_321),
.B(n_380),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_357),
.C(n_372),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_323),
.B(n_394),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_341),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_324),
.B(n_342),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_331),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_330),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_329),
.Y(n_462)
);

OAI21xp33_ASAP7_75t_L g453 ( 
.A1(n_331),
.A2(n_454),
.B(n_459),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_L g410 ( 
.A(n_332),
.B(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_348),
.Y(n_356)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_357),
.B(n_372),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_358),
.Y(n_398)
);

BUFx4f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_387),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_382),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_383),
.B(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_384),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_384),
.B(n_385),
.C(n_479),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_387),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_413),
.B(n_445),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_392),
.B(n_446),
.C(n_449),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.Y(n_392)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_393),
.Y(n_415)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_399),
.C(n_400),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2x1_ASAP7_75t_L g444 ( 
.A(n_397),
.B(n_399),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_444),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g472 ( 
.A(n_401),
.Y(n_472)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx2_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_406),
.B(n_419),
.Y(n_418)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_406),
.Y(n_430)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_416),
.B2(n_443),
.Y(n_413)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_438),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_417),
.B(n_438),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_426),
.B1(n_430),
.B2(n_431),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_428),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_443),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_469),
.C(n_473),
.Y(n_449)
);

OA21x2_ASAP7_75t_SL g450 ( 
.A1(n_451),
.A2(n_463),
.B(n_468),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_452),
.B(n_453),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_454),
.Y(n_470)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_456),
.B(n_466),
.Y(n_465)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_460),
.Y(n_467)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_480),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_480),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_529),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_494),
.B(n_496),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_499),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_514),
.B2(n_528),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_501),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_503),
.B1(n_507),
.B2(n_513),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

BUFx4f_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_507),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_514),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_519),
.Y(n_516)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVxp33_ASAP7_75t_SL g529 ( 
.A(n_530),
.Y(n_529)
);


endmodule