module fake_jpeg_18939_n_327 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_327);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_18),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_26),
.B1(n_21),
.B2(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_20),
.B1(n_41),
.B2(n_43),
.Y(n_64)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_56),
.B(n_18),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_64),
.A2(n_85),
.B1(n_49),
.B2(n_59),
.Y(n_104)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_73),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_62),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_60),
.B(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_42),
.B1(n_43),
.B2(n_26),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_77),
.A2(n_52),
.B1(n_45),
.B2(n_38),
.Y(n_109)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_78),
.Y(n_98)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_25),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_26),
.B1(n_21),
.B2(n_34),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_91),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_43),
.B1(n_44),
.B2(n_37),
.Y(n_85)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_20),
.B1(n_38),
.B2(n_36),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g124 ( 
.A1(n_87),
.A2(n_45),
.B1(n_36),
.B2(n_38),
.Y(n_124)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_66),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_38),
.C(n_36),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_38),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_49),
.B1(n_21),
.B2(n_20),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_104),
.B1(n_78),
.B2(n_94),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_35),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_100),
.A2(n_113),
.B(n_120),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_85),
.B(n_77),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_124),
.B1(n_65),
.B2(n_88),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_72),
.B1(n_75),
.B2(n_92),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_69),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_112),
.B(n_118),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_SL g120 ( 
.A1(n_83),
.A2(n_87),
.B(n_80),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_76),
.B(n_27),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_129),
.Y(n_163)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_63),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_105),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_66),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_136),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_38),
.C(n_36),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_133),
.B(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_86),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_140),
.A2(n_96),
.B1(n_90),
.B2(n_18),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_68),
.B1(n_35),
.B2(n_44),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_147),
.B1(n_154),
.B2(n_98),
.Y(n_160)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_37),
.B(n_44),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_152),
.B(n_147),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_108),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_35),
.B1(n_37),
.B2(n_22),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_101),
.A2(n_34),
.B1(n_27),
.B2(n_30),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_28),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2x1p5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_53),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_86),
.C(n_24),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_98),
.A2(n_30),
.B1(n_13),
.B2(n_14),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_164),
.B1(n_172),
.B2(n_175),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_170),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_114),
.B1(n_107),
.B2(n_103),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_143),
.B(n_132),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_165),
.A2(n_169),
.B(n_143),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_168),
.B1(n_176),
.B2(n_187),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_103),
.B1(n_114),
.B2(n_107),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_131),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_178),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_125),
.B1(n_108),
.B2(n_115),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_153),
.A2(n_115),
.B1(n_105),
.B2(n_123),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_12),
.B1(n_14),
.B2(n_11),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_183),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_135),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_18),
.B1(n_24),
.B2(n_25),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_154),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_127),
.A2(n_31),
.B1(n_29),
.B2(n_19),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_140),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_188)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_129),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_189)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_172),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_165),
.A2(n_136),
.B(n_148),
.Y(n_193)
);

AOI211xp5_ASAP7_75t_L g236 ( 
.A1(n_193),
.A2(n_187),
.B(n_175),
.C(n_160),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_151),
.C(n_141),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_204),
.C(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_161),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_206),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_167),
.B1(n_168),
.B2(n_158),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_139),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_202),
.B(n_203),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_28),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_138),
.C(n_25),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_161),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_28),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

AOI21x1_ASAP7_75t_SL g208 ( 
.A1(n_169),
.A2(n_17),
.B(n_1),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_5),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_218),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_159),
.B(n_6),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_211),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_214),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_178),
.B(n_6),
.C(n_9),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_181),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_176),
.B(n_6),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_11),
.C(n_4),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_218),
.C(n_209),
.Y(n_239)
);

BUFx12f_ASAP7_75t_SL g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2x1_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_234),
.Y(n_259)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_225),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_230),
.B(n_237),
.Y(n_245)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_189),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_198),
.A2(n_164),
.B1(n_158),
.B2(n_181),
.Y(n_238)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_182),
.B1(n_166),
.B2(n_157),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_241),
.A2(n_243),
.B1(n_213),
.B2(n_212),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_190),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_247),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_196),
.B1(n_192),
.B2(n_217),
.Y(n_252)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_203),
.C(n_192),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_257),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_199),
.B1(n_208),
.B2(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_215),
.C(n_219),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_240),
.B(n_221),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_188),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_182),
.C(n_171),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_263),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_157),
.C(n_210),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_265),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_256),
.B(n_230),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_266),
.A2(n_271),
.B(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_222),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_245),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_246),
.B(n_221),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_275),
.A2(n_261),
.B(n_233),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_263),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_276),
.Y(n_289)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_262),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_247),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_272),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_282),
.B(n_288),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_280),
.B1(n_267),
.B2(n_252),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_290),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_245),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_253),
.C(n_255),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_244),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_280),
.C(n_270),
.Y(n_304)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_273),
.Y(n_293)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_293),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g294 ( 
.A1(n_265),
.A2(n_257),
.B1(n_239),
.B2(n_235),
.C(n_260),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_235),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_270),
.C(n_275),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_293),
.Y(n_297)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_303),
.B(n_4),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_271),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_4),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_287),
.B(n_283),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_7),
.B(n_8),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_266),
.B1(n_291),
.B2(n_282),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_296),
.B1(n_299),
.B2(n_156),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_8),
.B1(n_9),
.B2(n_2),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_7),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_311),
.B(n_299),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_315),
.A2(n_316),
.B(n_318),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_309),
.B(n_308),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_307),
.B(n_312),
.Y(n_320)
);

A2O1A1O1Ixp25_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_321),
.B(n_8),
.C(n_3),
.D(n_1),
.Y(n_323)
);

AO22x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_0),
.C(n_1),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_0),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_3),
.B(n_273),
.Y(n_327)
);


endmodule