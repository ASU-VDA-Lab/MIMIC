module real_aes_10116_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_87;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_649;
wire n_193;
wire n_162;
wire n_293;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_639;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
NAND2xp5_ASAP7_75t_L g151 ( .A(n_0), .B(n_152), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_1), .A2(n_66), .B1(n_150), .B2(n_202), .Y(n_201) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_2), .Y(n_596) );
INVx1_ASAP7_75t_L g632 ( .A(n_2), .Y(n_632) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_3), .Y(n_156) );
INVx1_ASAP7_75t_L g578 ( .A(n_4), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_4), .A2(n_58), .B1(n_652), .B2(n_654), .Y(n_651) );
INVx2_ASAP7_75t_L g496 ( .A(n_5), .Y(n_496) );
BUFx2_ASAP7_75t_L g544 ( .A(n_6), .Y(n_544) );
BUFx2_ASAP7_75t_L g593 ( .A(n_6), .Y(n_593) );
INVx1_ASAP7_75t_L g630 ( .A(n_6), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_7), .A2(n_30), .B1(n_170), .B2(n_171), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_8), .A2(n_47), .B1(n_171), .B2(n_173), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_9), .B(n_139), .C(n_171), .Y(n_195) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_9), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_10), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_11), .A2(n_76), .B1(n_612), .B2(n_613), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_11), .A2(n_76), .B1(n_639), .B2(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g504 ( .A(n_12), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_12), .A2(n_41), .B1(n_617), .B2(n_620), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_13), .B(n_117), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_14), .B(n_89), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g190 ( .A(n_15), .B(n_93), .C(n_142), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_16), .A2(n_20), .B1(n_142), .B2(n_170), .Y(n_200) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_16), .Y(n_706) );
INVx1_ASAP7_75t_L g521 ( .A(n_17), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_17), .A2(n_34), .B1(n_622), .B2(n_626), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_18), .B(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
HB1xp67_ASAP7_75t_L g715 ( .A(n_20), .Y(n_715) );
BUFx6f_ASAP7_75t_L g90 ( .A(n_21), .Y(n_90) );
INVx1_ASAP7_75t_L g678 ( .A(n_22), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_23), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_24), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g542 ( .A(n_25), .Y(n_542) );
INVx1_ASAP7_75t_L g704 ( .A(n_25), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_26), .A2(n_38), .B1(n_173), .B2(n_176), .Y(n_172) );
XNOR2xp5_ASAP7_75t_L g487 ( .A(n_27), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_28), .B(n_93), .Y(n_188) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_29), .A2(n_51), .B(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g217 ( .A(n_31), .B(n_128), .Y(n_217) );
AND2x6_ASAP7_75t_L g83 ( .A(n_32), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_32), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_32), .B(n_662), .Y(n_719) );
NAND2x1p5_ASAP7_75t_L g196 ( .A(n_33), .B(n_128), .Y(n_196) );
INVx1_ASAP7_75t_L g492 ( .A(n_34), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_35), .B(n_89), .Y(n_121) );
INVx1_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_36), .Y(n_662) );
INVx1_ASAP7_75t_L g555 ( .A(n_37), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_37), .A2(n_63), .B1(n_646), .B2(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_39), .B(n_128), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_40), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g515 ( .A(n_41), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_42), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_43), .A2(n_53), .B1(n_604), .B2(n_608), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_43), .A2(n_53), .B1(n_644), .B2(n_646), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_44), .B(n_142), .Y(n_230) );
NAND2x1_ASAP7_75t_L g127 ( .A(n_45), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_46), .B(n_139), .Y(n_149) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_48), .Y(n_674) );
INVx2_ASAP7_75t_L g554 ( .A(n_49), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_50), .B(n_224), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_52), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_54), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g525 ( .A(n_55), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_55), .A2(n_67), .B1(n_562), .B2(n_567), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_56), .A2(n_60), .B1(n_142), .B2(n_170), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_57), .Y(n_160) );
INVx1_ASAP7_75t_L g583 ( .A(n_58), .Y(n_583) );
BUFx10_ASAP7_75t_L g698 ( .A(n_59), .Y(n_698) );
INVx1_ASAP7_75t_SL g205 ( .A(n_61), .Y(n_205) );
INVx2_ASAP7_75t_L g560 ( .A(n_62), .Y(n_560) );
INVx1_ASAP7_75t_L g565 ( .A(n_62), .Y(n_565) );
INVx1_ASAP7_75t_L g589 ( .A(n_63), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_64), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_65), .Y(n_125) );
INVx1_ASAP7_75t_L g532 ( .A(n_67), .Y(n_532) );
INVx2_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_69), .B(n_139), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_70), .B(n_114), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_71), .Y(n_671) );
INVx2_ASAP7_75t_L g552 ( .A(n_72), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_73), .B(n_118), .Y(n_228) );
BUFx3_ASAP7_75t_L g501 ( .A(n_74), .Y(n_501) );
INVx1_ASAP7_75t_L g519 ( .A(n_74), .Y(n_519) );
BUFx3_ASAP7_75t_L g503 ( .A(n_75), .Y(n_503) );
INVx1_ASAP7_75t_L g509 ( .A(n_75), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_486), .Y(n_77) );
BUFx3_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_81), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_82), .A2(n_151), .B(n_162), .Y(n_161) );
INVx8_ASAP7_75t_L g166 ( .A(n_82), .Y(n_166) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx2_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_83), .A2(n_134), .B(n_137), .Y(n_133) );
OAI21x1_ASAP7_75t_L g186 ( .A1(n_83), .A2(n_187), .B(n_191), .Y(n_186) );
INVx1_ASAP7_75t_L g234 ( .A(n_83), .Y(n_234) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g717 ( .A1(n_86), .A2(n_718), .B(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_91), .Y(n_86) );
HB1xp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx1_ASAP7_75t_L g123 ( .A(n_89), .Y(n_123) );
INVx2_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx2_ASAP7_75t_L g158 ( .A(n_89), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_89), .B(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_90), .Y(n_118) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_90), .Y(n_171) );
INVx1_ASAP7_75t_L g175 ( .A(n_90), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_91), .A2(n_169), .B1(n_172), .B2(n_177), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_92), .Y(n_91) );
AOI21x1_ASAP7_75t_L g120 ( .A1(n_92), .A2(n_121), .B(n_122), .Y(n_120) );
INVx3_ASAP7_75t_L g203 ( .A(n_92), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_92), .A2(n_230), .B(n_231), .Y(n_229) );
BUFx12f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx5_ASAP7_75t_L g119 ( .A(n_93), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_93), .A2(n_138), .B1(n_140), .B2(n_141), .Y(n_137) );
INVx5_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
OAI321xp33_ASAP7_75t_L g147 ( .A1(n_93), .A2(n_142), .A3(n_148), .B1(n_149), .B2(n_150), .C(n_151), .Y(n_147) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NOR3x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_363), .C(n_458), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_306), .Y(n_96) );
NAND3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_252), .C(n_285), .Y(n_97) );
AOI221xp5_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_181), .B1(n_206), .B2(n_235), .C(n_239), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_144), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_101), .B(n_362), .Y(n_419) );
INVx2_ASAP7_75t_SL g430 ( .A(n_101), .Y(n_430) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_130), .Y(n_101) );
INVx1_ASAP7_75t_L g288 ( .A(n_102), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_102), .B(n_130), .Y(n_338) );
AND2x2_ASAP7_75t_L g432 ( .A(n_102), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_L g335 ( .A(n_103), .B(n_163), .Y(n_335) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_103), .Y(n_358) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g256 ( .A(n_104), .Y(n_256) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_111), .B(n_127), .Y(n_104) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_105), .A2(n_133), .B(n_143), .Y(n_132) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_105), .A2(n_111), .B(n_127), .Y(n_246) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_105), .A2(n_133), .B(n_143), .Y(n_269) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AO31x2_ASAP7_75t_L g198 ( .A1(n_106), .A2(n_166), .A3(n_199), .B(n_204), .Y(n_198) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g167 ( .A(n_107), .Y(n_167) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_107), .Y(n_275) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g129 ( .A(n_108), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_108), .B(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_120), .B(n_126), .Y(n_111) );
AOI21x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_119), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g176 ( .A(n_115), .Y(n_176) );
INVxp67_ASAP7_75t_L g189 ( .A(n_117), .Y(n_189) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g170 ( .A(n_118), .Y(n_170) );
INVx2_ASAP7_75t_L g232 ( .A(n_118), .Y(n_232) );
AOI21x1_ASAP7_75t_L g134 ( .A1(n_119), .A2(n_135), .B(n_136), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_119), .A2(n_154), .B(n_159), .Y(n_153) );
CKINVDCx6p67_ASAP7_75t_R g177 ( .A(n_119), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g324 ( .A(n_131), .Y(n_324) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g320 ( .A(n_132), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_139), .A2(n_142), .B(n_227), .C(n_228), .Y(n_226) );
INVx2_ASAP7_75t_SL g194 ( .A(n_142), .Y(n_194) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g283 ( .A(n_145), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g304 ( .A(n_145), .B(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g327 ( .A(n_145), .Y(n_327) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_163), .Y(n_145) );
INVx2_ASAP7_75t_L g238 ( .A(n_146), .Y(n_238) );
INVx1_ASAP7_75t_L g248 ( .A(n_146), .Y(n_248) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B(n_161), .Y(n_146) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx1_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
BUFx5_ASAP7_75t_L g212 ( .A(n_152), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g258 ( .A(n_163), .Y(n_258) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g237 ( .A(n_164), .Y(n_237) );
AOI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_178), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g202 ( .A(n_175), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_177), .A2(n_200), .B1(n_201), .B2(n_203), .Y(n_199) );
OA22x2_ASAP7_75t_L g213 ( .A1(n_177), .A2(n_203), .B1(n_214), .B2(n_215), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_180), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g224 ( .A(n_180), .Y(n_224) );
INVxp67_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_197), .Y(n_182) );
INVx2_ASAP7_75t_L g301 ( .A(n_183), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_183), .B(n_410), .Y(n_409) );
NAND2xp33_ASAP7_75t_SL g452 ( .A(n_183), .B(n_376), .Y(n_452) );
BUFx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g220 ( .A(n_184), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g295 ( .A(n_184), .B(n_222), .Y(n_295) );
OAI21x1_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_196), .Y(n_184) );
OAI21x1_ASAP7_75t_L g263 ( .A1(n_185), .A2(n_186), .B(n_196), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_190), .Y(n_187) );
OAI21xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2x1_ASAP7_75t_L g218 ( .A(n_197), .B(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g442 ( .A(n_197), .Y(n_442) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_197), .Y(n_466) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g264 ( .A(n_198), .Y(n_264) );
INVx1_ASAP7_75t_L g292 ( .A(n_198), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_198), .B(n_274), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_198), .B(n_209), .Y(n_377) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_198), .Y(n_456) );
OAI22xp33_ASAP7_75t_SL g460 ( .A1(n_206), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_460) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_218), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_207), .B(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g329 ( .A(n_207), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g440 ( .A(n_207), .Y(n_440) );
AND2x2_ASAP7_75t_L g485 ( .A(n_207), .B(n_339), .Y(n_485) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g348 ( .A(n_208), .B(n_339), .Y(n_348) );
AND2x2_ASAP7_75t_L g420 ( .A(n_208), .B(n_421), .Y(n_420) );
NOR2x1_ASAP7_75t_L g434 ( .A(n_208), .B(n_291), .Y(n_434) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
INVx1_ASAP7_75t_L g282 ( .A(n_209), .Y(n_282) );
INVxp67_ASAP7_75t_SL g297 ( .A(n_209), .Y(n_297) );
HB1xp67_ASAP7_75t_L g484 ( .A(n_209), .Y(n_484) );
OAI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_213), .B(n_216), .Y(n_209) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_213), .A2(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVxp67_ASAP7_75t_L g276 ( .A(n_217), .Y(n_276) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g250 ( .A(n_220), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g341 ( .A(n_220), .Y(n_341) );
INVx2_ASAP7_75t_L g273 ( .A(n_221), .Y(n_273) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g281 ( .A(n_222), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_223), .B(n_225), .Y(n_222) );
OAI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_229), .B(n_233), .Y(n_225) );
NAND3xp33_ASAP7_75t_L g439 ( .A(n_235), .B(n_440), .C(n_441), .Y(n_439) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g287 ( .A(n_236), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g317 ( .A(n_236), .B(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_236), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g412 ( .A(n_236), .B(n_244), .Y(n_412) );
OR2x2_ASAP7_75t_L g438 ( .A(n_236), .B(n_338), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_236), .B(n_305), .Y(n_457) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g247 ( .A(n_237), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_237), .B(n_284), .Y(n_345) );
AND2x2_ASAP7_75t_L g267 ( .A(n_238), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g384 ( .A(n_238), .B(n_269), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_247), .Y(n_241) );
OR2x2_ASAP7_75t_L g451 ( .A(n_242), .B(n_345), .Y(n_451) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g388 ( .A(n_243), .B(n_324), .Y(n_388) );
AND2x2_ASAP7_75t_L g424 ( .A(n_243), .B(n_267), .Y(n_424) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g270 ( .A(n_244), .B(n_257), .Y(n_270) );
AND2x2_ASAP7_75t_L g396 ( .A(n_244), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g404 ( .A(n_244), .B(n_331), .Y(n_404) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_244), .Y(n_417) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_258), .Y(n_323) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g370 ( .A(n_246), .B(n_248), .Y(n_370) );
AND2x2_ASAP7_75t_L g333 ( .A(n_247), .B(n_319), .Y(n_333) );
INVx2_ASAP7_75t_L g362 ( .A(n_247), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_247), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g402 ( .A(n_248), .Y(n_402) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g312 ( .A(n_251), .Y(n_312) );
AND2x2_ASAP7_75t_L g475 ( .A(n_251), .B(n_280), .Y(n_475) );
AOI322xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_259), .A3(n_265), .B1(n_270), .B2(n_271), .C1(n_277), .C2(n_283), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_254), .A2(n_479), .B(n_481), .C(n_485), .Y(n_478) );
BUFx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AOI32xp33_ASAP7_75t_L g453 ( .A1(n_255), .A2(n_383), .A3(n_421), .B1(n_454), .B2(n_457), .Y(n_453) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
BUFx2_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_256), .Y(n_326) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_258), .Y(n_369) );
NOR2x1p5_ASAP7_75t_L g379 ( .A(n_260), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g271 ( .A(n_261), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g331 ( .A(n_262), .B(n_273), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_262), .B(n_281), .Y(n_394) );
INVx1_ASAP7_75t_L g433 ( .A(n_262), .Y(n_433) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g355 ( .A(n_263), .B(n_274), .Y(n_355) );
AND2x4_ASAP7_75t_L g280 ( .A(n_264), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g411 ( .A(n_264), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_265), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_266), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g284 ( .A(n_269), .Y(n_284) );
INVx1_ASAP7_75t_L g385 ( .A(n_270), .Y(n_385) );
AND2x4_ASAP7_75t_L g462 ( .A(n_270), .B(n_324), .Y(n_462) );
INVx2_ASAP7_75t_L g386 ( .A(n_272), .Y(n_386) );
AND2x4_ASAP7_75t_L g408 ( .A(n_272), .B(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
AND2x2_ASAP7_75t_L g339 ( .A(n_273), .B(n_292), .Y(n_339) );
INVx2_ASAP7_75t_L g354 ( .A(n_273), .Y(n_354) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_278), .A2(n_406), .B1(n_407), .B2(n_412), .Y(n_405) );
OR2x6_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x4_ASAP7_75t_L g313 ( .A(n_280), .B(n_301), .Y(n_313) );
INVx1_ASAP7_75t_L g389 ( .A(n_280), .Y(n_389) );
AND2x2_ASAP7_75t_L g421 ( .A(n_281), .B(n_411), .Y(n_421) );
AND2x2_ASAP7_75t_L g381 ( .A(n_282), .B(n_354), .Y(n_381) );
AND2x2_ASAP7_75t_L g449 ( .A(n_282), .B(n_295), .Y(n_449) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_283), .Y(n_349) );
INVx2_ASAP7_75t_L g305 ( .A(n_284), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_289), .B1(n_298), .B2(n_302), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_288), .B(n_384), .Y(n_406) );
AOI221xp5_ASAP7_75t_SL g342 ( .A1(n_289), .A2(n_343), .B1(n_346), .B2(n_349), .C(n_350), .Y(n_342) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp67_ASAP7_75t_L g353 ( .A(n_292), .B(n_354), .Y(n_353) );
BUFx2_ASAP7_75t_L g423 ( .A(n_293), .Y(n_423) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_294), .B(n_329), .C(n_347), .Y(n_346) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g375 ( .A(n_295), .Y(n_375) );
AND2x2_ASAP7_75t_L g454 ( .A(n_295), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
AND2x4_ASAP7_75t_L g401 ( .A(n_305), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_342), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_314), .B(n_328), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_310), .B(n_313), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_310), .A2(n_391), .B(n_405), .Y(n_390) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g360 ( .A(n_312), .B(n_331), .Y(n_360) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_321), .C(n_325), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_318), .Y(n_480) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g418 ( .A(n_320), .B(n_402), .Y(n_418) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g463 ( .A(n_322), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g448 ( .A(n_323), .Y(n_448) );
AND2x2_ASAP7_75t_L g365 ( .A(n_324), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g471 ( .A(n_324), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_332), .B(n_336), .Y(n_328) );
INVx2_ASAP7_75t_L g445 ( .A(n_330), .Y(n_445) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_333), .A2(n_337), .B1(n_339), .B2(n_340), .Y(n_336) );
INVx2_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g467 ( .A1(n_335), .A2(n_468), .B1(n_473), .B2(n_476), .C(n_478), .Y(n_467) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g397 ( .A(n_345), .Y(n_397) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_356), .B1(n_359), .B2(n_361), .Y(n_350) );
INVx1_ASAP7_75t_L g461 ( .A(n_351), .Y(n_461) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
AND2x4_ASAP7_75t_L g435 ( .A(n_355), .B(n_421), .Y(n_435) );
OR2x2_ASAP7_75t_L g361 ( .A(n_357), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g367 ( .A(n_359), .Y(n_367) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g465 ( .A(n_360), .B(n_466), .Y(n_465) );
NAND4xp75_ASAP7_75t_L g363 ( .A(n_364), .B(n_390), .C(n_413), .D(n_436), .Y(n_363) );
AOI221x1_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B1(n_368), .B2(n_371), .C(n_382), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_368), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_378), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_376), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_376), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g469 ( .A(n_376), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_377), .B(n_394), .Y(n_472) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OAI32xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_385), .A3(n_386), .B1(n_387), .B2(n_389), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_384), .A2(n_432), .B(n_434), .C(n_435), .Y(n_431) );
AND2x2_ASAP7_75t_L g446 ( .A(n_384), .B(n_447), .Y(n_446) );
OAI22xp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B1(n_398), .B2(n_403), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx4_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_401), .Y(n_477) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_412), .A2(n_451), .B(n_452), .C(n_453), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g413 ( .A(n_414), .B(n_425), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_422), .Y(n_414) );
OAI21xp33_ASAP7_75t_SL g415 ( .A1(n_416), .A2(n_419), .B(n_420), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_431), .Y(n_425) );
NAND2x1_ASAP7_75t_SL g426 ( .A(n_427), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g470 ( .A(n_429), .Y(n_470) );
AND2x2_ASAP7_75t_L g474 ( .A(n_432), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_433), .B(n_484), .Y(n_483) );
AOI221x1_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_443), .B1(n_446), .B2(n_449), .C(n_450), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g482 ( .A(n_442), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_467), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_472), .Y(n_468) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVxp67_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B1(n_660), .B2(n_665), .C(n_711), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_488), .A2(n_712), .B1(n_715), .B2(n_716), .Y(n_711) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI211x1_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_539), .B(n_545), .C(n_597), .Y(n_489) );
NAND4xp25_ASAP7_75t_SL g490 ( .A(n_491), .B(n_510), .C(n_520), .D(n_535), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B1(n_504), .B2(n_505), .Y(n_491) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
AND2x6_ASAP7_75t_L g516 ( .A(n_494), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g507 ( .A(n_496), .Y(n_507) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_496), .Y(n_514) );
AND2x2_ASAP7_75t_L g637 ( .A(n_496), .B(n_542), .Y(n_637) );
INVx2_ASAP7_75t_L g659 ( .A(n_496), .Y(n_659) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g645 ( .A(n_498), .Y(n_645) );
INVx6_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g512 ( .A(n_499), .B(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g650 ( .A(n_499), .Y(n_650) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g534 ( .A(n_500), .Y(n_534) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g508 ( .A(n_501), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g524 ( .A(n_501), .B(n_503), .Y(n_524) );
INVx1_ASAP7_75t_L g531 ( .A(n_502), .Y(n_531) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x4_ASAP7_75t_L g518 ( .A(n_503), .B(n_519), .Y(n_518) );
AND2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g537 ( .A(n_506), .Y(n_537) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x6_ASAP7_75t_L g533 ( .A(n_507), .B(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_508), .Y(n_640) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_508), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_515), .B2(n_516), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_511), .A2(n_585), .B1(n_589), .B2(n_590), .Y(n_584) );
AND2x4_ASAP7_75t_L g528 ( .A(n_513), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g642 ( .A(n_517), .Y(n_642) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g655 ( .A(n_518), .Y(n_655) );
AOI222xp33_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_525), .B2(n_526), .C1(n_532), .C2(n_533), .Y(n_520) );
BUFx4f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_SL g647 ( .A(n_523), .Y(n_647) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_524), .Y(n_538) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g696 ( .A(n_531), .Y(n_696) );
INVx5_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x4_ASAP7_75t_L g658 ( .A(n_542), .B(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g601 ( .A(n_544), .Y(n_601) );
AOI31xp33_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_570), .A3(n_584), .B(n_592), .Y(n_545) );
AOI211xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_555), .B(n_556), .C(n_561), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g556 ( .A(n_550), .B(n_557), .Y(n_556) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_550), .Y(n_610) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g569 ( .A(n_552), .Y(n_569) );
INVx2_ASAP7_75t_L g575 ( .A(n_552), .Y(n_575) );
AND2x4_ASAP7_75t_L g582 ( .A(n_552), .B(n_553), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_552), .B(n_554), .Y(n_588) );
AND2x2_ASAP7_75t_L g607 ( .A(n_552), .B(n_554), .Y(n_607) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g566 ( .A(n_554), .Y(n_566) );
INVx1_ASAP7_75t_L g577 ( .A(n_554), .Y(n_577) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g631 ( .A(n_559), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g573 ( .A(n_560), .Y(n_573) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_566), .Y(n_563) );
OR2x6_ASAP7_75t_L g586 ( .A(n_564), .B(n_587), .Y(n_586) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g567 ( .A(n_565), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g602 ( .A(n_565), .B(n_595), .Y(n_602) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_578), .B1(n_579), .B2(n_583), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
AND2x4_ASAP7_75t_L g579 ( .A(n_572), .B(n_580), .Y(n_579) );
OR2x6_ASAP7_75t_L g591 ( .A(n_572), .B(n_587), .Y(n_591) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g612 ( .A(n_574), .Y(n_612) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_574), .Y(n_619) );
AND2x4_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_582), .Y(n_615) );
INVx8_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx4_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x6_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x4_ASAP7_75t_L g657 ( .A(n_593), .B(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_633), .Y(n_597) );
AOI33xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_603), .A3(n_611), .B1(n_616), .B2(n_621), .B3(n_627), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
OR2x6_ASAP7_75t_L g635 ( .A(n_601), .B(n_636), .Y(n_635) );
BUFx3_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_607), .Y(n_625) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g626 ( .A(n_609), .Y(n_626) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
INVx4_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx3_ASAP7_75t_L g620 ( .A(n_615), .Y(n_620) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx6_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x6_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AOI33xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_638), .A3(n_643), .B1(n_648), .B2(n_651), .B3(n_656), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g692 ( .A(n_637), .Y(n_692) );
BUFx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx3_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx4f_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AND2x4_ASAP7_75t_L g702 ( .A(n_659), .B(n_703), .Y(n_702) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_662), .B(n_664), .Y(n_688) );
INVx1_ASAP7_75t_SL g718 ( .A(n_662), .Y(n_718) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_684), .B1(n_706), .B2(n_707), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_666), .A2(n_706), .B1(n_713), .B2(n_714), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_672), .B1(n_682), .B2(n_683), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_667), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_672), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B1(n_676), .B2(n_681), .Y(n_672) );
CKINVDCx14_ASAP7_75t_R g681 ( .A(n_673), .Y(n_681) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_679), .B2(n_680), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_679), .Y(n_680) );
INVx8_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx8_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_687), .Y(n_713) );
OR2x6_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OR2x4_ASAP7_75t_L g710 ( .A(n_688), .B(n_690), .Y(n_710) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AOI31xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .A3(n_697), .B(n_699), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g705 ( .A(n_696), .Y(n_705) );
INVx6_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx4_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx8_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g714 ( .A(n_709), .Y(n_714) );
INVx8_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx2_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
endmodule