module fake_jpeg_29945_n_471 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_49),
.Y(n_146)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_0),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_52),
.B(n_70),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g102 ( 
.A(n_54),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_56),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_31),
.B(n_8),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_61),
.B(n_65),
.Y(n_124)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_68),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_18),
.B(n_8),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_32),
.B(n_1),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_72),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_76),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_74),
.B(n_84),
.Y(n_123)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_9),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_32),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_90),
.Y(n_139)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_86),
.Y(n_135)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_17),
.Y(n_87)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_89),
.Y(n_128)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_27),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_92),
.B(n_93),
.Y(n_133)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_17),
.Y(n_93)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_20),
.B1(n_17),
.B2(n_44),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_96),
.A2(n_97),
.B1(n_103),
.B2(n_107),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_88),
.B1(n_84),
.B2(n_74),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_20),
.B1(n_17),
.B2(n_44),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_20),
.B1(n_46),
.B2(n_33),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_104),
.A2(n_117),
.B1(n_127),
.B2(n_137),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_44),
.B1(n_43),
.B2(n_27),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_108),
.A2(n_111),
.B1(n_113),
.B2(n_121),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_28),
.B1(n_46),
.B2(n_42),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_49),
.A2(n_26),
.B1(n_47),
.B2(n_39),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_51),
.A2(n_30),
.B1(n_28),
.B2(n_42),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_70),
.A2(n_48),
.B1(n_47),
.B2(n_39),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_70),
.A2(n_48),
.B1(n_39),
.B2(n_38),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_52),
.B(n_30),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_136),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_52),
.B(n_41),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_71),
.A2(n_41),
.B1(n_25),
.B2(n_29),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_85),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_142),
.B1(n_75),
.B2(n_1),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_50),
.A2(n_38),
.B1(n_34),
.B2(n_26),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_81),
.A2(n_35),
.B1(n_38),
.B2(n_34),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_59),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_95),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_183),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

BUFx16f_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_56),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_157),
.Y(n_200)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_55),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_163),
.Y(n_206)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_112),
.A2(n_69),
.B1(n_83),
.B2(n_58),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_160),
.A2(n_172),
.B1(n_191),
.B2(n_135),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_117),
.A2(n_72),
.B1(n_64),
.B2(n_92),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_98),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_166),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_78),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_167),
.B(n_177),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_90),
.B1(n_63),
.B2(n_57),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_170),
.A2(n_135),
.B1(n_99),
.B2(n_126),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_123),
.B(n_26),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_171),
.B(n_193),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_114),
.A2(n_34),
.B1(n_86),
.B2(n_87),
.Y(n_172)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_175),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_102),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_176),
.B(n_189),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_136),
.B(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_180),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_116),
.B(n_62),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_181),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_93),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_35),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_77),
.B(n_94),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_185),
.A2(n_133),
.B(n_135),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_35),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_192),
.Y(n_208)
);

INVx5_ASAP7_75t_SL g187 ( 
.A(n_102),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_188),
.Y(n_231)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_125),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_190),
.Y(n_236)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_94),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_54),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_196),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_130),
.B(n_86),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_195),
.B(n_147),
.Y(n_226)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_86),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_7),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_152),
.B(n_127),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_202),
.B(n_215),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_158),
.B(n_102),
.Y(n_212)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_212),
.B(n_154),
.CI(n_159),
.CON(n_266),
.SN(n_266)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_158),
.B(n_121),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_219),
.B(n_234),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_231),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_163),
.B(n_148),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_197),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_232),
.B(n_237),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_235),
.B1(n_169),
.B2(n_154),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g234 ( 
.A1(n_183),
.A2(n_145),
.B(n_99),
.C(n_132),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_161),
.A2(n_134),
.B1(n_115),
.B2(n_145),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_150),
.B(n_132),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_173),
.A2(n_146),
.B1(n_118),
.B2(n_99),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_238),
.A2(n_185),
.B(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_150),
.B(n_134),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_240),
.B(n_161),
.Y(n_243)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_242),
.B(n_263),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_243),
.B(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_245),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_230),
.Y(n_247)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_247),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_218),
.B(n_186),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_192),
.C(n_194),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_251),
.B(n_209),
.C(n_236),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_199),
.B(n_174),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_252),
.B(n_227),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_228),
.A2(n_171),
.B1(n_184),
.B2(n_151),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_253),
.A2(n_269),
.B1(n_219),
.B2(n_214),
.Y(n_280)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_207),
.Y(n_254)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_254),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_187),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_256),
.Y(n_306)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_213),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_200),
.B(n_176),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_261),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_233),
.B1(n_222),
.B2(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_213),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_206),
.A2(n_175),
.B1(n_181),
.B2(n_196),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_224),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_265),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_267),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_191),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_221),
.B(n_177),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_270),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_228),
.A2(n_206),
.B1(n_214),
.B2(n_238),
.Y(n_269)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_220),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_271),
.Y(n_291)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_206),
.B(n_164),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_222),
.B(n_234),
.Y(n_294)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_276),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_221),
.B(n_188),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_278),
.A2(n_231),
.B1(n_224),
.B2(n_217),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_220),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_281),
.A2(n_282),
.B1(n_290),
.B2(n_304),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_243),
.A2(n_215),
.B1(n_232),
.B2(n_212),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_208),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_288),
.B(n_308),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_262),
.A2(n_214),
.B1(n_212),
.B2(n_235),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_289),
.A2(n_294),
.B(n_302),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_240),
.B1(n_237),
.B2(n_202),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_293),
.B(n_264),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_252),
.A2(n_210),
.B1(n_234),
.B2(n_199),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_297),
.A2(n_274),
.B1(n_248),
.B2(n_267),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_273),
.A2(n_210),
.B(n_226),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_242),
.A2(n_209),
.B1(n_217),
.B2(n_227),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_249),
.A2(n_231),
.B(n_224),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_313),
.B(n_315),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_251),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_249),
.A2(n_224),
.B(n_156),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_266),
.A2(n_190),
.B(n_205),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_317),
.Y(n_353)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_295),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_340),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_299),
.A2(n_266),
.B(n_272),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_320),
.A2(n_309),
.B(n_313),
.Y(n_359)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_321),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_277),
.Y(n_322)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_322),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_323),
.B(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_291),
.B(n_265),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_336),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g372 ( 
.A1(n_328),
.A2(n_310),
.B(n_306),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_299),
.A2(n_279),
.B1(n_273),
.B2(n_271),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_329),
.A2(n_337),
.B1(n_349),
.B2(n_294),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_308),
.B(n_272),
.C(n_263),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_332),
.C(n_282),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_268),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_289),
.A2(n_301),
.B1(n_280),
.B2(n_297),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_333),
.A2(n_290),
.B1(n_304),
.B2(n_281),
.Y(n_356)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_285),
.Y(n_335)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_264),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_299),
.A2(n_260),
.B1(n_241),
.B2(n_244),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_291),
.B(n_245),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_339),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_247),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_284),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_278),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_343),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_300),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_342),
.B(n_344),
.Y(n_368)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_286),
.B(n_312),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_284),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_346),
.B(n_347),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_275),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_298),
.B(n_250),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_292),
.B1(n_310),
.B2(n_306),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_299),
.A2(n_256),
.B1(n_261),
.B2(n_258),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_327),
.B1(n_337),
.B2(n_329),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_308),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_352),
.B(n_354),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_301),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_361),
.C(n_378),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_356),
.A2(n_365),
.B1(n_371),
.B2(n_375),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_359),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_331),
.B(n_288),
.C(n_289),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_345),
.A2(n_315),
.B(n_312),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_340),
.Y(n_363)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_334),
.A2(n_288),
.B1(n_316),
.B2(n_287),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_338),
.Y(n_383)
);

AOI21x1_ASAP7_75t_L g370 ( 
.A1(n_325),
.A2(n_302),
.B(n_314),
.Y(n_370)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_322),
.A2(n_292),
.B1(n_293),
.B2(n_303),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_336),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_346),
.A2(n_303),
.B1(n_296),
.B2(n_305),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_333),
.A2(n_296),
.B1(n_305),
.B2(n_257),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_379),
.B1(n_365),
.B2(n_358),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_330),
.B(n_254),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_324),
.A2(n_270),
.B1(n_276),
.B2(n_205),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_374),
.B(n_347),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_381),
.B(n_388),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_319),
.B1(n_345),
.B2(n_324),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_384),
.A2(n_396),
.B1(n_397),
.B2(n_400),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_404),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_350),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_350),
.B(n_339),
.Y(n_389)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_368),
.B(n_373),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_390),
.B(n_391),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_357),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_332),
.C(n_320),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_392),
.B(n_395),
.C(n_401),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_327),
.C(n_323),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_328),
.B1(n_349),
.B2(n_343),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_361),
.B(n_341),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_385),
.Y(n_412)
);

OAI22x1_ASAP7_75t_L g400 ( 
.A1(n_370),
.A2(n_348),
.B1(n_335),
.B2(n_321),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_318),
.C(n_317),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_372),
.B1(n_355),
.B2(n_367),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_236),
.C(n_225),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_403),
.B(n_376),
.C(n_364),
.Y(n_410)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_380),
.A2(n_359),
.B(n_379),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_405),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_407),
.A2(n_414),
.B1(n_421),
.B2(n_397),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_410),
.B(n_411),
.C(n_417),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_364),
.C(n_353),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_229),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_360),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_394),
.A2(n_367),
.B1(n_353),
.B2(n_203),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_166),
.Y(n_415)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_165),
.C(n_120),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_387),
.A2(n_201),
.B1(n_162),
.B2(n_153),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_100),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_393),
.A2(n_120),
.B1(n_109),
.B2(n_105),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_406),
.A2(n_387),
.B1(n_404),
.B2(n_394),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_423),
.A2(n_424),
.B1(n_427),
.B2(n_146),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_419),
.A2(n_380),
.B1(n_398),
.B2(n_384),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_399),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_425),
.A2(n_409),
.B(n_416),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_426),
.A2(n_434),
.B1(n_430),
.B2(n_423),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_416),
.A2(n_383),
.B1(n_395),
.B2(n_392),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_422),
.B(n_385),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_428),
.B(n_432),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_430),
.B(n_434),
.C(n_417),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_418),
.B(n_14),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_433),
.B(n_15),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_229),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_439),
.B(n_443),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_438),
.B(n_446),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_429),
.B(n_411),
.C(n_408),
.Y(n_439)
);

AOI21x1_ASAP7_75t_SL g440 ( 
.A1(n_435),
.A2(n_415),
.B(n_413),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_441),
.A2(n_444),
.B1(n_424),
.B2(n_105),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_431),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_442),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_408),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_223),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_223),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_454),
.Y(n_461)
);

AOI322xp5_ASAP7_75t_L g457 ( 
.A1(n_450),
.A2(n_437),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_12),
.C2(n_13),
.Y(n_457)
);

AOI21xp33_ASAP7_75t_L g451 ( 
.A1(n_442),
.A2(n_10),
.B(n_2),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_451),
.A2(n_436),
.B(n_5),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_446),
.A2(n_110),
.B1(n_126),
.B2(n_129),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_452),
.A2(n_453),
.B1(n_13),
.B2(n_15),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_440),
.A2(n_110),
.B1(n_2),
.B2(n_3),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_444),
.A2(n_7),
.B1(n_2),
.B2(n_5),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_456),
.B(n_459),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_458),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_455),
.B(n_439),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_438),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_449),
.A2(n_7),
.B(n_10),
.C(n_12),
.Y(n_460)
);

AOI322xp5_ASAP7_75t_L g466 ( 
.A1(n_460),
.A2(n_1),
.A3(n_223),
.B1(n_291),
.B2(n_325),
.C1(n_154),
.C2(n_338),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_462),
.A2(n_449),
.B1(n_452),
.B2(n_453),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_464),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_466),
.Y(n_468)
);

OA21x2_ASAP7_75t_SL g469 ( 
.A1(n_468),
.A2(n_465),
.B(n_463),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_469),
.B(n_470),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_467),
.B(n_463),
.C(n_461),
.Y(n_470)
);


endmodule