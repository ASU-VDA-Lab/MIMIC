module fake_jpeg_6426_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx12_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_15),
.A2(n_3),
.B1(n_7),
.B2(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_17),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_19),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

AO21x2_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_22),
.B(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_15),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_29),
.B1(n_17),
.B2(n_12),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_24),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_28),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_6),
.B(n_8),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_27),
.C(n_29),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_37),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_28),
.C(n_6),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_32),
.B1(n_28),
.B2(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_40),
.Y(n_41)
);

MAJx2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_37),
.C(n_6),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_SL g44 ( 
.A(n_42),
.B(n_14),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_3),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_45),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_41),
.B(n_42),
.Y(n_47)
);


endmodule