module fake_jpeg_19248_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx12_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_0),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_31),
.C(n_32),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_27),
.A2(n_29),
.B1(n_11),
.B2(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_7),
.Y(n_29)
);

INVxp67_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_34),
.A2(n_42),
.B1(n_32),
.B2(n_31),
.Y(n_50)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_25),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_26),
.B(n_24),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_26),
.A2(n_17),
.B1(n_15),
.B2(n_12),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_13),
.B1(n_12),
.B2(n_22),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_43),
.A2(n_13),
.B1(n_20),
.B2(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_56),
.Y(n_58)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_22),
.C(n_29),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_43),
.C(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_22),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_43),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_58),
.B(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_34),
.B1(n_38),
.B2(n_42),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_56),
.A2(n_38),
.B1(n_33),
.B2(n_35),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_35),
.B1(n_43),
.B2(n_14),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_43),
.C(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_54),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_70),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_64),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_58),
.B1(n_60),
.B2(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_48),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_63),
.B(n_62),
.C(n_57),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_86),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_85),
.A2(n_72),
.B(n_3),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_57),
.B1(n_36),
.B2(n_40),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_83),
.C(n_84),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_89),
.Y(n_95)
);

A2O1A1O1Ixp25_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_76),
.B(n_71),
.C(n_73),
.D(n_69),
.Y(n_88)
);

OAI211xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_90),
.B(n_92),
.C(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_69),
.Y(n_90)
);

NOR2xp67_ASAP7_75t_SL g93 ( 
.A(n_91),
.B(n_86),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_2),
.B(n_4),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_96),
.Y(n_97)
);

OAI221xp5_ASAP7_75t_L g96 ( 
.A1(n_91),
.A2(n_83),
.B1(n_85),
.B2(n_36),
.C(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_97),
.B(n_8),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_9),
.C(n_10),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_102),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_10),
.Y(n_106)
);


endmodule