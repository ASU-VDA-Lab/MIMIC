module fake_jpeg_18905_n_99 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_99);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx4f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_2),
.B(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_26),
.Y(n_31)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_21),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_38),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_23),
.A2(n_19),
.B1(n_17),
.B2(n_22),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_40),
.B1(n_35),
.B2(n_33),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_19),
.B1(n_17),
.B2(n_12),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_13),
.B1(n_15),
.B2(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_38),
.B(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_42),
.B(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_26),
.B1(n_30),
.B2(n_13),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_46),
.B1(n_54),
.B2(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_45),
.B(n_53),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_15),
.B1(n_11),
.B2(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_11),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_50),
.B(n_54),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_14),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_37),
.B1(n_33),
.B2(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_57),
.B1(n_8),
.B2(n_10),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_56),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_4),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_59),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_7),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_65),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_53),
.B(n_45),
.C(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_71),
.B(n_59),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_49),
.B(n_57),
.C(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_50),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_70),
.C(n_68),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_69),
.Y(n_81)
);

NOR4xp25_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_60),
.C(n_61),
.D(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_84),
.Y(n_88)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_73),
.B1(n_62),
.B2(n_75),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_90),
.B1(n_82),
.B2(n_85),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_87),
.C(n_86),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_93),
.A2(n_64),
.B(n_91),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.C(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);


endmodule