module fake_jpeg_6516_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_26),
.Y(n_61)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_61),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_32),
.B1(n_26),
.B2(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_32),
.B1(n_17),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_73),
.B1(n_28),
.B2(n_24),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_32),
.B1(n_26),
.B2(n_18),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_60),
.B(n_30),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_32),
.B1(n_18),
.B2(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_21),
.B1(n_22),
.B2(n_16),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_70),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_20),
.B1(n_28),
.B2(n_30),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_21),
.B1(n_22),
.B2(n_16),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_45),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_46),
.B1(n_41),
.B2(n_37),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_52),
.B1(n_64),
.B2(n_71),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_88),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_45),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_54),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_45),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_88),
.C(n_78),
.Y(n_111)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_60),
.B1(n_59),
.B2(n_24),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_92),
.B1(n_93),
.B2(n_81),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_25),
.B1(n_27),
.B2(n_23),
.Y(n_157)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_116),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_48),
.B1(n_53),
.B2(n_59),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_75),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_52),
.B1(n_72),
.B2(n_37),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_124),
.B1(n_94),
.B2(n_91),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_115),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_95),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_84),
.B1(n_97),
.B2(n_75),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_85),
.B1(n_97),
.B2(n_96),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_119),
.A2(n_122),
.B1(n_123),
.B2(n_79),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_46),
.B1(n_41),
.B2(n_31),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_76),
.A2(n_27),
.B(n_33),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_127),
.B(n_79),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_46),
.B(n_41),
.C(n_27),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_83),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_135),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_101),
.B(n_89),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_140),
.C(n_129),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_146),
.B1(n_149),
.B2(n_156),
.Y(n_159)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_84),
.B(n_90),
.C(n_75),
.D(n_27),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_136),
.A2(n_112),
.B(n_126),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_84),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_144),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_139),
.A2(n_153),
.B(n_137),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_157),
.B1(n_127),
.B2(n_116),
.Y(n_164)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_77),
.B1(n_65),
.B2(n_49),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_113),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_77),
.B1(n_65),
.B2(n_49),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_151),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_100),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_122),
.A2(n_80),
.B(n_27),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_80),
.B1(n_67),
.B2(n_23),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_111),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_147),
.B(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_25),
.B1(n_33),
.B2(n_105),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_133),
.A2(n_103),
.B(n_125),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_165),
.A2(n_178),
.B(n_187),
.Y(n_211)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_181),
.C(n_186),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_174),
.A2(n_176),
.B(n_182),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_123),
.A3(n_114),
.B1(n_102),
.B2(n_23),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_185),
.B1(n_119),
.B2(n_104),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_150),
.B1(n_140),
.B2(n_157),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_154),
.B1(n_152),
.B2(n_25),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_50),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_135),
.B(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_67),
.B1(n_112),
.B2(n_23),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_50),
.C(n_54),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_33),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_141),
.B(n_134),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_162),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_149),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_202),
.C(n_205),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_185),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_130),
.B1(n_144),
.B2(n_152),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_152),
.B1(n_102),
.B2(n_115),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_208),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_172),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_50),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_54),
.C(n_154),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_166),
.C(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_180),
.B1(n_164),
.B2(n_187),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_170),
.A2(n_154),
.B1(n_54),
.B2(n_2),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_0),
.Y(n_214)
);

NOR2x1_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_185),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_169),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_216),
.B(n_226),
.Y(n_257)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_214),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_182),
.B1(n_171),
.B2(n_174),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_219),
.A2(n_238),
.B1(n_239),
.B2(n_242),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_187),
.B1(n_159),
.B2(n_162),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_221),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_179),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_224),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_199),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_223),
.A2(n_228),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_186),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_237),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

XOR2x2_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_185),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_229),
.B(n_205),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_204),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g247 ( 
.A(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_241),
.C(n_193),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_189),
.B(n_161),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_175),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_240),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_158),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_207),
.A2(n_175),
.B1(n_158),
.B2(n_2),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_246),
.Y(n_267)
);

XOR2x1_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_204),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_4),
.B(n_5),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_211),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_245),
.B(n_266),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_248),
.B(n_253),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_265),
.Y(n_270)
);

NOR3xp33_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_188),
.C(n_196),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_196),
.B1(n_203),
.B2(n_206),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_254),
.A2(n_256),
.B1(n_3),
.B2(n_4),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_208),
.B1(n_201),
.B2(n_193),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_3),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_237),
.C(n_218),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_225),
.B1(n_227),
.B2(n_8),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_220),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_218),
.B(n_15),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_272),
.C(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_221),
.B1(n_220),
.B2(n_217),
.Y(n_271)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_241),
.C(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_250),
.Y(n_287)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_277),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_8),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_251),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_259),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_13),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_4),
.C(n_5),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_252),
.B(n_248),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_286),
.A2(n_298),
.B(n_276),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_253),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_13),
.B(n_6),
.Y(n_314)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_245),
.B1(n_255),
.B2(n_263),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_271),
.B1(n_269),
.B2(n_285),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_274),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_273),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_272),
.B(n_263),
.C(n_266),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_276),
.C(n_281),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_301),
.B(n_10),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_309),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_277),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_304),
.A2(n_307),
.B(n_313),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_278),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_315),
.C(n_300),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_10),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_293),
.B(n_298),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_10),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_289),
.A2(n_11),
.B(n_12),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_290),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_286),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_320),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_295),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_309),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_322),
.C(n_295),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_315),
.B(n_292),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_291),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_327),
.B(n_328),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_302),
.C(n_288),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_330),
.A2(n_333),
.B(n_324),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_314),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_311),
.C(n_6),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_337),
.B(n_338),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_329),
.B(n_317),
.Y(n_337)
);

AO21x2_ASAP7_75t_L g340 ( 
.A1(n_336),
.A2(n_325),
.B(n_6),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_334),
.C(n_339),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_342),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_343),
.A2(n_7),
.B(n_334),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);


endmodule