module fake_aes_7212_n_1153 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1153);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1153;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_384;
wire n_434;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1098;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1125;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_1101;
wire n_630;
wire n_1078;
wire n_511;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_725;
wire n_769;
wire n_844;
wire n_818;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_1138;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_771;
wire n_696;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_1089;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_1110;
wire n_327;
wire n_944;
wire n_325;
wire n_1131;
wire n_1102;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_912;
wire n_924;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1117;
wire n_859;
wire n_1007;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_251), .Y(n_278) );
INVxp67_ASAP7_75t_L g279 ( .A(n_177), .Y(n_279) );
BUFx10_ASAP7_75t_L g280 ( .A(n_243), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_89), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_233), .Y(n_282) );
BUFx2_ASAP7_75t_SL g283 ( .A(n_69), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_178), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_5), .Y(n_285) );
CKINVDCx16_ASAP7_75t_R g286 ( .A(n_276), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_15), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_53), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_208), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_202), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_5), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_193), .Y(n_292) );
CKINVDCx14_ASAP7_75t_R g293 ( .A(n_277), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_131), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_122), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_69), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_230), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_248), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_253), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_20), .Y(n_300) );
INVxp33_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_192), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_90), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_109), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_225), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_34), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_222), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_212), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_124), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_181), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_170), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_119), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_142), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_125), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_167), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_22), .Y(n_316) );
INVxp67_ASAP7_75t_L g317 ( .A(n_38), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_273), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_197), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_191), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_132), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_267), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_102), .Y(n_323) );
CKINVDCx20_ASAP7_75t_R g324 ( .A(n_78), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_224), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_150), .Y(n_326) );
INVxp33_ASAP7_75t_L g327 ( .A(n_262), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_30), .Y(n_328) );
INVxp67_ASAP7_75t_SL g329 ( .A(n_43), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_226), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_97), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_59), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_220), .Y(n_333) );
INVxp33_ASAP7_75t_L g334 ( .A(n_199), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_218), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_201), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_213), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_274), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_44), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_183), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_74), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_143), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_237), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_171), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_241), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_203), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_101), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_114), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_235), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_250), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_244), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_259), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_257), .Y(n_353) );
INVxp33_ASAP7_75t_L g354 ( .A(n_242), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_146), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_51), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_258), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_151), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_84), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_145), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_264), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_8), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_166), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_271), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_1), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_117), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_25), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_60), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_169), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_140), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_82), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_196), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_13), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_263), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_16), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_200), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_190), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_223), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_82), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_186), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_36), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_12), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_2), .Y(n_383) );
BUFx5_ASAP7_75t_L g384 ( .A(n_275), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_121), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_165), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_174), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_184), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g389 ( .A(n_204), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_112), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_182), .Y(n_391) );
BUFx3_ASAP7_75t_L g392 ( .A(n_80), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_260), .Y(n_393) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_168), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_231), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_207), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_187), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_159), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_136), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_101), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_54), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_12), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_185), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_240), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_139), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_228), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_65), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_127), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_130), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_49), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_249), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_60), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_272), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_138), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_211), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_110), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g417 ( .A(n_26), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g418 ( .A(n_198), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_214), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_148), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_102), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_80), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_133), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_56), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_219), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_64), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_61), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_127), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_17), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g430 ( .A(n_128), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_24), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_104), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_383), .B(n_0), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_303), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_292), .B(n_0), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_297), .B(n_1), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_322), .B(n_2), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_303), .B(n_3), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_384), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_303), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_337), .B(n_4), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_330), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_367), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g444 ( .A1(n_291), .A2(n_7), .B1(n_4), .B2(n_6), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_384), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_367), .B(n_6), .Y(n_446) );
INVx5_ASAP7_75t_L g447 ( .A(n_374), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_367), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_286), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_420), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_330), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_374), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_338), .B(n_420), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_316), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_374), .B(n_343), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_384), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_280), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_330), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_326), .Y(n_460) );
OAI21x1_ASAP7_75t_L g461 ( .A1(n_282), .A2(n_164), .B(n_163), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_316), .Y(n_462) );
XOR2x2_ASAP7_75t_SL g463 ( .A(n_331), .B(n_379), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_330), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_343), .B(n_7), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_355), .A2(n_10), .B1(n_8), .B2(n_9), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_375), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_375), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_381), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_430), .A2(n_13), .B1(n_10), .B2(n_11), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_384), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_347), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_384), .Y(n_473) );
BUFx8_ASAP7_75t_L g474 ( .A(n_384), .Y(n_474) );
OR2x6_ASAP7_75t_L g475 ( .A(n_444), .B(n_283), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_460), .B(n_285), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_433), .A2(n_281), .B1(n_294), .B2(n_287), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_453), .B(n_425), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_458), .B(n_301), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_460), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_458), .B(n_327), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_440), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_440), .Y(n_484) );
AND2x6_ASAP7_75t_L g485 ( .A(n_438), .B(n_284), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_453), .B(n_285), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_453), .B(n_334), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_458), .B(n_354), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_472), .B(n_280), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_439), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_440), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_439), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_458), .B(n_288), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_463), .B(n_280), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_456), .B(n_331), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_445), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_445), .Y(n_500) );
NOR2x1p5_ASAP7_75t_L g501 ( .A(n_449), .B(n_304), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_456), .B(n_279), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_433), .A2(n_319), .B1(n_352), .B2(n_305), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_445), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_472), .B(n_312), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_457), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_456), .B(n_340), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_457), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_456), .B(n_312), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_471), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_433), .B(n_347), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_471), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_471), .Y(n_515) );
INVx3_ASAP7_75t_L g516 ( .A(n_438), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_516), .B(n_463), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_516), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_490), .B(n_436), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_492), .B(n_436), .Y(n_520) );
INVx2_ASAP7_75t_SL g521 ( .A(n_492), .Y(n_521) );
OR2x6_ASAP7_75t_L g522 ( .A(n_475), .B(n_466), .Y(n_522) );
AND2x4_ASAP7_75t_L g523 ( .A(n_513), .B(n_436), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_487), .B(n_456), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_516), .B(n_465), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_479), .B(n_435), .Y(n_526) );
NOR2x1p5_ASAP7_75t_L g527 ( .A(n_476), .B(n_435), .Y(n_527) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_475), .A2(n_324), .B1(n_328), .B2(n_291), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_483), .A2(n_461), .B(n_465), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_498), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_485), .A2(n_438), .B1(n_446), .B2(n_474), .Y(n_531) );
AND2x2_ASAP7_75t_SL g532 ( .A(n_503), .B(n_438), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_511), .B(n_437), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_480), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_498), .Y(n_535) );
AND2x6_ASAP7_75t_L g536 ( .A(n_498), .B(n_465), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_485), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_482), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_485), .A2(n_438), .B1(n_446), .B2(n_474), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_513), .Y(n_540) );
AO22x1_ASAP7_75t_L g541 ( .A1(n_485), .A2(n_470), .B1(n_466), .B2(n_474), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_485), .A2(n_446), .B1(n_474), .B2(n_465), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_506), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_481), .B(n_441), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_497), .A2(n_446), .B1(n_319), .B2(n_389), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_482), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_486), .B(n_358), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_478), .B(n_358), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_496), .B(n_474), .Y(n_549) );
OR2x6_ASAP7_75t_L g550 ( .A(n_475), .B(n_470), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_483), .B(n_446), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_502), .B(n_434), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_508), .B(n_434), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_485), .B(n_443), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_484), .B(n_443), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_503), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_484), .A2(n_461), .B(n_473), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_488), .Y(n_558) );
BUFx8_ASAP7_75t_L g559 ( .A(n_495), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_501), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_489), .B(n_448), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_488), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_501), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_477), .A2(n_365), .B1(n_371), .B2(n_360), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_495), .A2(n_452), .B1(n_448), .B2(n_450), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_491), .B(n_450), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_491), .B(n_454), .Y(n_568) );
OR2x6_ASAP7_75t_L g569 ( .A(n_505), .B(n_379), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_499), .B(n_360), .Y(n_570) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
BUFx6f_ASAP7_75t_SL g572 ( .A(n_500), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_494), .B(n_447), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_507), .B(n_447), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_504), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_493), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_509), .A2(n_461), .B(n_452), .C(n_455), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_510), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_510), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_512), .B(n_447), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_512), .B(n_447), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_514), .B(n_447), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_514), .B(n_447), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_515), .B(n_278), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_505), .B(n_289), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_505), .B(n_473), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_480), .B(n_401), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_490), .B(n_289), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_516), .B(n_473), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_534), .B(n_407), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_542), .A2(n_293), .B1(n_416), .B2(n_407), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_529), .A2(n_452), .B(n_394), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_522), .A2(n_416), .B1(n_421), .B2(n_417), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_559), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_559), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_530), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_531), .B(n_539), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_517), .A2(n_408), .B(n_317), .C(n_329), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_571), .Y(n_600) );
NOR2xp33_ASAP7_75t_SL g601 ( .A(n_572), .B(n_423), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_517), .A2(n_431), .B(n_424), .C(n_296), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_572), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_547), .B(n_423), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g605 ( .A1(n_552), .A2(n_382), .B(n_392), .C(n_356), .Y(n_605) );
AOI21x1_ASAP7_75t_L g606 ( .A1(n_557), .A2(n_307), .B(n_302), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_519), .B(n_426), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_542), .A2(n_427), .B1(n_426), .B2(n_298), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_520), .A2(n_300), .B(n_306), .C(n_295), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_551), .A2(n_320), .B(n_310), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_532), .A2(n_527), .B1(n_521), .B2(n_548), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_540), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_555), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_518), .Y(n_614) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_537), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_589), .A2(n_336), .B(n_335), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_524), .A2(n_313), .B(n_314), .C(n_309), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_523), .B(n_321), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_577), .A2(n_346), .B(n_345), .Y(n_619) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_560), .A2(n_350), .B(n_349), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_523), .B(n_341), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_564), .B(n_348), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_536), .A2(n_382), .B1(n_392), .B2(n_356), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_575), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_543), .B(n_422), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_SL g626 ( .A1(n_549), .A2(n_351), .B(n_357), .C(n_353), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_589), .A2(n_369), .B(n_363), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_570), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_561), .B(n_366), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_578), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_536), .A2(n_402), .B1(n_429), .B2(n_400), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_536), .A2(n_402), .B1(n_429), .B2(n_400), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_573), .A2(n_377), .B(n_376), .Y(n_633) );
INVx3_ASAP7_75t_L g634 ( .A(n_569), .Y(n_634) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_545), .B(n_311), .C(n_308), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_587), .Y(n_636) );
OR2x6_ASAP7_75t_L g637 ( .A(n_522), .B(n_381), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_526), .A2(n_325), .B1(n_333), .B2(n_315), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_578), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_562), .A2(n_568), .B(n_567), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_522), .A2(n_332), .B1(n_339), .B2(n_323), .Y(n_641) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_569), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_565), .B(n_462), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_544), .A2(n_359), .B(n_362), .C(n_342), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_579), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_588), .B(n_361), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_579), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_553), .A2(n_370), .B(n_373), .C(n_368), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_528), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_554), .A2(n_380), .B(n_378), .Y(n_650) );
NOR3xp33_ASAP7_75t_SL g651 ( .A(n_541), .B(n_386), .C(n_364), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_550), .A2(n_387), .B1(n_388), .B2(n_386), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_585), .B(n_387), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_586), .A2(n_396), .B(n_391), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_584), .B(n_388), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_566), .B(n_393), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_538), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_586), .A2(n_403), .B(n_397), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_546), .B(n_393), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_581), .A2(n_406), .B(n_404), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_550), .B(n_385), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_546), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_558), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_563), .A2(n_398), .B1(n_399), .B2(n_390), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_583), .A2(n_409), .B(n_410), .C(n_405), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_576), .B(n_413), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_574), .B(n_418), .Y(n_667) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_574), .Y(n_668) );
INVx4_ASAP7_75t_SL g669 ( .A(n_583), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_580), .A2(n_419), .B1(n_418), .B2(n_414), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_582), .A2(n_415), .B(n_411), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_525), .A2(n_290), .B(n_282), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_532), .A2(n_428), .B1(n_432), .B2(n_412), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_533), .B(n_467), .Y(n_674) );
AND3x1_ASAP7_75t_SL g675 ( .A(n_527), .B(n_468), .C(n_467), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_533), .B(n_468), .Y(n_676) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_542), .B(n_344), .C(n_318), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_534), .B(n_469), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_571), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_525), .A2(n_299), .B(n_290), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_559), .Y(n_681) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_571), .Y(n_682) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_571), .Y(n_683) );
CKINVDCx5p33_ASAP7_75t_R g684 ( .A(n_559), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_684), .Y(n_685) );
AOI31xp67_ASAP7_75t_L g686 ( .A1(n_598), .A2(n_451), .A3(n_459), .B(n_442), .Y(n_686) );
AO32x2_ASAP7_75t_L g687 ( .A1(n_591), .A2(n_442), .A3(n_464), .B1(n_459), .B2(n_451), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_662), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_612), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_640), .A2(n_644), .B(n_617), .C(n_648), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_624), .Y(n_691) );
AND2x4_ASAP7_75t_L g692 ( .A(n_594), .B(n_14), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_636), .B(n_15), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g694 ( .A(n_601), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_613), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_611), .B(n_17), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_592), .A2(n_395), .B(n_372), .Y(n_697) );
OAI21x1_ASAP7_75t_L g698 ( .A1(n_606), .A2(n_395), .B(n_442), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_643), .B(n_18), .Y(n_699) );
AO21x1_ASAP7_75t_L g700 ( .A1(n_619), .A2(n_451), .B(n_442), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_673), .B(n_18), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_662), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_673), .A2(n_451), .B1(n_459), .B2(n_442), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_681), .B(n_19), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_674), .Y(n_705) );
AO32x2_ASAP7_75t_L g706 ( .A1(n_652), .A2(n_464), .A3(n_459), .B1(n_451), .B2(n_23), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_593), .B(n_21), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_609), .A2(n_464), .B(n_459), .C(n_23), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_593), .B(n_21), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_604), .B(n_24), .Y(n_710) );
AO31x2_ASAP7_75t_L g711 ( .A1(n_605), .A2(n_29), .A3(n_27), .B(n_28), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_676), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_678), .B(n_31), .Y(n_713) );
BUFx3_ASAP7_75t_L g714 ( .A(n_603), .Y(n_714) );
INVx1_ASAP7_75t_SL g715 ( .A(n_642), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_663), .A2(n_173), .B(n_172), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_590), .B(n_31), .Y(n_717) );
OR2x6_ASAP7_75t_L g718 ( .A(n_637), .B(n_32), .Y(n_718) );
A2O1A1Ixp33_ASAP7_75t_L g719 ( .A1(n_602), .A2(n_36), .B(n_33), .C(n_35), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_600), .A2(n_176), .B(n_175), .Y(n_720) );
AND2x6_ASAP7_75t_L g721 ( .A(n_634), .B(n_37), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_679), .A2(n_180), .B(n_179), .Y(n_722) );
INVx5_ASAP7_75t_L g723 ( .A(n_634), .Y(n_723) );
BUFx10_ASAP7_75t_L g724 ( .A(n_661), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_607), .B(n_39), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_641), .B(n_40), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_657), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_L g728 ( .A1(n_665), .A2(n_42), .B(n_40), .C(n_41), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_682), .Y(n_729) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_641), .A2(n_45), .B1(n_43), .B2(n_44), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_669), .B(n_46), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_630), .Y(n_732) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_625), .A2(n_621), .B1(n_618), .B2(n_664), .C(n_649), .Y(n_733) );
AOI221xp5_ASAP7_75t_SL g734 ( .A1(n_599), .A2(n_47), .B1(n_48), .B2(n_49), .C(n_50), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_596), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_597), .Y(n_736) );
AO31x2_ASAP7_75t_L g737 ( .A1(n_672), .A2(n_53), .A3(n_51), .B(n_52), .Y(n_737) );
AO31x2_ASAP7_75t_L g738 ( .A1(n_680), .A2(n_55), .A3(n_52), .B(n_54), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_622), .B(n_55), .Y(n_739) );
OAI22x1_ASAP7_75t_L g740 ( .A1(n_675), .A2(n_58), .B1(n_56), .B2(n_57), .Y(n_740) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_639), .A2(n_189), .B(n_188), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_645), .A2(n_195), .B(n_194), .Y(n_742) );
A2O1A1Ixp33_ASAP7_75t_L g743 ( .A1(n_610), .A2(n_59), .B(n_57), .C(n_58), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_647), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g745 ( .A1(n_660), .A2(n_63), .B(n_61), .C(n_62), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_650), .A2(n_62), .B(n_63), .C(n_64), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_614), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_664), .B(n_66), .Y(n_748) );
O2A1O1Ixp33_ASAP7_75t_L g749 ( .A1(n_626), .A2(n_67), .B(n_68), .C(n_70), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_L g750 ( .A1(n_654), .A2(n_68), .B(n_70), .C(n_71), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_651), .Y(n_751) );
AO31x2_ASAP7_75t_L g752 ( .A1(n_658), .A2(n_71), .A3(n_72), .B(n_73), .Y(n_752) );
AO31x2_ASAP7_75t_L g753 ( .A1(n_616), .A2(n_75), .A3(n_76), .B(n_77), .Y(n_753) );
BUFx12f_ASAP7_75t_L g754 ( .A(n_668), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_635), .A2(n_76), .B1(n_77), .B2(n_78), .Y(n_755) );
A2O1A1Ixp33_ASAP7_75t_L g756 ( .A1(n_627), .A2(n_79), .B(n_81), .C(n_83), .Y(n_756) );
AO31x2_ASAP7_75t_L g757 ( .A1(n_633), .A2(n_83), .A3(n_84), .B(n_85), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_620), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g759 ( .A1(n_671), .A2(n_85), .B(n_86), .C(n_87), .Y(n_759) );
AOI221xp5_ASAP7_75t_SL g760 ( .A1(n_608), .A2(n_86), .B1(n_87), .B2(n_88), .C(n_89), .Y(n_760) );
NOR2xp33_ASAP7_75t_SL g761 ( .A(n_677), .B(n_88), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_638), .B(n_91), .Y(n_762) );
AND2x6_ASAP7_75t_L g763 ( .A(n_615), .B(n_91), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_659), .Y(n_764) );
OAI21x1_ASAP7_75t_L g765 ( .A1(n_623), .A2(n_206), .B(n_205), .Y(n_765) );
BUFx5_ASAP7_75t_L g766 ( .A(n_682), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_666), .Y(n_767) );
BUFx6f_ASAP7_75t_L g768 ( .A(n_682), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_655), .A2(n_210), .B(n_209), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g770 ( .A1(n_632), .A2(n_92), .B(n_93), .C(n_94), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_656), .B(n_92), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_629), .B(n_93), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_667), .Y(n_773) );
OAI21xp5_ASAP7_75t_L g774 ( .A1(n_631), .A2(n_216), .B(n_215), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_670), .A2(n_95), .B1(n_96), .B2(n_98), .Y(n_775) );
BUFx3_ASAP7_75t_L g776 ( .A(n_683), .Y(n_776) );
A2O1A1Ixp33_ASAP7_75t_L g777 ( .A1(n_653), .A2(n_99), .B(n_100), .C(n_103), .Y(n_777) );
A2O1A1Ixp33_ASAP7_75t_L g778 ( .A1(n_646), .A2(n_99), .B(n_100), .C(n_103), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g779 ( .A1(n_675), .A2(n_270), .B(n_269), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_669), .Y(n_780) );
AOI21xp5_ASAP7_75t_L g781 ( .A1(n_615), .A2(n_245), .B(n_265), .Y(n_781) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_615), .Y(n_782) );
AOI22xp33_ASAP7_75t_SL g783 ( .A1(n_615), .A2(n_105), .B1(n_106), .B2(n_107), .Y(n_783) );
AO31x2_ASAP7_75t_L g784 ( .A1(n_669), .A2(n_106), .A3(n_107), .B(n_108), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_640), .A2(n_266), .B(n_261), .Y(n_785) );
INVx4_ASAP7_75t_L g786 ( .A(n_595), .Y(n_786) );
OR2x2_ASAP7_75t_L g787 ( .A(n_715), .B(n_111), .Y(n_787) );
OAI21xp33_ASAP7_75t_L g788 ( .A1(n_761), .A2(n_113), .B(n_115), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_707), .A2(n_116), .B1(n_117), .B2(n_118), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_709), .A2(n_118), .B1(n_119), .B2(n_120), .Y(n_790) );
BUFx3_ASAP7_75t_L g791 ( .A(n_786), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_689), .Y(n_792) );
A2O1A1Ixp33_ASAP7_75t_L g793 ( .A1(n_758), .A2(n_123), .B(n_126), .C(n_129), .Y(n_793) );
OA21x2_ASAP7_75t_L g794 ( .A1(n_700), .A2(n_256), .B(n_255), .Y(n_794) );
OA21x2_ASAP7_75t_L g795 ( .A1(n_779), .A2(n_254), .B(n_252), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_691), .Y(n_796) );
CKINVDCx11_ASAP7_75t_R g797 ( .A(n_786), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_726), .A2(n_134), .B1(n_135), .B2(n_137), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_692), .B(n_135), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_735), .Y(n_800) );
AO21x2_ASAP7_75t_L g801 ( .A1(n_774), .A2(n_247), .B(n_246), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_688), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_702), .Y(n_803) );
OR2x6_ASAP7_75t_L g804 ( .A(n_692), .B(n_141), .Y(n_804) );
INVx4_ASAP7_75t_SL g805 ( .A(n_721), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_736), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_693), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_772), .A2(n_144), .B1(n_146), .B2(n_147), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g809 ( .A(n_694), .Y(n_809) );
BUFx5_ASAP7_75t_L g810 ( .A(n_776), .Y(n_810) );
OA21x2_ASAP7_75t_L g811 ( .A1(n_760), .A2(n_217), .B(n_238), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_740), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_721), .Y(n_813) );
BUFx2_ASAP7_75t_L g814 ( .A(n_754), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_721), .Y(n_815) );
AO31x2_ASAP7_75t_L g816 ( .A1(n_708), .A2(n_149), .A3(n_151), .B(n_152), .Y(n_816) );
BUFx6f_ASAP7_75t_L g817 ( .A(n_729), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_717), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_713), .B(n_153), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_730), .A2(n_154), .B1(n_155), .B2(n_156), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_721), .Y(n_821) );
OA21x2_ASAP7_75t_L g822 ( .A1(n_765), .A2(n_221), .B(n_236), .Y(n_822) );
INVx3_ASAP7_75t_L g823 ( .A(n_731), .Y(n_823) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_785), .A2(n_239), .B(n_234), .Y(n_824) );
NAND2x1_ASAP7_75t_L g825 ( .A(n_763), .B(n_232), .Y(n_825) );
INVx6_ASAP7_75t_L g826 ( .A(n_724), .Y(n_826) );
INVx4_ASAP7_75t_SL g827 ( .A(n_763), .Y(n_827) );
BUFx4f_ASAP7_75t_SL g828 ( .A(n_714), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_755), .A2(n_157), .B1(n_158), .B2(n_159), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_704), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_724), .B(n_160), .Y(n_831) );
A2O1A1Ixp33_ASAP7_75t_L g832 ( .A1(n_739), .A2(n_161), .B(n_162), .C(n_227), .Y(n_832) );
A2O1A1Ixp33_ASAP7_75t_L g833 ( .A1(n_749), .A2(n_229), .B(n_755), .C(n_771), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_747), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_748), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_699), .A2(n_731), .B1(n_701), .B2(n_696), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_710), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_752), .Y(n_838) );
BUFx12f_ASAP7_75t_L g839 ( .A(n_685), .Y(n_839) );
INVx3_ASAP7_75t_L g840 ( .A(n_763), .Y(n_840) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_727), .Y(n_841) );
NOR2xp33_ASAP7_75t_SL g842 ( .A(n_780), .B(n_751), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_725), .B(n_762), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_752), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_764), .B(n_767), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_752), .Y(n_846) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_729), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_723), .B(n_732), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_753), .Y(n_849) );
O2A1O1Ixp33_ASAP7_75t_L g850 ( .A1(n_719), .A2(n_778), .B(n_728), .C(n_777), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_773), .B(n_723), .Y(n_851) );
NOR2x1_ASAP7_75t_SL g852 ( .A(n_723), .B(n_729), .Y(n_852) );
OAI22xp5_ASAP7_75t_L g853 ( .A1(n_703), .A2(n_775), .B1(n_770), .B2(n_783), .Y(n_853) );
BUFx8_ASAP7_75t_L g854 ( .A(n_706), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_744), .B(n_734), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_753), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_769), .A2(n_746), .B(n_750), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_753), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_711), .B(n_757), .Y(n_859) );
AOI21x1_ASAP7_75t_L g860 ( .A1(n_716), .A2(n_686), .B(n_742), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_757), .Y(n_861) );
NAND2x1p5_ASAP7_75t_L g862 ( .A(n_768), .B(n_782), .Y(n_862) );
NAND2x1_ASAP7_75t_L g863 ( .A(n_782), .B(n_781), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_745), .A2(n_743), .B(n_756), .C(n_759), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_757), .Y(n_865) );
OA21x2_ASAP7_75t_L g866 ( .A1(n_741), .A2(n_722), .B(n_720), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_711), .B(n_737), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_706), .Y(n_868) );
INVx4_ASAP7_75t_L g869 ( .A(n_766), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g870 ( .A(n_766), .B(n_784), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g871 ( .A1(n_766), .A2(n_784), .B1(n_737), .B2(n_738), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_766), .A2(n_687), .B1(n_784), .B2(n_737), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_738), .B(n_766), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_697), .A2(n_592), .B(n_529), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_695), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_697), .A2(n_592), .B(n_529), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_695), .Y(n_877) );
OA21x2_ASAP7_75t_L g878 ( .A1(n_698), .A2(n_700), .B(n_697), .Y(n_878) );
A2O1A1Ixp33_ASAP7_75t_L g879 ( .A1(n_690), .A2(n_712), .B(n_705), .C(n_758), .Y(n_879) );
INVx6_ASAP7_75t_L g880 ( .A(n_786), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_705), .B(n_712), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_705), .B(n_712), .Y(n_882) );
OA21x2_ASAP7_75t_L g883 ( .A1(n_698), .A2(n_700), .B(n_697), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g884 ( .A(n_733), .B(n_556), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_697), .A2(n_592), .B(n_529), .Y(n_885) );
AND2x2_ASAP7_75t_L g886 ( .A(n_695), .B(n_628), .Y(n_886) );
AO31x2_ASAP7_75t_L g887 ( .A1(n_700), .A2(n_697), .A3(n_577), .B(n_758), .Y(n_887) );
OA21x2_ASAP7_75t_L g888 ( .A1(n_698), .A2(n_700), .B(n_697), .Y(n_888) );
AND2x2_ASAP7_75t_L g889 ( .A(n_695), .B(n_628), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g890 ( .A1(n_718), .A2(n_673), .B1(n_637), .B2(n_758), .Y(n_890) );
OR2x6_ASAP7_75t_L g891 ( .A(n_804), .B(n_890), .Y(n_891) );
AND2x2_ASAP7_75t_L g892 ( .A(n_835), .B(n_841), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_881), .B(n_882), .Y(n_893) );
AO21x2_ASAP7_75t_L g894 ( .A1(n_872), .A2(n_873), .B(n_844), .Y(n_894) );
AO21x2_ASAP7_75t_L g895 ( .A1(n_838), .A2(n_849), .B(n_846), .Y(n_895) );
INVx1_ASAP7_75t_L g896 ( .A(n_856), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_834), .B(n_792), .Y(n_897) );
OA21x2_ASAP7_75t_L g898 ( .A1(n_858), .A2(n_865), .B(n_861), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_880), .Y(n_899) );
HB1xp67_ASAP7_75t_L g900 ( .A(n_886), .Y(n_900) );
OA21x2_ASAP7_75t_L g901 ( .A1(n_868), .A2(n_859), .B(n_867), .Y(n_901) );
HB1xp67_ASAP7_75t_L g902 ( .A(n_889), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g903 ( .A1(n_833), .A2(n_879), .B(n_864), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_800), .B(n_806), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_870), .Y(n_905) );
OA21x2_ASAP7_75t_L g906 ( .A1(n_874), .A2(n_885), .B(n_876), .Y(n_906) );
INVx3_ASAP7_75t_L g907 ( .A(n_869), .Y(n_907) );
INVx1_ASAP7_75t_SL g908 ( .A(n_814), .Y(n_908) );
OR2x6_ASAP7_75t_L g909 ( .A(n_840), .B(n_823), .Y(n_909) );
AO21x2_ASAP7_75t_L g910 ( .A1(n_860), .A2(n_857), .B(n_855), .Y(n_910) );
INVx2_ASAP7_75t_SL g911 ( .A(n_880), .Y(n_911) );
AND2x2_ASAP7_75t_L g912 ( .A(n_796), .B(n_875), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_887), .Y(n_913) );
INVxp67_ASAP7_75t_L g914 ( .A(n_791), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_878), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_812), .B(n_877), .Y(n_916) );
AO21x2_ASAP7_75t_L g917 ( .A1(n_836), .A2(n_853), .B(n_801), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_798), .B(n_837), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_813), .Y(n_919) );
AOI21xp5_ASAP7_75t_SL g920 ( .A1(n_795), .A2(n_788), .B(n_827), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_815), .Y(n_921) );
AO21x2_ASAP7_75t_L g922 ( .A1(n_836), .A2(n_853), .B(n_801), .Y(n_922) );
AO21x2_ASAP7_75t_L g923 ( .A1(n_821), .A2(n_843), .B(n_850), .Y(n_923) );
INVx3_ASAP7_75t_L g924 ( .A(n_869), .Y(n_924) );
INVx2_ASAP7_75t_L g925 ( .A(n_883), .Y(n_925) );
INVx3_ASAP7_75t_L g926 ( .A(n_840), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_827), .Y(n_927) );
INVx2_ASAP7_75t_SL g928 ( .A(n_826), .Y(n_928) );
AOI21xp5_ASAP7_75t_SL g929 ( .A1(n_795), .A2(n_805), .B(n_829), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_883), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_871), .Y(n_931) );
BUFx2_ASAP7_75t_L g932 ( .A(n_805), .Y(n_932) );
AND2x4_ASAP7_75t_L g933 ( .A(n_852), .B(n_817), .Y(n_933) );
AND2x2_ASAP7_75t_L g934 ( .A(n_798), .B(n_848), .Y(n_934) );
OR2x6_ASAP7_75t_L g935 ( .A(n_825), .B(n_820), .Y(n_935) );
INVx2_ASAP7_75t_L g936 ( .A(n_888), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_816), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_816), .Y(n_938) );
INVx3_ASAP7_75t_L g939 ( .A(n_847), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_816), .Y(n_940) );
OR2x2_ASAP7_75t_L g941 ( .A(n_845), .B(n_819), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_854), .Y(n_942) );
AOI33xp33_ASAP7_75t_L g943 ( .A1(n_789), .A2(n_790), .A3(n_799), .B1(n_818), .B2(n_807), .B3(n_808), .Y(n_943) );
OA21x2_ASAP7_75t_L g944 ( .A1(n_793), .A2(n_824), .B(n_832), .Y(n_944) );
OR2x6_ASAP7_75t_L g945 ( .A(n_862), .B(n_851), .Y(n_945) );
AND2x2_ASAP7_75t_L g946 ( .A(n_811), .B(n_831), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_794), .Y(n_947) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_863), .Y(n_948) );
AO21x2_ASAP7_75t_L g949 ( .A1(n_822), .A2(n_866), .B(n_787), .Y(n_949) );
INVx6_ASAP7_75t_SL g950 ( .A(n_828), .Y(n_950) );
OA21x2_ASAP7_75t_L g951 ( .A1(n_810), .A2(n_842), .B(n_809), .Y(n_951) );
AND2x2_ASAP7_75t_L g952 ( .A(n_810), .B(n_842), .Y(n_952) );
AND2x2_ASAP7_75t_L g953 ( .A(n_810), .B(n_839), .Y(n_953) );
INVx2_ASAP7_75t_L g954 ( .A(n_810), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_810), .Y(n_955) );
BUFx12f_ASAP7_75t_L g956 ( .A(n_797), .Y(n_956) );
BUFx2_ASAP7_75t_L g957 ( .A(n_827), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_884), .B(n_556), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_802), .B(n_803), .Y(n_959) );
INVxp67_ASAP7_75t_SL g960 ( .A(n_830), .Y(n_960) );
AND2x4_ASAP7_75t_L g961 ( .A(n_805), .B(n_827), .Y(n_961) );
OR2x6_ASAP7_75t_L g962 ( .A(n_804), .B(n_890), .Y(n_962) );
INVx5_ASAP7_75t_SL g963 ( .A(n_804), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_802), .B(n_803), .Y(n_964) );
OR2x6_ASAP7_75t_L g965 ( .A(n_804), .B(n_890), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_838), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_896), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_891), .B(n_962), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_896), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_893), .B(n_904), .Y(n_970) );
NOR2xp33_ASAP7_75t_L g971 ( .A(n_908), .B(n_958), .Y(n_971) );
INVx5_ASAP7_75t_L g972 ( .A(n_961), .Y(n_972) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_900), .Y(n_973) );
INVx3_ASAP7_75t_L g974 ( .A(n_907), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_891), .B(n_962), .Y(n_975) );
NOR2xp67_ASAP7_75t_L g976 ( .A(n_956), .B(n_914), .Y(n_976) );
BUFx12f_ASAP7_75t_L g977 ( .A(n_956), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_965), .B(n_901), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_966), .Y(n_979) );
AND2x2_ASAP7_75t_L g980 ( .A(n_965), .B(n_901), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_897), .B(n_912), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_912), .B(n_918), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_902), .Y(n_983) );
INVx3_ASAP7_75t_L g984 ( .A(n_907), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_901), .B(n_931), .Y(n_985) );
OR2x2_ASAP7_75t_L g986 ( .A(n_942), .B(n_916), .Y(n_986) );
INVxp67_ASAP7_75t_SL g987 ( .A(n_907), .Y(n_987) );
INVx4_ASAP7_75t_L g988 ( .A(n_961), .Y(n_988) );
NAND2x1_ASAP7_75t_L g989 ( .A(n_929), .B(n_920), .Y(n_989) );
NOR2x1_ASAP7_75t_SL g990 ( .A(n_935), .B(n_909), .Y(n_990) );
INVx4_ASAP7_75t_L g991 ( .A(n_961), .Y(n_991) );
OR2x2_ASAP7_75t_L g992 ( .A(n_942), .B(n_916), .Y(n_992) );
NAND2x1p5_ASAP7_75t_L g993 ( .A(n_932), .B(n_924), .Y(n_993) );
INVx3_ASAP7_75t_L g994 ( .A(n_924), .Y(n_994) );
INVx2_ASAP7_75t_SL g995 ( .A(n_933), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_959), .B(n_964), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_964), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_898), .Y(n_998) );
INVx4_ASAP7_75t_L g999 ( .A(n_932), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_898), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_963), .B(n_934), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_923), .B(n_917), .Y(n_1002) );
OR2x6_ASAP7_75t_L g1003 ( .A(n_935), .B(n_920), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_963), .B(n_941), .Y(n_1004) );
NAND2x1p5_ASAP7_75t_SL g1005 ( .A(n_946), .B(n_952), .Y(n_1005) );
AND2x2_ASAP7_75t_L g1006 ( .A(n_923), .B(n_917), .Y(n_1006) );
INVx3_ASAP7_75t_L g1007 ( .A(n_924), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1008 ( .A(n_917), .B(n_922), .Y(n_1008) );
NAND2x1p5_ASAP7_75t_SL g1009 ( .A(n_946), .B(n_952), .Y(n_1009) );
AND2x4_ASAP7_75t_L g1010 ( .A(n_905), .B(n_919), .Y(n_1010) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_933), .Y(n_1011) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_905), .B(n_919), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_922), .B(n_937), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_895), .Y(n_1014) );
AND2x2_ASAP7_75t_L g1015 ( .A(n_922), .B(n_937), .Y(n_1015) );
INVx1_ASAP7_75t_SL g1016 ( .A(n_950), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_938), .B(n_940), .Y(n_1017) );
NAND4xp25_ASAP7_75t_L g1018 ( .A(n_943), .B(n_892), .C(n_941), .D(n_903), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_938), .B(n_940), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_921), .B(n_892), .Y(n_1020) );
HB1xp67_ASAP7_75t_L g1021 ( .A(n_960), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g1022 ( .A(n_955), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1023 ( .A(n_963), .B(n_895), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_921), .B(n_895), .Y(n_1024) );
NOR2xp67_ASAP7_75t_L g1025 ( .A(n_899), .B(n_911), .Y(n_1025) );
NAND2x1_ASAP7_75t_L g1026 ( .A(n_935), .B(n_954), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_913), .B(n_894), .Y(n_1027) );
AND2x4_ASAP7_75t_L g1028 ( .A(n_990), .B(n_925), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_1021), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_967), .Y(n_1030) );
INVx2_ASAP7_75t_SL g1031 ( .A(n_999), .Y(n_1031) );
NOR2x1p5_ASAP7_75t_L g1032 ( .A(n_989), .B(n_926), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_986), .B(n_894), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_969), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_985), .B(n_936), .Y(n_1035) );
INVx3_ASAP7_75t_L g1036 ( .A(n_989), .Y(n_1036) );
NOR2x1p5_ASAP7_75t_L g1037 ( .A(n_1026), .B(n_926), .Y(n_1037) );
NAND2xp5_ASAP7_75t_L g1038 ( .A(n_996), .B(n_899), .Y(n_1038) );
OR2x2_ASAP7_75t_L g1039 ( .A(n_992), .B(n_906), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_979), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_985), .B(n_936), .Y(n_1041) );
AOI221x1_ASAP7_75t_L g1042 ( .A1(n_1018), .A2(n_947), .B1(n_926), .B2(n_948), .C(n_954), .Y(n_1042) );
NOR2xp33_ASAP7_75t_L g1043 ( .A(n_971), .B(n_928), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_978), .B(n_915), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_980), .B(n_915), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_980), .B(n_930), .Y(n_1046) );
NOR2xp33_ASAP7_75t_R g1047 ( .A(n_977), .B(n_950), .Y(n_1047) );
NAND2x1_ASAP7_75t_L g1048 ( .A(n_1003), .B(n_951), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_1024), .B(n_1013), .Y(n_1049) );
INVxp33_ASAP7_75t_L g1050 ( .A(n_976), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1015), .B(n_906), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1052 ( .A(n_1017), .B(n_910), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1019), .B(n_910), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1019), .B(n_910), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_998), .Y(n_1055) );
HB1xp67_ASAP7_75t_L g1056 ( .A(n_973), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_983), .Y(n_1057) );
INVx6_ASAP7_75t_L g1058 ( .A(n_972), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_981), .B(n_951), .Y(n_1059) );
OR2x2_ASAP7_75t_L g1060 ( .A(n_982), .B(n_951), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1000), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_997), .B(n_949), .Y(n_1062) );
AND2x4_ASAP7_75t_L g1063 ( .A(n_1003), .B(n_948), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1049), .B(n_968), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1029), .B(n_1020), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1049), .B(n_975), .Y(n_1066) );
INVx1_ASAP7_75t_SL g1067 ( .A(n_1047), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_1055), .Y(n_1068) );
OR2x2_ASAP7_75t_L g1069 ( .A(n_1039), .B(n_970), .Y(n_1069) );
CKINVDCx16_ASAP7_75t_R g1070 ( .A(n_1043), .Y(n_1070) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_1050), .B(n_977), .Y(n_1071) );
NOR2x1_ASAP7_75t_SL g1072 ( .A(n_1031), .B(n_999), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_1056), .Y(n_1073) );
NOR2xp33_ASAP7_75t_L g1074 ( .A(n_1057), .B(n_1016), .Y(n_1074) );
AND2x4_ASAP7_75t_L g1075 ( .A(n_1028), .B(n_1003), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_1044), .B(n_1027), .Y(n_1076) );
INVx2_ASAP7_75t_SL g1077 ( .A(n_1031), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1061), .Y(n_1078) );
OR2x6_ASAP7_75t_L g1079 ( .A(n_1048), .B(n_1003), .Y(n_1079) );
AND2x2_ASAP7_75t_L g1080 ( .A(n_1045), .B(n_1002), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1030), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1046), .B(n_1006), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1039), .B(n_1005), .Y(n_1083) );
NAND2x1_ASAP7_75t_SL g1084 ( .A(n_1036), .B(n_999), .Y(n_1084) );
NAND3x1_ASAP7_75t_L g1085 ( .A(n_1036), .B(n_1008), .C(n_953), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1034), .Y(n_1086) );
OAI22xp33_ASAP7_75t_SL g1087 ( .A1(n_1070), .A2(n_1058), .B1(n_1048), .B2(n_993), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1069), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1089 ( .A(n_1069), .B(n_1059), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1073), .Y(n_1090) );
OR2x2_ASAP7_75t_L g1091 ( .A(n_1065), .B(n_1059), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_1080), .B(n_1051), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_1080), .B(n_1051), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_1082), .B(n_1035), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1083), .B(n_1033), .Y(n_1095) );
INVxp67_ASAP7_75t_SL g1096 ( .A(n_1072), .Y(n_1096) );
AOI21xp5_ASAP7_75t_L g1097 ( .A1(n_1072), .A2(n_987), .B(n_1042), .Y(n_1097) );
NAND2xp5_ASAP7_75t_SL g1098 ( .A(n_1077), .B(n_1036), .Y(n_1098) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1068), .Y(n_1099) );
AOI22x1_ASAP7_75t_L g1100 ( .A1(n_1067), .A2(n_991), .B1(n_988), .B2(n_957), .Y(n_1100) );
INVx1_ASAP7_75t_SL g1101 ( .A(n_1077), .Y(n_1101) );
OAI21xp5_ASAP7_75t_L g1102 ( .A1(n_1085), .A2(n_1025), .B(n_1042), .Y(n_1102) );
O2A1O1Ixp33_ASAP7_75t_L g1103 ( .A1(n_1074), .A2(n_1004), .B(n_1038), .C(n_1001), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1083), .B(n_1060), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1076), .B(n_1041), .Y(n_1105) );
INVx2_ASAP7_75t_SL g1106 ( .A(n_1084), .Y(n_1106) );
AOI21xp33_ASAP7_75t_L g1107 ( .A1(n_1071), .A2(n_1023), .B(n_1062), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1092), .B(n_1064), .Y(n_1108) );
OR3x1_ASAP7_75t_L g1109 ( .A(n_1107), .B(n_1079), .C(n_1040), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1104), .Y(n_1110) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_1096), .A2(n_1079), .B1(n_1058), .B2(n_972), .Y(n_1111) );
NOR3xp33_ASAP7_75t_L g1112 ( .A(n_1102), .B(n_1087), .C(n_1090), .Y(n_1112) );
NAND3xp33_ASAP7_75t_SL g1113 ( .A(n_1101), .B(n_993), .C(n_957), .Y(n_1113) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1089), .Y(n_1114) );
INVx2_ASAP7_75t_L g1115 ( .A(n_1099), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1088), .B(n_1066), .Y(n_1116) );
NAND2xp5_ASAP7_75t_L g1117 ( .A(n_1104), .B(n_1066), .Y(n_1117) );
BUFx6f_ASAP7_75t_L g1118 ( .A(n_1106), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1091), .Y(n_1119) );
AND2x4_ASAP7_75t_L g1120 ( .A(n_1098), .B(n_1079), .Y(n_1120) );
NAND2xp5_ASAP7_75t_SL g1121 ( .A(n_1100), .B(n_1075), .Y(n_1121) );
AOI21xp5_ASAP7_75t_L g1122 ( .A1(n_1121), .A2(n_1098), .B(n_1097), .Y(n_1122) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_1112), .B(n_1095), .C(n_1103), .Y(n_1123) );
NOR2xp67_ASAP7_75t_L g1124 ( .A(n_1121), .B(n_1093), .Y(n_1124) );
HB1xp67_ASAP7_75t_L g1125 ( .A(n_1110), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1119), .Y(n_1126) );
OAI21xp33_ASAP7_75t_SL g1127 ( .A1(n_1108), .A2(n_1105), .B(n_1094), .Y(n_1127) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_1127), .A2(n_1113), .B1(n_1118), .B2(n_1114), .C(n_1117), .Y(n_1128) );
AOI221xp5_ASAP7_75t_L g1129 ( .A1(n_1123), .A2(n_1109), .B1(n_1120), .B2(n_1111), .C(n_1116), .Y(n_1129) );
AOI211xp5_ASAP7_75t_L g1130 ( .A1(n_1124), .A2(n_1120), .B(n_1118), .C(n_927), .Y(n_1130) );
NAND3xp33_ASAP7_75t_L g1131 ( .A(n_1122), .B(n_1118), .C(n_1115), .Y(n_1131) );
NOR2xp33_ASAP7_75t_R g1132 ( .A(n_1126), .B(n_950), .Y(n_1132) );
AOI22x1_ASAP7_75t_L g1133 ( .A1(n_1125), .A2(n_988), .B1(n_991), .B2(n_1032), .Y(n_1133) );
OR5x1_ASAP7_75t_L g1134 ( .A(n_1128), .B(n_1009), .C(n_972), .D(n_988), .E(n_1037), .Y(n_1134) );
NAND5xp2_ASAP7_75t_L g1135 ( .A(n_1129), .B(n_1014), .C(n_1052), .D(n_1053), .E(n_1054), .Y(n_1135) );
NAND4xp25_ASAP7_75t_L g1136 ( .A(n_1130), .B(n_1063), .C(n_1010), .D(n_1012), .Y(n_1136) );
NOR3x1_ASAP7_75t_L g1137 ( .A(n_1131), .B(n_1026), .C(n_1011), .Y(n_1137) );
NOR5xp2_ASAP7_75t_L g1138 ( .A(n_1132), .B(n_1014), .C(n_1078), .D(n_1086), .E(n_1022), .Y(n_1138) );
INVxp67_ASAP7_75t_L g1139 ( .A(n_1135), .Y(n_1139) );
XNOR2xp5_ASAP7_75t_L g1140 ( .A(n_1134), .B(n_1133), .Y(n_1140) );
NOR3xp33_ASAP7_75t_SL g1141 ( .A(n_1136), .B(n_1086), .C(n_1081), .Y(n_1141) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1140), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_1141), .B(n_1137), .Y(n_1143) );
AOI22x1_ASAP7_75t_L g1144 ( .A1(n_1139), .A2(n_1138), .B1(n_1037), .B2(n_1012), .Y(n_1144) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_1142), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1144), .Y(n_1146) );
AOI21xp5_ASAP7_75t_L g1147 ( .A1(n_1146), .A2(n_1143), .B(n_909), .Y(n_1147) );
AOI22xp5_ASAP7_75t_L g1148 ( .A1(n_1145), .A2(n_995), .B1(n_909), .B2(n_1063), .Y(n_1148) );
XNOR2xp5_ASAP7_75t_L g1149 ( .A(n_1147), .B(n_944), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1150 ( .A1(n_1148), .A2(n_984), .B1(n_994), .B2(n_1007), .C(n_974), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1149), .Y(n_1151) );
OAI21xp5_ASAP7_75t_L g1152 ( .A1(n_1151), .A2(n_1150), .B(n_945), .Y(n_1152) );
AOI21xp5_ASAP7_75t_L g1153 ( .A1(n_1152), .A2(n_945), .B(n_939), .Y(n_1153) );
endmodule