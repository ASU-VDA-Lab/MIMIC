module fake_netlist_6_50_n_5792 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_695, n_507, n_580, n_209, n_367, n_465, n_680, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_694, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_676, n_327, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_532, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_689, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_692, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_675, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_681, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_5792);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_680;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_694;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_675;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_681;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_5792;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_1351;
wire n_5254;
wire n_1212;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_3849;
wire n_5138;
wire n_4395;
wire n_4388;
wire n_1061;
wire n_3089;
wire n_783;
wire n_5653;
wire n_4978;
wire n_5409;
wire n_5301;
wire n_1854;
wire n_3088;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_2317;
wire n_5524;
wire n_5345;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_2179;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_5267;
wire n_4249;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_3030;
wire n_830;
wire n_5725;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_2926;
wire n_1078;
wire n_4273;
wire n_5545;
wire n_2321;
wire n_2019;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_4724;
wire n_945;
wire n_5598;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_4696;
wire n_4347;
wire n_5259;
wire n_2480;
wire n_3877;
wire n_3929;
wire n_3048;
wire n_1455;
wire n_5279;
wire n_2786;
wire n_5239;
wire n_1781;
wire n_1971;
wire n_5354;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_3107;
wire n_4956;
wire n_1421;
wire n_3664;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_3047;
wire n_4414;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_2843;
wire n_3760;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_1894;
wire n_3347;
wire n_5136;
wire n_907;
wire n_5638;
wire n_4110;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_2011;
wire n_5684;
wire n_5729;
wire n_5680;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_4671;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_4314;
wire n_2080;
wire n_5099;
wire n_1381;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_2770;
wire n_2101;
wire n_4507;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_3900;
wire n_3488;
wire n_939;
wire n_3732;
wire n_2811;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_1910;
wire n_3980;
wire n_1075;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_3859;
wire n_2692;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_3575;
wire n_2469;
wire n_3927;
wire n_5452;
wire n_3888;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_733;
wire n_2922;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_4331;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_4375;
wire n_1701;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_5532;
wire n_1726;
wire n_4613;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_2641;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_5046;
wire n_2749;
wire n_3298;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_1747;
wire n_5667;
wire n_780;
wire n_2624;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_2092;
wire n_1654;
wire n_1750;
wire n_1462;
wire n_2514;
wire n_5314;
wire n_1588;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_5144;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_3434;
wire n_4510;
wire n_4473;
wire n_5552;
wire n_5226;
wire n_890;
wire n_5457;
wire n_2812;
wire n_4518;
wire n_1709;
wire n_2393;
wire n_2657;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_760;
wire n_1546;
wire n_4394;
wire n_2279;
wire n_1296;
wire n_3352;
wire n_3073;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_1779;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_3021;
wire n_2558;
wire n_1164;
wire n_4697;
wire n_4289;
wire n_4288;
wire n_3763;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_1487;
wire n_3614;
wire n_874;
wire n_5183;
wire n_2145;
wire n_898;
wire n_4964;
wire n_4228;
wire n_3423;
wire n_925;
wire n_1932;
wire n_1101;
wire n_4636;
wire n_4322;
wire n_3644;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_963;
wire n_2767;
wire n_4576;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_4345;
wire n_996;
wire n_1376;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_977;
wire n_3158;
wire n_1788;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_1835;
wire n_3470;
wire n_5076;
wire n_4713;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_3700;
wire n_4995;
wire n_3166;
wire n_3104;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_4310;
wire n_1432;
wire n_5212;
wire n_989;
wire n_2689;
wire n_1473;
wire n_5286;
wire n_2191;
wire n_1246;
wire n_4528;
wire n_899;
wire n_1035;
wire n_4914;
wire n_4939;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_3631;
wire n_5599;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_2103;
wire n_3770;
wire n_2772;
wire n_4440;
wire n_4402;
wire n_927;
wire n_5052;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_4551;
wire n_2857;
wire n_5326;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_3342;
wire n_998;
wire n_5035;
wire n_717;
wire n_1383;
wire n_3390;
wire n_3656;
wire n_1424;
wire n_1000;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_2199;
wire n_2661;
wire n_731;
wire n_5359;
wire n_1955;
wire n_931;
wire n_1791;
wire n_958;
wire n_5137;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_5741;
wire n_2773;
wire n_5405;
wire n_5288;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_2788;
wire n_964;
wire n_4756;
wire n_2797;
wire n_4746;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_2331;
wire n_2292;
wire n_3441;
wire n_3534;
wire n_3964;
wire n_2416;
wire n_1877;
wire n_3944;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_2209;
wire n_3605;
wire n_1602;
wire n_4633;
wire n_3306;
wire n_3026;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_4428;
wire n_1533;
wire n_3323;
wire n_2274;
wire n_5761;
wire n_4618;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_4805;
wire n_1679;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_2146;
wire n_2131;
wire n_5472;
wire n_3547;
wire n_5679;
wire n_2575;
wire n_5100;
wire n_4410;
wire n_1933;
wire n_1179;
wire n_3816;
wire n_4807;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_2928;
wire n_5166;
wire n_1917;
wire n_1580;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_5740;
wire n_1731;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_858;
wire n_2049;
wire n_5182;
wire n_956;
wire n_5534;
wire n_4880;
wire n_3566;
wire n_2781;
wire n_4126;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_1594;
wire n_1869;
wire n_3804;
wire n_4207;
wire n_5196;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_4028;
wire n_2448;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_3406;
wire n_820;
wire n_951;
wire n_952;
wire n_3919;
wire n_2263;
wire n_5185;
wire n_974;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_1934;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_3973;
wire n_2756;
wire n_5334;
wire n_807;
wire n_4761;
wire n_1275;
wire n_2884;
wire n_1510;
wire n_5783;
wire n_3120;
wire n_3797;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_1749;
wire n_3474;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_5556;
wire n_4932;
wire n_5456;
wire n_2302;
wire n_1667;
wire n_1037;
wire n_5143;
wire n_3592;
wire n_5500;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_3967;
wire n_3195;
wire n_2526;
wire n_4274;
wire n_5215;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_4189;
wire n_3817;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_3648;
wire n_1686;
wire n_3042;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_5433;
wire n_3228;
wire n_3657;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_5618;
wire n_1586;
wire n_2264;
wire n_3464;
wire n_3723;
wire n_1190;
wire n_4380;
wire n_4990;
wire n_4996;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_5082;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_5689;
wire n_1043;
wire n_4090;
wire n_4165;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_4144;
wire n_2964;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1361;
wire n_3262;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_937;
wire n_4689;
wire n_1682;
wire n_4547;
wire n_5731;
wire n_3329;
wire n_3826;
wire n_4905;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_1186;
wire n_4623;
wire n_5007;
wire n_3320;
wire n_2518;
wire n_5754;
wire n_3988;
wire n_1720;
wire n_3476;
wire n_4842;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_2688;
wire n_1845;
wire n_1489;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_4859;
wire n_2626;
wire n_1567;
wire n_4037;
wire n_3562;
wire n_2973;
wire n_5218;
wire n_3665;
wire n_3007;
wire n_3528;
wire n_4571;
wire n_3698;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_4215;
wire n_2154;
wire n_1484;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_1373;
wire n_3958;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_5149;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_1385;
wire n_3713;
wire n_1931;
wire n_2668;
wire n_1257;
wire n_3197;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_3124;
wire n_1741;
wire n_1002;
wire n_1949;
wire n_3759;
wire n_2671;
wire n_4516;
wire n_2715;
wire n_1804;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_1337;
wire n_1477;
wire n_2614;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5607;
wire n_3694;
wire n_2937;
wire n_4789;
wire n_4376;
wire n_1001;
wire n_2241;
wire n_4708;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_4462;
wire n_1716;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_749;
wire n_1824;
wire n_3954;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_5577;
wire n_1255;
wire n_5124;
wire n_3951;
wire n_823;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_4639;
wire n_5413;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_1810;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_814;
wire n_5779;
wire n_1643;
wire n_2020;
wire n_4171;
wire n_3652;
wire n_4023;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_3617;
wire n_2076;
wire n_3567;
wire n_1598;
wire n_4344;
wire n_2935;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_918;
wire n_1114;
wire n_4027;
wire n_763;
wire n_3154;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_4391;
wire n_946;
wire n_1303;
wire n_4095;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_1944;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_3215;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_1561;
wire n_1112;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_1460;
wire n_911;
wire n_5159;
wire n_2862;
wire n_2615;
wire n_4068;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_4166;
wire n_1821;
wire n_1058;
wire n_3378;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3176;
wire n_5541;
wire n_5568;
wire n_2505;
wire n_4817;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_3680;
wire n_5381;
wire n_2408;
wire n_5723;
wire n_3468;
wire n_5045;
wire n_1972;
wire n_4383;
wire n_4491;
wire n_5696;
wire n_4486;
wire n_1816;
wire n_3024;
wire n_4612;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_5163;
wire n_4529;
wire n_3361;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_2723;
wire n_5485;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_4390;
wire n_3096;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_3902;
wire n_4062;
wire n_3295;
wire n_4396;
wire n_1998;
wire n_3101;
wire n_1574;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_3125;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_849;
wire n_4684;
wire n_3116;
wire n_4091;
wire n_1753;
wire n_5027;
wire n_3095;
wire n_2471;
wire n_4412;
wire n_2807;
wire n_1921;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_4148;
wire n_2461;
wire n_4057;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_2308;
wire n_2333;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_5018;
wire n_3815;
wire n_3896;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_4457;
wire n_4093;
wire n_1616;
wire n_1862;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_4482;
wire n_1621;
wire n_2547;
wire n_2415;
wire n_5073;
wire n_827;
wire n_4834;
wire n_4762;
wire n_5581;
wire n_3113;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_4504;
wire n_3844;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_3741;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_5601;
wire n_5784;
wire n_3443;
wire n_4819;
wire n_1209;
wire n_5248;
wire n_1708;
wire n_805;
wire n_2051;
wire n_4370;
wire n_2359;
wire n_5112;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_3668;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_5528;
wire n_4302;
wire n_5111;
wire n_3340;
wire n_5227;
wire n_873;
wire n_3946;
wire n_2989;
wire n_5778;
wire n_3395;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_3275;
wire n_836;
wire n_3678;
wire n_3440;
wire n_2094;
wire n_1511;
wire n_2356;
wire n_1422;
wire n_1772;
wire n_4692;
wire n_3165;
wire n_1119;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_2864;
wire n_4311;
wire n_1180;
wire n_2703;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_3261;
wire n_4187;
wire n_940;
wire n_2058;
wire n_2660;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_4962;
wire n_4563;
wire n_5056;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_3532;
wire n_5716;
wire n_3948;
wire n_2124;
wire n_4619;
wire n_5762;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_3803;
wire n_2085;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_3351;
wire n_808;
wire n_5519;
wire n_4047;
wire n_5753;
wire n_3413;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_3791;
wire n_3164;
wire n_4575;
wire n_699;
wire n_4320;
wire n_3884;
wire n_5436;
wire n_5139;
wire n_757;
wire n_5231;
wire n_2190;
wire n_3438;
wire n_4141;
wire n_5193;
wire n_2850;
wire n_1481;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_3883;
wire n_3728;
wire n_2925;
wire n_4499;
wire n_5195;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_5364;
wire n_3315;
wire n_5533;
wire n_3798;
wire n_788;
wire n_1543;
wire n_1599;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_1873;
wire n_3630;
wire n_3518;
wire n_1866;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_3714;
wire n_2228;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_3099;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_1663;
wire n_4172;
wire n_3403;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_3686;
wire n_4502;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4277;
wire n_4526;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_4319;
wire n_3369;
wire n_3581;
wire n_3069;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_3725;
wire n_3933;
wire n_5554;
wire n_1175;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_4066;
wire n_903;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_816;
wire n_1188;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_2467;
wire n_5549;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_5757;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_2377;
wire n_701;
wire n_950;
wire n_3009;
wire n_3719;
wire n_2525;
wire n_4361;
wire n_5488;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_4367;
wire n_5637;
wire n_1987;
wire n_968;
wire n_2271;
wire n_1008;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_2431;
wire n_2078;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_3450;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_5423;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_3436;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_3240;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_4851;
wire n_3293;
wire n_872;
wire n_3922;
wire n_5204;
wire n_5333;
wire n_847;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_5551;
wire n_3150;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_5257;
wire n_765;
wire n_1492;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_4058;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_5059;
wire n_843;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_3799;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_2675;
wire n_5631;
wire n_3537;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_2119;
wire n_947;
wire n_1117;
wire n_1992;
wire n_5686;
wire n_3223;
wire n_3140;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_1698;
wire n_4100;
wire n_4264;
wire n_3788;
wire n_4891;
wire n_777;
wire n_1299;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_4464;
wire n_4624;
wire n_4818;
wire n_4659;
wire n_3600;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_4339;
wire n_3324;
wire n_2338;
wire n_1178;
wire n_796;
wire n_1195;
wire n_1811;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_1048;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_4937;
wire n_5277;
wire n_3615;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_4976;
wire n_2389;
wire n_2132;
wire n_2892;
wire n_4120;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_3718;
wire n_1787;
wire n_1993;
wire n_2281;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_3909;
wire n_5676;
wire n_1220;
wire n_1893;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_4223;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_5121;
wire n_1286;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_4489;
wire n_4839;
wire n_2596;
wire n_3163;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_1531;
wire n_2828;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_759;
wire n_2724;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_1901;
wire n_3869;
wire n_2556;
wire n_4747;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_4801;
wire n_3260;
wire n_2550;
wire n_3175;
wire n_3736;
wire n_5475;
wire n_4448;
wire n_1096;
wire n_2227;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_2159;
wire n_4386;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_1437;
wire n_4844;
wire n_4438;
wire n_4836;
wire n_5439;
wire n_4955;
wire n_4149;
wire n_4355;
wire n_2276;
wire n_3234;
wire n_2803;
wire n_856;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_1129;
wire n_2181;
wire n_2911;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_3429;
wire n_2379;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1635;
wire n_5431;
wire n_4067;
wire n_4357;
wire n_3462;
wire n_2851;
wire n_4374;
wire n_5132;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_3722;
wire n_4400;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_4024;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_732;
wire n_2983;
wire n_2240;
wire n_2538;
wire n_724;
wire n_3250;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_1871;
wire n_4860;
wire n_845;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_768;
wire n_3651;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_4488;
wire n_3767;
wire n_2544;
wire n_3550;
wire n_4211;
wire n_1206;
wire n_4016;
wire n_750;
wire n_5508;
wire n_4656;
wire n_3839;
wire n_2823;
wire n_5597;
wire n_4915;
wire n_4328;
wire n_1057;
wire n_2785;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_1298;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_1589;
wire n_4712;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_3672;
wire n_5318;
wire n_3533;
wire n_1622;
wire n_4725;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_5053;
wire n_2171;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_4109;
wire n_4192;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_5150;
wire n_782;
wire n_809;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_1870;
wire n_1171;
wire n_5179;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_1152;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5585;
wire n_711;
wire n_3105;
wire n_2872;
wire n_3692;
wire n_4616;
wire n_4982;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_2738;
wire n_972;
wire n_5348;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_2346;
wire n_4831;
wire n_3045;
wire n_3821;
wire n_936;
wire n_885;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_3676;
wire n_4896;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_2940;
wire n_4739;
wire n_1974;
wire n_4122;
wire n_934;
wire n_4209;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_5461;
wire n_3003;
wire n_4128;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_1355;
wire n_2258;
wire n_5503;
wire n_804;
wire n_2390;
wire n_959;
wire n_2562;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_5600;
wire n_5755;
wire n_707;
wire n_1900;
wire n_5048;
wire n_3246;
wire n_3381;
wire n_1548;
wire n_1155;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_4715;
wire n_4935;
wire n_4694;
wire n_4672;
wire n_5054;
wire n_2962;
wire n_5448;
wire n_2939;
wire n_5749;
wire n_1672;
wire n_1925;
wire n_4407;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_3258;
wire n_4524;
wire n_3143;
wire n_4084;
wire n_3149;
wire n_3365;
wire n_3379;
wire n_4850;
wire n_4424;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_3939;
wire n_4776;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_1650;
wire n_3506;
wire n_1962;
wire n_3855;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_4723;
wire n_4269;
wire n_5418;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_1019;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_4719;
wire n_5173;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_4735;
wire n_3602;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_2827;
wire n_1177;
wire n_3515;
wire n_1150;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_3806;
wire n_5514;
wire n_2931;
wire n_2569;
wire n_3866;
wire n_5351;
wire n_4543;
wire n_740;
wire n_703;
wire n_4157;
wire n_4229;
wire n_5293;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_1401;
wire n_1516;
wire n_3846;
wire n_3512;
wire n_5201;
wire n_2029;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_832;
wire n_3049;
wire n_5389;
wire n_5142;
wire n_3830;
wire n_3679;
wire n_3541;
wire n_3117;
wire n_4930;
wire n_5623;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_2149;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_895;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_4416;
wire n_4593;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_5114;
wire n_4980;
wire n_1392;
wire n_5693;
wire n_4495;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_2463;
wire n_3363;
wire n_1677;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_4559;
wire n_838;
wire n_3969;
wire n_3336;
wire n_4160;
wire n_4231;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_5203;
wire n_930;
wire n_2620;
wire n_5162;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_1414;
wire n_5285;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_2683;
wire n_5365;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_990;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_870;
wire n_5395;
wire n_1253;
wire n_5709;
wire n_1693;
wire n_3802;
wire n_3256;
wire n_2118;
wire n_2111;
wire n_2915;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_2802;
wire n_3643;
wire n_2425;
wire n_4265;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_3060;
wire n_3098;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_4064;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_5266;
wire n_5580;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_1789;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_3863;
wire n_3669;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_5764;
wire n_2282;
wire n_4628;
wire n_2047;
wire n_5385;
wire n_1609;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_1763;
wire n_5322;
wire n_3989;
wire n_2490;
wire n_4460;
wire n_4108;
wire n_3786;
wire n_3841;
wire n_4254;
wire n_1996;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_1158;
wire n_2248;
wire n_5011;
wire n_3147;
wire n_2662;
wire n_4909;
wire n_753;
wire n_3925;
wire n_3180;
wire n_2795;
wire n_3472;
wire n_5376;
wire n_5106;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_3717;
wire n_5561;
wire n_5410;
wire n_2215;
wire n_1884;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_2038;
wire n_4447;
wire n_4826;
wire n_3445;
wire n_1833;
wire n_3903;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_5378;
wire n_1417;
wire n_3673;
wire n_4281;
wire n_4648;
wire n_3094;
wire n_965;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_4957;
wire n_3079;
wire n_4360;
wire n_4039;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_4853;
wire n_1748;
wire n_3504;
wire n_4272;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_3111;
wire n_1885;
wire n_5269;
wire n_3054;
wire n_1538;
wire n_1240;
wire n_5468;
wire n_4730;
wire n_5399;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_2353;
wire n_4099;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_5550;
wire n_3911;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_2997;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5509;
wire n_5382;
wire n_5659;
wire n_3619;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_4065;
wire n_2645;
wire n_3904;
wire n_1393;
wire n_1867;
wire n_1517;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_4733;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_1056;
wire n_758;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_4879;
wire n_772;
wire n_2806;
wire n_770;
wire n_3028;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_886;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_4117;
wire n_4687;
wire n_2836;
wire n_1404;
wire n_5492;
wire n_2378;
wire n_887;
wire n_2655;
wire n_4600;
wire n_1467;
wire n_4250;
wire n_3906;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_3963;
wire n_3368;
wire n_2370;
wire n_2612;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_913;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_5525;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_4305;
wire n_824;
wire n_4297;
wire n_2907;
wire n_5374;
wire n_5575;
wire n_1843;
wire n_5675;
wire n_4227;
wire n_2778;
wire n_1909;
wire n_5020;
wire n_5297;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_1970;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_4364;
wire n_1957;
wire n_4354;
wire n_4732;
wire n_3912;
wire n_3118;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_860;
wire n_1530;
wire n_4745;
wire n_938;
wire n_1302;
wire n_5642;
wire n_4581;
wire n_4377;
wire n_2143;
wire n_905;
wire n_4792;
wire n_1680;
wire n_3842;
wire n_993;
wire n_2031;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_2654;
wire n_3036;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_2711;
wire n_4199;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_1312;
wire n_5668;
wire n_5038;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_5463;
wire n_3022;
wire n_5489;
wire n_1165;
wire n_4773;
wire n_5654;
wire n_2008;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_1386;
wire n_4427;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_2804;
wire n_2453;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_4822;
wire n_1214;
wire n_850;
wire n_5692;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_825;
wire n_3785;
wire n_2963;
wire n_5366;
wire n_2602;
wire n_3873;
wire n_2980;
wire n_4886;
wire n_1317;
wire n_1082;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_4055;
wire n_2178;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_1796;
wire n_2082;
wire n_3519;
wire n_5078;
wire n_3707;
wire n_3578;
wire n_909;
wire n_4737;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_2943;
wire n_5205;
wire n_1634;
wire n_3252;
wire n_3253;
wire n_1465;
wire n_2622;
wire n_2658;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_4603;
wire n_1523;
wire n_1627;
wire n_5080;
wire n_3128;
wire n_1527;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_2230;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_1565;
wire n_1493;
wire n_5690;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_1514;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_4994;
wire n_2537;
wire n_4483;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_3171;
wire n_3608;
wire n_4540;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_3499;
wire n_4284;
wire n_1005;
wire n_1947;
wire n_3426;
wire n_4971;
wire n_5656;
wire n_1469;
wire n_5125;
wire n_2650;
wire n_5652;
wire n_987;
wire n_5499;
wire n_720;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_738;
wire n_2012;
wire n_3497;
wire n_5066;
wire n_3580;
wire n_2842;
wire n_2335;
wire n_2307;
wire n_3704;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_4280;
wire n_1181;
wire n_5190;
wire n_3173;
wire n_3677;
wire n_3996;
wire n_1049;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_2868;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_5442;
wire n_4459;
wire n_4545;
wire n_2896;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_5295;
wire n_2368;
wire n_4175;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_1073;
wire n_4514;
wire n_3191;
wire n_5584;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_2682;
wire n_3032;
wire n_5160;
wire n_2877;
wire n_5098;
wire n_1021;
wire n_811;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_5497;
wire n_880;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_2432;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3641;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_1382;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_2701;
wire n_2511;
wire n_4167;
wire n_1427;
wire n_2745;
wire n_1080;
wire n_5271;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_5234;
wire n_4431;
wire n_2421;
wire n_1136;
wire n_4387;
wire n_2618;
wire n_3265;
wire n_2464;
wire n_3755;
wire n_4042;
wire n_1125;
wire n_5128;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_5467;
wire n_4299;
wire n_4890;
wire n_1784;
wire n_3571;
wire n_1775;
wire n_2410;
wire n_1093;
wire n_1783;
wire n_2929;
wire n_4176;
wire n_5199;
wire n_3407;
wire n_5313;
wire n_3856;
wire n_4236;
wire n_1185;
wire n_3425;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_5079;
wire n_1453;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3188;
wire n_1459;
wire n_3243;
wire n_2462;
wire n_1135;
wire n_2889;
wire n_4034;
wire n_4056;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_4887;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_906;
wire n_1390;
wire n_2289;
wire n_1733;
wire n_2955;
wire n_5592;
wire n_2158;
wire n_4609;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_736;
wire n_5278;
wire n_3525;
wire n_3314;
wire n_2100;
wire n_5157;
wire n_3016;
wire n_4754;
wire n_2993;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_4003;
wire n_5708;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_1905;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_5287;
wire n_1079;
wire n_2139;
wire n_5083;
wire n_4509;
wire n_2875;
wire n_3907;
wire n_1103;
wire n_3338;
wire n_4217;
wire n_4906;
wire n_2219;
wire n_1203;
wire n_3636;
wire n_2327;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_4897;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_3572;
wire n_3886;
wire n_4710;
wire n_4420;
wire n_892;
wire n_3637;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_1718;
wire n_5174;
wire n_4234;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_1847;
wire n_3634;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_4945;
wire n_3417;
wire n_5677;
wire n_4124;
wire n_5570;
wire n_785;
wire n_5153;
wire n_4611;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_2607;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_3249;
wire n_1320;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_5486;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_4832;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_5391;
wire n_1938;
wire n_2472;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_4554;
wire n_3040;
wire n_3279;
wire n_5240;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1692;
wire n_1084;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3501;
wire n_3475;
wire n_1705;
wire n_3905;
wire n_4680;
wire n_3013;
wire n_921;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_2200;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_3878;
wire n_2670;
wire n_2700;
wire n_1041;
wire n_3134;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_896;
wire n_4553;
wire n_3278;
wire n_2084;
wire n_4875;
wire n_5682;
wire n_5387;
wire n_5557;
wire n_2458;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_4321;
wire n_4183;
wire n_5681;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4821;
wire n_4145;
wire n_3121;
wire n_4040;
wire n_1640;
wire n_2406;
wire n_806;
wire n_2141;
wire n_5316;
wire n_5703;
wire n_833;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_2561;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_1241;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_4338;
wire n_3457;
wire n_3762;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_3558;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_4726;
wire n_1045;
wire n_786;
wire n_1559;
wire n_1872;
wire n_5040;
wire n_1325;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_1727;
wire n_4301;
wire n_3744;
wire n_4788;
wire n_2041;
wire n_1360;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_3543;
wire n_3621;
wire n_2903;
wire n_3216;
wire n_3808;
wire n_4365;
wire n_1882;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_3758;
wire n_5417;
wire n_2587;
wire n_3199;
wire n_3339;
wire n_4923;
wire n_2400;
wire n_1953;
wire n_4741;
wire n_3343;
wire n_2752;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_4652;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_2814;
wire n_5253;
wire n_5209;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_4295;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_5777;
wire n_4225;
wire n_747;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_5064;
wire n_5610;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_1994;
wire n_957;
wire n_2566;
wire n_744;
wire n_971;
wire n_2702;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_4568;
wire n_1205;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_5786;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_1016;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_1083;
wire n_5768;
wire n_3553;
wire n_2465;
wire n_2275;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_1721;
wire n_3494;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_4409;
wire n_4629;
wire n_4638;
wire n_708;
wire n_1973;
wire n_3181;
wire n_5700;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_904;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3328;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_2466;
wire n_2530;
wire n_1085;
wire n_2042;
wire n_771;
wire n_924;
wire n_1582;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_2035;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_4104;
wire n_4845;
wire n_1770;
wire n_878;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_981;
wire n_4089;
wire n_5478;
wire n_2071;
wire n_1144;
wire n_3219;
wire n_3702;
wire n_2233;
wire n_4779;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_1198;
wire n_4061;
wire n_2174;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_1133;
wire n_4429;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_4865;
wire n_1039;
wire n_2043;
wire n_1480;
wire n_3206;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_4562;
wire n_3383;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_4186;
wire n_2540;
wire n_973;
wire n_5743;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_2065;
wire n_2879;
wire n_967;
wire n_4522;
wire n_2001;
wire n_4341;
wire n_1629;
wire n_5368;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_3555;
wire n_915;
wire n_812;
wire n_1131;
wire n_3155;
wire n_1006;
wire n_3110;
wire n_1632;
wire n_1888;
wire n_1311;
wire n_4780;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_3467;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_1322;
wire n_1958;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_4984;
wire n_2579;
wire n_2105;
wire n_1423;
wire n_3387;
wire n_5782;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1612;
wire n_4809;
wire n_1199;
wire n_3392;
wire n_3773;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_798;
wire n_2324;
wire n_5563;
wire n_1348;
wire n_2977;
wire n_1739;
wire n_1380;
wire n_2847;
wire n_2557;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_2647;
wire n_883;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_2521;
wire n_1099;
wire n_4578;
wire n_2211;
wire n_4777;
wire n_5720;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_1285;
wire n_1985;
wire n_1172;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_3031;
wire n_4029;
wire n_2447;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_1649;
wire n_4555;
wire n_5650;
wire n_4969;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_822;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_2212;
wire n_3063;
wire n_2729;
wire n_1163;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_3998;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_3655;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_2108;
wire n_5158;
wire n_1211;
wire n_5022;
wire n_5670;
wire n_1280;
wire n_3296;
wire n_5276;
wire n_1445;
wire n_2551;
wire n_1526;
wire n_5047;
wire n_2985;
wire n_1978;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_4403;
wire n_5238;
wire n_3269;
wire n_3531;
wire n_1054;
wire n_1956;
wire n_4139;
wire n_4549;
wire n_1986;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_5429;
wire n_813;
wire n_3822;
wire n_4163;
wire n_818;
wire n_5535;
wire n_3812;
wire n_3910;
wire n_2633;
wire n_2207;
wire n_4948;
wire n_5268;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_2198;
wire n_3319;
wire n_2073;
wire n_2273;
wire n_3748;
wire n_3272;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_3396;
wire n_4393;
wire n_1162;
wire n_821;
wire n_4372;
wire n_1068;
wire n_982;
wire n_5640;
wire n_932;
wire n_4318;
wire n_2831;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_2123;
wire n_1697;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_2941;
wire n_1278;
wire n_5108;
wire n_4032;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_4147;
wire n_4477;
wire n_3168;
wire n_2751;
wire n_4337;
wire n_4130;
wire n_2009;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_3092;
wire n_1289;
wire n_3055;
wire n_3966;
wire n_2866;
wire n_4742;
wire n_3734;
wire n_1014;
wire n_1703;
wire n_2580;
wire n_882;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_3384;
wire n_1950;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5202;
wire n_702;
wire n_4965;
wire n_3346;
wire n_1896;
wire n_2965;
wire n_3058;
wire n_3861;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_4523;
wire n_1655;
wire n_1886;
wire n_4371;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_3689;
wire n_877;
wire n_4673;
wire n_2519;
wire n_728;
wire n_3415;
wire n_1063;
wire n_4607;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_4169;
wire n_697;
wire n_3271;
wire n_5088;
wire n_4248;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_1825;
wire n_1757;
wire n_1792;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_3993;
wire n_4685;
wire n_4031;
wire n_4675;
wire n_2663;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_2750;
wire n_2775;
wire n_1295;
wire n_3477;
wire n_2349;
wire n_5596;
wire n_2684;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_4653;
wire n_4435;
wire n_5604;
wire n_1756;
wire n_1128;
wire n_5411;
wire n_4019;
wire n_1071;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_4922;
wire n_865;
wire n_3616;
wire n_4191;
wire n_5695;
wire n_2870;
wire n_2151;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_826;
wire n_4350;
wire n_3747;
wire n_1714;
wire n_718;
wire n_5331;
wire n_4330;
wire n_5311;
wire n_2089;
wire n_3522;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_704;
wire n_2148;
wire n_4162;
wire n_5565;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_5520;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_1838;
wire n_2638;
wire n_4785;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_2002;
wire n_2138;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5669;
wire n_5772;
wire n_2208;
wire n_4775;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_1304;
wire n_3775;
wire n_4669;
wire n_2134;
wire n_1176;
wire n_5603;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_2489;
wire n_1087;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_1505;
wire n_5712;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_3620;
wire n_3832;
wire n_2520;
wire n_4484;
wire n_3693;
wire n_4497;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_2251;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_2403;
wire n_1070;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_2589;
wire n_4535;
wire n_755;
wire n_2442;
wire n_3627;
wire n_3480;
wire n_1368;
wire n_1137;
wire n_3612;
wire n_4695;
wire n_2545;
wire n_3509;
wire n_4368;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_1314;
wire n_3196;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_1534;
wire n_5005;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_723;
wire n_3144;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_3640;
wire n_1159;
wire n_3481;
wire n_995;
wire n_2250;
wire n_3033;
wire n_5775;
wire n_2374;
wire n_1681;
wire n_4597;
wire n_3364;
wire n_3226;
wire n_4020;
wire n_2780;
wire n_5220;
wire n_1618;
wire n_4867;
wire n_5061;
wire n_1653;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_2920;
wire n_773;
wire n_920;
wire n_1374;
wire n_2648;
wire n_3212;
wire n_1169;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_4721;
wire n_3093;
wire n_848;
wire n_4247;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_2023;
wire n_2204;
wire n_2720;
wire n_4614;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_4001;
wire n_1323;
wire n_2627;
wire n_4422;
wire n_960;
wire n_778;
wire n_3004;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_5037;
wire n_2515;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_2201;
wire n_725;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_4635;
wire n_994;
wire n_5735;
wire n_2278;
wire n_1020;
wire n_1273;
wire n_4214;
wire n_3448;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_3991;
wire n_3516;
wire n_3926;
wire n_1095;
wire n_1270;
wire n_4405;
wire n_4413;
wire n_1852;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_4667;
wire n_5081;
wire n_4182;
wire n_3230;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_1409;
wire n_5189;
wire n_1503;
wire n_2819;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3635;
wire n_5118;
wire n_4155;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_5632;
wire n_5582;
wire n_5425;
wire n_1216;
wire n_2716;
wire n_2452;
wire n_3650;
wire n_5446;
wire n_3010;
wire n_3043;
wire n_5224;
wire n_4590;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_3529;
wire n_3238;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_2790;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_5437;
wire n_4586;
wire n_1608;
wire n_2373;
wire n_1472;
wire n_3628;
wire n_5454;
wire n_800;
wire n_4734;
wire n_1491;
wire n_1840;
wire n_4434;
wire n_5307;
wire n_2244;
wire n_4290;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_3790;
wire n_2766;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_5230;
wire n_4888;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_2229;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_2099;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_4561;
wire n_4461;
wire n_3245;
wire n_3075;
wire n_4007;
wire n_4949;
wire n_2642;
wire n_4239;
wire n_2383;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_2536;
wire n_3915;
wire n_1633;
wire n_3489;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2727;
wire n_3377;
wire n_4782;
wire n_1321;
wire n_2533;
wire n_3530;
wire n_2869;
wire n_4378;
wire n_5349;
wire n_1235;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_790;
wire n_2901;
wire n_2611;
wire n_4358;
wire n_5616;
wire n_2653;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_4469;
wire n_5169;
wire n_3156;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_743;
wire n_766;
wire n_1746;
wire n_3524;
wire n_2885;
wire n_3097;
wire n_2062;
wire n_4539;
wire n_2975;
wire n_4421;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_1607;
wire n_1454;
wire n_4953;
wire n_2348;
wire n_2944;
wire n_3831;
wire n_869;
wire n_1154;
wire n_1329;
wire n_5167;
wire n_5661;
wire n_3589;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_3391;
wire n_1800;
wire n_1463;
wire n_3458;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_5558;
wire n_1826;
wire n_5687;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_5051;
wire n_5587;
wire n_5236;
wire n_853;
wire n_875;
wire n_5012;
wire n_1678;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5025;
wire n_933;
wire n_4173;
wire n_3135;
wire n_5651;
wire n_4630;
wire n_1217;
wire n_5645;
wire n_3990;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_988;
wire n_2796;
wire n_2507;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_1204;
wire n_1132;
wire n_1327;
wire n_955;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_5412;
wire n_769;
wire n_2380;
wire n_4786;
wire n_1120;
wire n_4579;
wire n_2290;
wire n_4811;
wire n_2048;
wire n_2005;
wire n_4857;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_863;
wire n_3774;
wire n_5733;
wire n_2910;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_2584;
wire n_1812;
wire n_866;
wire n_2287;
wire n_5791;
wire n_5727;
wire n_761;
wire n_2492;
wire n_3778;
wire n_5328;
wire n_5657;
wire n_1173;
wire n_4974;
wire n_4911;
wire n_4436;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_3334;
wire n_5602;
wire n_5097;
wire n_844;
wire n_4985;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_3114;
wire n_2741;
wire n_888;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_4309;
wire n_4363;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_4025;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_4313;
wire n_3309;
wire n_3671;
wire n_4142;
wire n_2015;
wire n_3982;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_3796;
wire n_3840;
wire n_3461;
wire n_3408;
wire n_4246;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_1525;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_4244;
wire n_2147;
wire n_2503;
wire n_4049;
wire n_1156;
wire n_2600;
wire n_984;
wire n_5626;
wire n_3508;
wire n_868;
wire n_4353;
wire n_735;
wire n_4787;
wire n_5633;
wire n_1218;
wire n_5664;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_4351;
wire n_2429;
wire n_985;
wire n_2440;
wire n_3521;
wire n_802;
wire n_980;
wire n_2681;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_4784;
wire n_4075;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_3066;
wire n_2844;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_5280;
wire n_4451;
wire n_4332;
wire n_810;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_3563;
wire n_2367;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_2909;
wire n_754;
wire n_5369;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_3187;
wire n_3218;
wire n_861;
wire n_857;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_2221;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_2709;
wire n_1578;
wire n_1861;
wire n_3955;
wire n_2280;
wire n_1557;
wire n_3945;
wire n_730;
wire n_5214;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_3433;
wire n_4463;
wire n_2185;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_5032;
wire n_1899;
wire n_784;
wire n_4804;
wire n_5619;
wire n_3965;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_1449;
wire n_4703;
wire n_2419;
wire n_5683;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_614),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_361),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_581),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_54),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_381),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_127),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_538),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_155),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_108),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_99),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_605),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_400),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_673),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_48),
.Y(n_710)
);

CKINVDCx20_ASAP7_75t_R g711 ( 
.A(n_95),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_146),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_127),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_180),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_691),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_245),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_104),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_117),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_392),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_380),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_17),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_477),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_560),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_122),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_209),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_251),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_427),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_512),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_617),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_181),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_448),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_348),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_616),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_584),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_453),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_516),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_447),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_277),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_37),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_158),
.Y(n_741)
);

BUFx5_ASAP7_75t_L g742 ( 
.A(n_405),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_184),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_518),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_379),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_426),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_466),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_373),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_568),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_40),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_624),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_350),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_406),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_387),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_81),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_179),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_368),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_345),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_503),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_289),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_496),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_87),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_119),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_237),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_511),
.Y(n_765)
);

CKINVDCx20_ASAP7_75t_R g766 ( 
.A(n_59),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_305),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_37),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_504),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_476),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_550),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_548),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_295),
.Y(n_773)
);

INVx1_ASAP7_75t_SL g774 ( 
.A(n_677),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_480),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_634),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_107),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_276),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_361),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_377),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_155),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_619),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_238),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_428),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_209),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_346),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_550),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_139),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_38),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_413),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_570),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_372),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_404),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_445),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_250),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_206),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_164),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_582),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_38),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_493),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_308),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_606),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_263),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_531),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_664),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_10),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_202),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_108),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_670),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_556),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_692),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_541),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_25),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_218),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_234),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_245),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_456),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_189),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_27),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_322),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_429),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_532),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_650),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_151),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_471),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_680),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_508),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_109),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_322),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_675),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_573),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_586),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_326),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_223),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_522),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_625),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_629),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_74),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_464),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_123),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_234),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_187),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_463),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_177),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_48),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_17),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_620),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_123),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_646),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_197),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_429),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_221),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_204),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_301),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_570),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_58),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_49),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_321),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_167),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_216),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_304),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_229),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_343),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_368),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_350),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_399),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_138),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_274),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_613),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_360),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_169),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_75),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_606),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_194),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_358),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_405),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_167),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_78),
.Y(n_878)
);

BUFx10_ASAP7_75t_L g879 ( 
.A(n_30),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_55),
.Y(n_880)
);

CKINVDCx16_ASAP7_75t_R g881 ( 
.A(n_343),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_365),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_451),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_653),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_467),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_296),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_281),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_288),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_70),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_598),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_336),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_346),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_684),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_434),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_485),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_353),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_256),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_369),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_192),
.Y(n_899)
);

CKINVDCx14_ASAP7_75t_R g900 ( 
.A(n_468),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_626),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_76),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_539),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_410),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_70),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_288),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_221),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_187),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_15),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_359),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_338),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_113),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_461),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_172),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_154),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_239),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_609),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_594),
.Y(n_918)
);

CKINVDCx14_ASAP7_75t_R g919 ( 
.A(n_69),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_390),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_433),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_438),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_422),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_163),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_215),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_609),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_508),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_310),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_480),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_342),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_400),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_217),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_404),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_639),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_307),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_316),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_284),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_587),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_313),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_591),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_378),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_528),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_69),
.Y(n_943)
);

CKINVDCx14_ASAP7_75t_R g944 ( 
.A(n_600),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_611),
.Y(n_945)
);

BUFx10_ASAP7_75t_L g946 ( 
.A(n_473),
.Y(n_946)
);

INVx2_ASAP7_75t_SL g947 ( 
.A(n_243),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_665),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_602),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_95),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_455),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_243),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_342),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_182),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_71),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_205),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_407),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_26),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_184),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_19),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_483),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_555),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_588),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_256),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_135),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_585),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_573),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_600),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_507),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_569),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_42),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_207),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_154),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_43),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_133),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_107),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_479),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_562),
.Y(n_978)
);

BUFx5_ASAP7_75t_L g979 ( 
.A(n_566),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_131),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_527),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_43),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_348),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_128),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_358),
.Y(n_985)
);

CKINVDCx16_ASAP7_75t_R g986 ( 
.A(n_627),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_72),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_274),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_667),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_556),
.Y(n_990)
);

CKINVDCx14_ASAP7_75t_R g991 ( 
.A(n_636),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_260),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_572),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_533),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_196),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_601),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_312),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_79),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_227),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_509),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_507),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_120),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_385),
.Y(n_1003)
);

INVx4_ASAP7_75t_R g1004 ( 
.A(n_169),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_118),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_224),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_359),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_65),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_555),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_185),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_571),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_418),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_540),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_199),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_115),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_60),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_618),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_591),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_483),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_540),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_323),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_604),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_387),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_253),
.Y(n_1024)
);

INVxp33_ASAP7_75t_L g1025 ( 
.A(n_247),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_392),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_397),
.Y(n_1027)
);

CKINVDCx16_ASAP7_75t_R g1028 ( 
.A(n_104),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_233),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_681),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_465),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_551),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_596),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_191),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_55),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_502),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_308),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_485),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_237),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_487),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_59),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_85),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_461),
.Y(n_1043)
);

CKINVDCx16_ASAP7_75t_R g1044 ( 
.A(n_302),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_302),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_688),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_306),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_402),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_385),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_282),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_213),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_134),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_138),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_553),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_463),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_110),
.Y(n_1056)
);

INVxp67_ASAP7_75t_SL g1057 ( 
.A(n_375),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_203),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_102),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_281),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_224),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_603),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_126),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_687),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_225),
.Y(n_1065)
);

INVx1_ASAP7_75t_SL g1066 ( 
.A(n_258),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_89),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_232),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_207),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_332),
.Y(n_1070)
);

CKINVDCx20_ASAP7_75t_R g1071 ( 
.A(n_468),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_170),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_253),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_251),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_538),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_189),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_120),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_496),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_320),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_422),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_439),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_2),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_161),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_445),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_171),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_217),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_2),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_427),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_455),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_62),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_568),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_156),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_524),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_336),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_14),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_92),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_125),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_547),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_644),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_504),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_289),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_165),
.Y(n_1102)
);

BUFx10_ASAP7_75t_L g1103 ( 
.A(n_370),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_226),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_536),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_194),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_402),
.Y(n_1107)
);

CKINVDCx14_ASAP7_75t_R g1108 ( 
.A(n_435),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_484),
.Y(n_1109)
);

BUFx10_ASAP7_75t_L g1110 ( 
.A(n_337),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_451),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_589),
.Y(n_1112)
);

BUFx10_ASAP7_75t_L g1113 ( 
.A(n_669),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_137),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_475),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_142),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_163),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_635),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_401),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_695),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_661),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_103),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_239),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_389),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_457),
.Y(n_1125)
);

BUFx10_ASAP7_75t_L g1126 ( 
.A(n_54),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_535),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_296),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_192),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_659),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_494),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_444),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_204),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_309),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_117),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_474),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_82),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_506),
.Y(n_1138)
);

INVx2_ASAP7_75t_SL g1139 ( 
.A(n_589),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_316),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_211),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_506),
.Y(n_1142)
);

CKINVDCx14_ASAP7_75t_R g1143 ( 
.A(n_539),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_113),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_587),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_112),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_579),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_494),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_306),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_395),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_188),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_135),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_497),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_34),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_206),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_562),
.Y(n_1156)
);

INVxp33_ASAP7_75t_R g1157 ( 
.A(n_247),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_551),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_7),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_517),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_28),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_32),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_263),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_375),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_323),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_185),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_142),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_481),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_501),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_406),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_233),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_655),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_363),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_671),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_486),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_310),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_314),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_5),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_258),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_157),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_132),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_278),
.Y(n_1182)
);

BUFx3_ASAP7_75t_L g1183 ( 
.A(n_131),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_638),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_583),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_548),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_593),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_260),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_219),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_571),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_662),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_102),
.Y(n_1192)
);

CKINVDCx16_ASAP7_75t_R g1193 ( 
.A(n_240),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_376),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_255),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_444),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_502),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_513),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_612),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_533),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_553),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_182),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_190),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_145),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_376),
.Y(n_1205)
);

BUFx10_ASAP7_75t_L g1206 ( 
.A(n_524),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_88),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_352),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_100),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_389),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_203),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_265),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_111),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_41),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_254),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_610),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_300),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_457),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_519),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_447),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_900),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_742),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_742),
.Y(n_1223)
);

INVxp67_ASAP7_75t_L g1224 ( 
.A(n_801),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_742),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_701),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1030),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_742),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_742),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_711),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_742),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_742),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_742),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_730),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_742),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_919),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1030),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_979),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_979),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_713),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1030),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_979),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_944),
.Y(n_1243)
);

INVxp33_ASAP7_75t_SL g1244 ( 
.A(n_740),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_979),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_979),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1108),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_801),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_979),
.Y(n_1249)
);

INVxp67_ASAP7_75t_SL g1250 ( 
.A(n_1179),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_979),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1179),
.Y(n_1252)
);

INVxp33_ASAP7_75t_SL g1253 ( 
.A(n_752),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_979),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_831),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_979),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_729),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_729),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_738),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_809),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_809),
.Y(n_1261)
);

CKINVDCx16_ASAP7_75t_R g1262 ( 
.A(n_831),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1179),
.B(n_0),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_849),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_755),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_849),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_884),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_766),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_884),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1017),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1017),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1120),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1120),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_713),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1121),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1121),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1172),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1172),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1174),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1174),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1179),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_775),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_713),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_714),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_881),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_714),
.Y(n_1286)
);

CKINVDCx16_ASAP7_75t_R g1287 ( 
.A(n_881),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_714),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_731),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_731),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1143),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_731),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_909),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_909),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_909),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_822),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_925),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_925),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1113),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_925),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_751),
.B(n_1),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1001),
.Y(n_1302)
);

CKINVDCx16_ASAP7_75t_R g1303 ( 
.A(n_1001),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_926),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_713),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_926),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_926),
.Y(n_1307)
);

CKINVDCx16_ASAP7_75t_R g1308 ( 
.A(n_1028),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_950),
.Y(n_1309)
);

CKINVDCx14_ASAP7_75t_R g1310 ( 
.A(n_991),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_950),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_950),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_969),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_713),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_969),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_969),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_697),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1029),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_744),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_709),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_847),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_L g1322 ( 
.A(n_822),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_713),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1029),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_776),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1029),
.Y(n_1326)
);

CKINVDCx16_ASAP7_75t_R g1327 ( 
.A(n_1028),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1183),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_782),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_805),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1183),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1183),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_811),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_791),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_823),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_773),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_847),
.Y(n_1337)
);

CKINVDCx14_ASAP7_75t_R g1338 ( 
.A(n_1113),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1189),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1189),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1189),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1207),
.Y(n_1342)
);

CKINVDCx16_ASAP7_75t_R g1343 ( 
.A(n_1044),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1207),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1207),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1216),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1044),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_862),
.B(n_0),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_826),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_862),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1216),
.Y(n_1351)
);

CKINVDCx14_ASAP7_75t_R g1352 ( 
.A(n_1113),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_804),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1216),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_847),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_773),
.Y(n_1356)
);

BUFx2_ASAP7_75t_SL g1357 ( 
.A(n_1184),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1160),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1113),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_773),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_773),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1160),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_773),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_773),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_808),
.Y(n_1365)
);

BUFx5_ASAP7_75t_L g1366 ( 
.A(n_699),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_1193),
.Y(n_1367)
);

INVxp33_ASAP7_75t_SL g1368 ( 
.A(n_763),
.Y(n_1368)
);

INVxp33_ASAP7_75t_L g1369 ( 
.A(n_896),
.Y(n_1369)
);

INVxp33_ASAP7_75t_SL g1370 ( 
.A(n_702),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_920),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_751),
.B(n_830),
.Y(n_1372)
);

BUFx5_ASAP7_75t_L g1373 ( 
.A(n_699),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_920),
.Y(n_1374)
);

INVxp33_ASAP7_75t_SL g1375 ( 
.A(n_705),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_920),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_920),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1193),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_726),
.B(n_1),
.Y(n_1379)
);

CKINVDCx16_ASAP7_75t_R g1380 ( 
.A(n_986),
.Y(n_1380)
);

CKINVDCx11_ASAP7_75t_R g1381 ( 
.A(n_744),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_920),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_920),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_999),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_999),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_837),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_869),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_999),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_999),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_708),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_893),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_934),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_700),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_999),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_999),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_1100),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1100),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_948),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1100),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_989),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1100),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1100),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_832),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1100),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1208),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_710),
.Y(n_1406)
);

CKINVDCx14_ASAP7_75t_R g1407 ( 
.A(n_1046),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1208),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_863),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1064),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_874),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1208),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1208),
.Y(n_1413)
);

INVxp67_ASAP7_75t_SL g1414 ( 
.A(n_1208),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1208),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1099),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1212),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1212),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1118),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1212),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1212),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1212),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1130),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_716),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1212),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_719),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1191),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1215),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1215),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1215),
.Y(n_1430)
);

HB1xp67_ASAP7_75t_L g1431 ( 
.A(n_720),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1215),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1199),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1215),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1215),
.Y(n_1435)
);

INVxp67_ASAP7_75t_SL g1436 ( 
.A(n_901),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_700),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_703),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_703),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_830),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_880),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_836),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_706),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_706),
.Y(n_1444)
);

CKINVDCx20_ASAP7_75t_R g1445 ( 
.A(n_916),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_959),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_721),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_707),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_707),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_722),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_712),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_712),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_723),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1151),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_717),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_717),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_734),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_734),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_747),
.Y(n_1459)
);

INVxp67_ASAP7_75t_SL g1460 ( 
.A(n_836),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_747),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_963),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_756),
.Y(n_1463)
);

CKINVDCx16_ASAP7_75t_R g1464 ( 
.A(n_986),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_698),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_756),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_767),
.B(n_3),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_758),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_758),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1025),
.B(n_4),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_761),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_761),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_724),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_744),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1057),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_725),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_765),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_765),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_698),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_771),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_771),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_698),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_790),
.Y(n_1483)
);

INVxp33_ASAP7_75t_L g1484 ( 
.A(n_790),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_733),
.B(n_715),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_793),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_793),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_727),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_704),
.Y(n_1489)
);

CKINVDCx14_ASAP7_75t_R g1490 ( 
.A(n_744),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_797),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_797),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_803),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_985),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_803),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_806),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_806),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_812),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_728),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_732),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_812),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_821),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_821),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_825),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_825),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_841),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_841),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_844),
.Y(n_1508)
);

BUFx5_ASAP7_75t_L g1509 ( 
.A(n_844),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1023),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_852),
.Y(n_1511)
);

INVxp33_ASAP7_75t_L g1512 ( 
.A(n_852),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_736),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_737),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_854),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_854),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_859),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_859),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_704),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_865),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_865),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_871),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_739),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_871),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_872),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1026),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_872),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_876),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1059),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_741),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_876),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_704),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_886),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_879),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_733),
.B(n_774),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_886),
.Y(n_1536)
);

INVxp33_ASAP7_75t_L g1537 ( 
.A(n_890),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_743),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_890),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_746),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_891),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_891),
.Y(n_1542)
);

NOR2xp67_ASAP7_75t_L g1543 ( 
.A(n_767),
.B(n_3),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_897),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_748),
.Y(n_1545)
);

INVxp33_ASAP7_75t_L g1546 ( 
.A(n_897),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_898),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_898),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_749),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_904),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_904),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_750),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_718),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_879),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_906),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_906),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_915),
.Y(n_1557)
);

NOR2xp67_ASAP7_75t_L g1558 ( 
.A(n_796),
.B(n_4),
.Y(n_1558)
);

CKINVDCx20_ASAP7_75t_R g1559 ( 
.A(n_1065),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_718),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_915),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_917),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_917),
.Y(n_1563)
);

INVxp33_ASAP7_75t_SL g1564 ( 
.A(n_753),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_921),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_921),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_930),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_757),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_930),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_759),
.Y(n_1570)
);

INVx1_ASAP7_75t_SL g1571 ( 
.A(n_1071),
.Y(n_1571)
);

INVxp67_ASAP7_75t_SL g1572 ( 
.A(n_718),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_745),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_945),
.Y(n_1574)
);

CKINVDCx20_ASAP7_75t_R g1575 ( 
.A(n_1076),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_745),
.Y(n_1576)
);

CKINVDCx20_ASAP7_75t_R g1577 ( 
.A(n_1083),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_945),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_960),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_960),
.Y(n_1580)
);

INVxp67_ASAP7_75t_SL g1581 ( 
.A(n_745),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_961),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1089),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_760),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_754),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_961),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_962),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1093),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_962),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_754),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_964),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_964),
.Y(n_1592)
);

INVxp33_ASAP7_75t_SL g1593 ( 
.A(n_764),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_768),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_976),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_976),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_977),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_977),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_770),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_772),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_777),
.Y(n_1601)
);

CKINVDCx14_ASAP7_75t_R g1602 ( 
.A(n_879),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_990),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_990),
.Y(n_1604)
);

INVxp33_ASAP7_75t_L g1605 ( 
.A(n_994),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_994),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_778),
.Y(n_1607)
);

NOR2xp67_ASAP7_75t_L g1608 ( 
.A(n_796),
.B(n_5),
.Y(n_1608)
);

CKINVDCx16_ASAP7_75t_R g1609 ( 
.A(n_879),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_997),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_754),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_997),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1008),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1094),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1008),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_780),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_781),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1010),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1010),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1011),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1011),
.Y(n_1621)
);

CKINVDCx16_ASAP7_75t_R g1622 ( 
.A(n_946),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1012),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_783),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_784),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1012),
.Y(n_1626)
);

CKINVDCx16_ASAP7_75t_R g1627 ( 
.A(n_946),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1015),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_785),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1015),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_946),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1136),
.Y(n_1632)
);

INVxp67_ASAP7_75t_L g1633 ( 
.A(n_1018),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_787),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1018),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1021),
.Y(n_1636)
);

CKINVDCx16_ASAP7_75t_R g1637 ( 
.A(n_946),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_762),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_788),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1021),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1032),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_789),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_792),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1032),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1036),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1036),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1039),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_794),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1039),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1040),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1040),
.Y(n_1651)
);

INVxp33_ASAP7_75t_L g1652 ( 
.A(n_1043),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_795),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_762),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1043),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1000),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_799),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1048),
.Y(n_1658)
);

CKINVDCx14_ASAP7_75t_R g1659 ( 
.A(n_1000),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1048),
.Y(n_1660)
);

INVxp67_ASAP7_75t_SL g1661 ( 
.A(n_762),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1323),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1317),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1320),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_1226),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1325),
.Y(n_1666)
);

CKINVDCx20_ASAP7_75t_R g1667 ( 
.A(n_1226),
.Y(n_1667)
);

CKINVDCx20_ASAP7_75t_R g1668 ( 
.A(n_1230),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1431),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1376),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1414),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1572),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1329),
.Y(n_1673)
);

CKINVDCx16_ASAP7_75t_R g1674 ( 
.A(n_1380),
.Y(n_1674)
);

CKINVDCx5p33_ASAP7_75t_R g1675 ( 
.A(n_1330),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1333),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1230),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1581),
.Y(n_1678)
);

INVxp67_ASAP7_75t_SL g1679 ( 
.A(n_1227),
.Y(n_1679)
);

CKINVDCx20_ASAP7_75t_R g1680 ( 
.A(n_1234),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1590),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1661),
.Y(n_1682)
);

CKINVDCx16_ASAP7_75t_R g1683 ( 
.A(n_1464),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1250),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1335),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1227),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1252),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1349),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1281),
.Y(n_1689)
);

CKINVDCx20_ASAP7_75t_R g1690 ( 
.A(n_1234),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_1386),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1356),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1259),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1387),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1360),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1391),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1361),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1363),
.Y(n_1698)
);

INVxp33_ASAP7_75t_L g1699 ( 
.A(n_1600),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1302),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1259),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1364),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1392),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1607),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1371),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1374),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1377),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1382),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1398),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1396),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1383),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_1400),
.Y(n_1712)
);

CKINVDCx5p33_ASAP7_75t_R g1713 ( 
.A(n_1416),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1419),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1384),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1423),
.Y(n_1716)
);

INVxp67_ASAP7_75t_SL g1717 ( 
.A(n_1237),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1385),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1265),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1302),
.Y(n_1720)
);

CKINVDCx16_ASAP7_75t_R g1721 ( 
.A(n_1255),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1388),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1265),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1571),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1268),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_1427),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1642),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1283),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1389),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1395),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1447),
.Y(n_1731)
);

CKINVDCx20_ASAP7_75t_R g1732 ( 
.A(n_1268),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1450),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1399),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1401),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_1282),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1402),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1408),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1412),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1413),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1415),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1417),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1453),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1347),
.Y(n_1744)
);

CKINVDCx20_ASAP7_75t_R g1745 ( 
.A(n_1282),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1418),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_1334),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1237),
.Y(n_1748)
);

CKINVDCx16_ASAP7_75t_R g1749 ( 
.A(n_1262),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1420),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_1334),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1357),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1421),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1485),
.B(n_798),
.Y(n_1754)
);

CKINVDCx20_ASAP7_75t_R g1755 ( 
.A(n_1353),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_1473),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_1473),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1476),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1476),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1347),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1488),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_SL g1762 ( 
.A(n_1299),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1358),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1241),
.Y(n_1764)
);

NOR2xp67_ASAP7_75t_L g1765 ( 
.A(n_1535),
.B(n_615),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1425),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1648),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1428),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1429),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1430),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1353),
.Y(n_1771)
);

INVxp67_ASAP7_75t_L g1772 ( 
.A(n_1390),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1488),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1432),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1434),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1365),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1435),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1284),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1286),
.Y(n_1779)
);

INVxp33_ASAP7_75t_SL g1780 ( 
.A(n_1221),
.Y(n_1780)
);

NOR2xp67_ASAP7_75t_L g1781 ( 
.A(n_1499),
.B(n_1500),
.Y(n_1781)
);

CKINVDCx20_ASAP7_75t_R g1782 ( 
.A(n_1365),
.Y(n_1782)
);

CKINVDCx20_ASAP7_75t_R g1783 ( 
.A(n_1403),
.Y(n_1783)
);

BUFx3_ASAP7_75t_L g1784 ( 
.A(n_1241),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1403),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_1409),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1288),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1289),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1396),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1409),
.Y(n_1790)
);

INVxp67_ASAP7_75t_SL g1791 ( 
.A(n_1410),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1290),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1411),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1292),
.Y(n_1794)
);

CKINVDCx20_ASAP7_75t_R g1795 ( 
.A(n_1411),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1293),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1499),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1294),
.Y(n_1798)
);

NOR2xp67_ASAP7_75t_L g1799 ( 
.A(n_1500),
.B(n_621),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1513),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1513),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1441),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1410),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1441),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1295),
.Y(n_1805)
);

CKINVDCx5p33_ASAP7_75t_R g1806 ( 
.A(n_1514),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1445),
.Y(n_1807)
);

CKINVDCx14_ASAP7_75t_R g1808 ( 
.A(n_1490),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1297),
.Y(n_1809)
);

CKINVDCx20_ASAP7_75t_R g1810 ( 
.A(n_1445),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1514),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1446),
.Y(n_1812)
);

CKINVDCx5p33_ASAP7_75t_R g1813 ( 
.A(n_1523),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1523),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1298),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1530),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1274),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1300),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1530),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1304),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1538),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1306),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1307),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1538),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1309),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1311),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1446),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_1462),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1460),
.B(n_798),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_1462),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1312),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1433),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1540),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1540),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1313),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1315),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1316),
.Y(n_1837)
);

NOR2xp67_ASAP7_75t_L g1838 ( 
.A(n_1545),
.B(n_622),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1318),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1494),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1324),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1358),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1326),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1328),
.Y(n_1844)
);

CKINVDCx20_ASAP7_75t_R g1845 ( 
.A(n_1494),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1331),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1545),
.Y(n_1847)
);

CKINVDCx20_ASAP7_75t_R g1848 ( 
.A(n_1510),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1332),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1339),
.Y(n_1850)
);

CKINVDCx20_ASAP7_75t_R g1851 ( 
.A(n_1510),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1340),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1283),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_L g1854 ( 
.A(n_1549),
.B(n_623),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_1549),
.Y(n_1855)
);

CKINVDCx5p33_ASAP7_75t_R g1856 ( 
.A(n_1552),
.Y(n_1856)
);

CKINVDCx20_ASAP7_75t_R g1857 ( 
.A(n_1526),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1305),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1552),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1341),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1568),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1568),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1362),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1570),
.Y(n_1864)
);

CKINVDCx20_ASAP7_75t_R g1865 ( 
.A(n_1526),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1342),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1344),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1570),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1594),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1345),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1529),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1406),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1362),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1594),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1378),
.Y(n_1875)
);

CKINVDCx20_ASAP7_75t_R g1876 ( 
.A(n_1529),
.Y(n_1876)
);

CKINVDCx5p33_ASAP7_75t_R g1877 ( 
.A(n_1599),
.Y(n_1877)
);

CKINVDCx20_ASAP7_75t_R g1878 ( 
.A(n_1559),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1599),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1632),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1601),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1601),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1616),
.Y(n_1883)
);

CKINVDCx20_ASAP7_75t_R g1884 ( 
.A(n_1559),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_1575),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1346),
.Y(n_1886)
);

INVxp33_ASAP7_75t_SL g1887 ( 
.A(n_1221),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1372),
.B(n_858),
.Y(n_1888)
);

CKINVDCx20_ASAP7_75t_R g1889 ( 
.A(n_1575),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1378),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1351),
.Y(n_1891)
);

INVxp67_ASAP7_75t_SL g1892 ( 
.A(n_1433),
.Y(n_1892)
);

CKINVDCx20_ASAP7_75t_R g1893 ( 
.A(n_1577),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1616),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1354),
.Y(n_1895)
);

CKINVDCx20_ASAP7_75t_R g1896 ( 
.A(n_1577),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1617),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1257),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1617),
.Y(n_1899)
);

CKINVDCx20_ASAP7_75t_R g1900 ( 
.A(n_1583),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1258),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1260),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1261),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_1624),
.Y(n_1904)
);

INVxp67_ASAP7_75t_SL g1905 ( 
.A(n_1475),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1624),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1264),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1625),
.Y(n_1908)
);

CKINVDCx16_ASAP7_75t_R g1909 ( 
.A(n_1285),
.Y(n_1909)
);

CKINVDCx20_ASAP7_75t_R g1910 ( 
.A(n_1583),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1266),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1625),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1274),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1267),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1269),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1270),
.Y(n_1916)
);

INVxp67_ASAP7_75t_L g1917 ( 
.A(n_1424),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1629),
.Y(n_1918)
);

CKINVDCx5p33_ASAP7_75t_R g1919 ( 
.A(n_1629),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1426),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1305),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_L g1922 ( 
.A(n_1370),
.B(n_858),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1271),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1634),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1272),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1370),
.B(n_929),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1588),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_1588),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1273),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1275),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1634),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1276),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1639),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1277),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1584),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1278),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1279),
.Y(n_1937)
);

CKINVDCx20_ASAP7_75t_R g1938 ( 
.A(n_1614),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1280),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1321),
.Y(n_1940)
);

INVxp67_ASAP7_75t_SL g1941 ( 
.A(n_1440),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1639),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1375),
.B(n_929),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1643),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1321),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1321),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1321),
.Y(n_1947)
);

BUFx6f_ASAP7_75t_SL g1948 ( 
.A(n_1299),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1643),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1375),
.B(n_947),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1337),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1653),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1653),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1337),
.Y(n_1954)
);

NOR2xp67_ASAP7_75t_L g1955 ( 
.A(n_1657),
.B(n_628),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1337),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1657),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1337),
.Y(n_1958)
);

INVxp67_ASAP7_75t_SL g1959 ( 
.A(n_1440),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_1614),
.Y(n_1960)
);

BUFx2_ASAP7_75t_L g1961 ( 
.A(n_1236),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1236),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1440),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1240),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1243),
.Y(n_1965)
);

INVxp67_ASAP7_75t_SL g1966 ( 
.A(n_1440),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1240),
.Y(n_1967)
);

CKINVDCx20_ASAP7_75t_R g1968 ( 
.A(n_1381),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_1407),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1407),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1240),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1404),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1404),
.Y(n_1973)
);

INVxp67_ASAP7_75t_SL g1974 ( 
.A(n_1442),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1404),
.Y(n_1975)
);

CKINVDCx20_ASAP7_75t_R g1976 ( 
.A(n_1381),
.Y(n_1976)
);

XOR2xp5_ASAP7_75t_L g1977 ( 
.A(n_1287),
.B(n_1149),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1243),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1247),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1310),
.B(n_1000),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1222),
.Y(n_1981)
);

CKINVDCx20_ASAP7_75t_R g1982 ( 
.A(n_1303),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1247),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1291),
.Y(n_1984)
);

INVxp67_ASAP7_75t_L g1985 ( 
.A(n_1534),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1223),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1291),
.Y(n_1987)
);

CKINVDCx14_ASAP7_75t_R g1988 ( 
.A(n_1490),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1564),
.B(n_947),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1225),
.Y(n_1990)
);

CKINVDCx20_ASAP7_75t_R g1991 ( 
.A(n_1308),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_1564),
.Y(n_1992)
);

INVx1_ASAP7_75t_SL g1993 ( 
.A(n_1359),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1228),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1229),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1593),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1593),
.B(n_1068),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1231),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1232),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1327),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1233),
.Y(n_2001)
);

INVxp67_ASAP7_75t_SL g2002 ( 
.A(n_1442),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1343),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1367),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1310),
.Y(n_2005)
);

NOR2xp67_ASAP7_75t_L g2006 ( 
.A(n_1319),
.B(n_630),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1436),
.B(n_1068),
.Y(n_2007)
);

INVxp67_ASAP7_75t_SL g2008 ( 
.A(n_1442),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1314),
.Y(n_2009)
);

CKINVDCx20_ASAP7_75t_R g2010 ( 
.A(n_1602),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1235),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_1609),
.Y(n_2012)
);

CKINVDCx20_ASAP7_75t_R g2013 ( 
.A(n_1602),
.Y(n_2013)
);

INVxp67_ASAP7_75t_SL g2014 ( 
.A(n_1442),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1238),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1239),
.Y(n_2016)
);

CKINVDCx20_ASAP7_75t_R g2017 ( 
.A(n_1659),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1245),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1246),
.Y(n_2019)
);

INVxp67_ASAP7_75t_SL g2020 ( 
.A(n_1534),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_1659),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1622),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1554),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1627),
.Y(n_2024)
);

CKINVDCx20_ASAP7_75t_R g2025 ( 
.A(n_1637),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1686),
.B(n_1263),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1728),
.Y(n_2027)
);

INVx4_ASAP7_75t_L g2028 ( 
.A(n_1710),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1778),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_2010),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1779),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1724),
.Y(n_2032)
);

CKINVDCx20_ASAP7_75t_R g2033 ( 
.A(n_1665),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_1728),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1880),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1993),
.B(n_1338),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1787),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1905),
.B(n_1244),
.Y(n_2038)
);

OA21x2_ASAP7_75t_L g2039 ( 
.A1(n_1981),
.A2(n_1251),
.B(n_1249),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1765),
.B(n_1366),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1662),
.B(n_1338),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1853),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1686),
.B(n_1479),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1788),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1792),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1784),
.B(n_1479),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1808),
.B(n_1352),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_1665),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1794),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1988),
.B(n_1352),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1796),
.Y(n_2051)
);

INVx3_ASAP7_75t_L g2052 ( 
.A(n_1710),
.Y(n_2052)
);

OA21x2_ASAP7_75t_L g2053 ( 
.A1(n_1986),
.A2(n_1256),
.B(n_1254),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1710),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1710),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1789),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1798),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1805),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1809),
.Y(n_2059)
);

OAI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1754),
.A2(n_1348),
.B1(n_1244),
.B2(n_1253),
.Y(n_2060)
);

INVx2_ASAP7_75t_L g2061 ( 
.A(n_1853),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1670),
.B(n_1314),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1784),
.B(n_1482),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1815),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1679),
.B(n_1482),
.Y(n_2065)
);

BUFx8_ASAP7_75t_L g2066 ( 
.A(n_1762),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1818),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1789),
.Y(n_2068)
);

CKINVDCx20_ASAP7_75t_R g2069 ( 
.A(n_1667),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_1982),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1789),
.Y(n_2071)
);

CKINVDCx5p33_ASAP7_75t_R g2072 ( 
.A(n_2010),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1858),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1717),
.B(n_1489),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1699),
.B(n_1350),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1820),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_2013),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1858),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1822),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1823),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1825),
.Y(n_2081)
);

HB1xp67_ASAP7_75t_L g2082 ( 
.A(n_2004),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_2013),
.Y(n_2083)
);

NAND2xp33_ASAP7_75t_SL g2084 ( 
.A(n_1888),
.B(n_1467),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1826),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1817),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1671),
.B(n_1336),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1748),
.B(n_1359),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_2017),
.Y(n_2089)
);

BUFx6f_ASAP7_75t_L g2090 ( 
.A(n_1940),
.Y(n_2090)
);

BUFx3_ASAP7_75t_L g2091 ( 
.A(n_1817),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1831),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1945),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_1921),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_2017),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1982),
.Y(n_2096)
);

AND2x6_ASAP7_75t_L g2097 ( 
.A(n_1980),
.B(n_1301),
.Y(n_2097)
);

OR2x6_ASAP7_75t_L g2098 ( 
.A(n_1700),
.B(n_1474),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1921),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1835),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1941),
.B(n_1336),
.Y(n_2101)
);

NOR2xp67_ASAP7_75t_L g2102 ( 
.A(n_1663),
.B(n_1224),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2009),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2009),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1836),
.Y(n_2105)
);

INVxp67_ASAP7_75t_L g2106 ( 
.A(n_2023),
.Y(n_2106)
);

CKINVDCx16_ASAP7_75t_R g2107 ( 
.A(n_1721),
.Y(n_2107)
);

BUFx2_ASAP7_75t_L g2108 ( 
.A(n_1991),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_2007),
.A2(n_1242),
.B(n_1394),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_1922),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1837),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_1990),
.A2(n_1242),
.B(n_1394),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_2021),
.Y(n_2113)
);

CKINVDCx20_ASAP7_75t_R g2114 ( 
.A(n_1667),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1764),
.B(n_1489),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1692),
.Y(n_2116)
);

INVx3_ASAP7_75t_L g2117 ( 
.A(n_1946),
.Y(n_2117)
);

NOR2xp33_ASAP7_75t_L g2118 ( 
.A(n_1684),
.B(n_1253),
.Y(n_2118)
);

AND2x6_ASAP7_75t_L g2119 ( 
.A(n_1687),
.B(n_779),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1839),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1841),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_1947),
.Y(n_2122)
);

INVx3_ASAP7_75t_L g2123 ( 
.A(n_1951),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1843),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1844),
.Y(n_2125)
);

INVxp67_ASAP7_75t_L g2126 ( 
.A(n_1926),
.Y(n_2126)
);

OAI21x1_ASAP7_75t_L g2127 ( 
.A1(n_1994),
.A2(n_1405),
.B(n_1397),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1846),
.Y(n_2128)
);

NAND2x1_ASAP7_75t_L g2129 ( 
.A(n_1995),
.B(n_1396),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1695),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_1791),
.B(n_1519),
.Y(n_2131)
);

AND2x2_ASAP7_75t_SL g2132 ( 
.A(n_1943),
.B(n_1470),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1849),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1799),
.B(n_1366),
.Y(n_2134)
);

CKINVDCx20_ASAP7_75t_R g2135 ( 
.A(n_1668),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1850),
.Y(n_2136)
);

CKINVDCx5p33_ASAP7_75t_R g2137 ( 
.A(n_2021),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1852),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1959),
.B(n_1397),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_1772),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1860),
.Y(n_2141)
);

BUFx6f_ASAP7_75t_L g2142 ( 
.A(n_1954),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1963),
.B(n_1405),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1866),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_1991),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_SL g2146 ( 
.A1(n_1977),
.A2(n_1177),
.B1(n_1182),
.B2(n_1176),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1867),
.Y(n_2147)
);

AND3x2_ASAP7_75t_L g2148 ( 
.A(n_1961),
.B(n_1322),
.C(n_1296),
.Y(n_2148)
);

OA21x2_ASAP7_75t_L g2149 ( 
.A1(n_1998),
.A2(n_1355),
.B(n_1422),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1870),
.Y(n_2150)
);

INVx3_ASAP7_75t_L g2151 ( 
.A(n_1956),
.Y(n_2151)
);

INVx5_ASAP7_75t_L g2152 ( 
.A(n_1913),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1886),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1891),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_1803),
.B(n_1519),
.Y(n_2155)
);

INVxp67_ASAP7_75t_L g2156 ( 
.A(n_1950),
.Y(n_2156)
);

AOI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_1781),
.A2(n_1997),
.B1(n_1989),
.B2(n_1704),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1895),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1898),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1697),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1966),
.B(n_1422),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1985),
.B(n_1554),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1698),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1901),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1902),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_1903),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1958),
.Y(n_2167)
);

CKINVDCx5p33_ASAP7_75t_R g2168 ( 
.A(n_1752),
.Y(n_2168)
);

INVx3_ASAP7_75t_L g2169 ( 
.A(n_1964),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1907),
.Y(n_2170)
);

NOR2xp33_ASAP7_75t_R g2171 ( 
.A(n_1969),
.B(n_1656),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1911),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1702),
.Y(n_2173)
);

BUFx2_ASAP7_75t_L g2174 ( 
.A(n_2000),
.Y(n_2174)
);

CKINVDCx20_ASAP7_75t_R g2175 ( 
.A(n_1668),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_1672),
.B(n_1678),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_1872),
.B(n_1631),
.Y(n_2177)
);

CKINVDCx5p33_ASAP7_75t_R g2178 ( 
.A(n_2005),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_2003),
.Y(n_2179)
);

CKINVDCx5p33_ASAP7_75t_R g2180 ( 
.A(n_1970),
.Y(n_2180)
);

NOR2xp33_ASAP7_75t_L g2181 ( 
.A(n_1681),
.B(n_1368),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_1917),
.B(n_1631),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1920),
.B(n_1935),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_1832),
.B(n_1532),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1669),
.B(n_1369),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1914),
.Y(n_2186)
);

NAND2xp33_ASAP7_75t_L g2187 ( 
.A(n_1999),
.B(n_1366),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1915),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_1916),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1923),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1925),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1929),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1930),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_1974),
.B(n_1396),
.Y(n_2194)
);

OA21x2_ASAP7_75t_L g2195 ( 
.A1(n_2001),
.A2(n_1553),
.B(n_1532),
.Y(n_2195)
);

CKINVDCx5p33_ASAP7_75t_R g2196 ( 
.A(n_1664),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1932),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2002),
.B(n_1366),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1705),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_1706),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1934),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1727),
.B(n_1369),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_1666),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1936),
.Y(n_2204)
);

INVx6_ASAP7_75t_L g2205 ( 
.A(n_1913),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1707),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1892),
.B(n_1553),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_1967),
.Y(n_2208)
);

INVx3_ASAP7_75t_L g2209 ( 
.A(n_1971),
.Y(n_2209)
);

BUFx3_ASAP7_75t_L g2210 ( 
.A(n_2011),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1937),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2008),
.B(n_1366),
.Y(n_2212)
);

HB1xp67_ASAP7_75t_L g2213 ( 
.A(n_1767),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_1939),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2014),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1708),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1711),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2015),
.Y(n_2218)
);

AOI22x1_ASAP7_75t_SL g2219 ( 
.A1(n_1968),
.A2(n_1204),
.B1(n_769),
.B2(n_1122),
.Y(n_2219)
);

NOR2xp33_ASAP7_75t_L g2220 ( 
.A(n_1682),
.B(n_1368),
.Y(n_2220)
);

CKINVDCx5p33_ASAP7_75t_R g2221 ( 
.A(n_1673),
.Y(n_2221)
);

CKINVDCx5p33_ASAP7_75t_R g2222 ( 
.A(n_1675),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1972),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2016),
.B(n_1366),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2018),
.Y(n_2225)
);

OR2x6_ASAP7_75t_L g2226 ( 
.A(n_1720),
.B(n_1248),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2019),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_1715),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1829),
.B(n_1454),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1689),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1718),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1722),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1729),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1730),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1734),
.Y(n_2235)
);

CKINVDCx5p33_ASAP7_75t_R g2236 ( 
.A(n_1676),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1735),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2020),
.B(n_1979),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_1973),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1737),
.B(n_1366),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1738),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1739),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1685),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1740),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1741),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1742),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1746),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1750),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1753),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1766),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1768),
.Y(n_2251)
);

INVx3_ASAP7_75t_L g2252 ( 
.A(n_1975),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1769),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1770),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1774),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1775),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1777),
.Y(n_2257)
);

INVxp33_ASAP7_75t_SL g2258 ( 
.A(n_1983),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_1762),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1838),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_1762),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1854),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1955),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1948),
.Y(n_2264)
);

OR2x6_ASAP7_75t_L g2265 ( 
.A(n_1875),
.B(n_1084),
.Y(n_2265)
);

INVx2_ASAP7_75t_L g2266 ( 
.A(n_1948),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_1948),
.Y(n_2267)
);

CKINVDCx5p33_ASAP7_75t_R g2268 ( 
.A(n_1688),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1894),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1906),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1952),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1691),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_1694),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_1984),
.B(n_1731),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2006),
.B(n_1373),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1696),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1744),
.Y(n_2277)
);

NOR2x1_ASAP7_75t_L g2278 ( 
.A(n_2025),
.B(n_1543),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1760),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1703),
.Y(n_2280)
);

INVx3_ASAP7_75t_L g2281 ( 
.A(n_1733),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_SL g2282 ( 
.A1(n_2025),
.A2(n_769),
.B1(n_1122),
.B2(n_1157),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1709),
.B(n_1373),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_1763),
.Y(n_2284)
);

CKINVDCx5p33_ASAP7_75t_R g2285 ( 
.A(n_1712),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1713),
.B(n_1373),
.Y(n_2286)
);

CKINVDCx5p33_ASAP7_75t_R g2287 ( 
.A(n_1714),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_1842),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1716),
.B(n_1373),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1863),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_SL g2291 ( 
.A1(n_1749),
.A2(n_1157),
.B1(n_786),
.B2(n_878),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1873),
.Y(n_2292)
);

CKINVDCx20_ASAP7_75t_R g2293 ( 
.A(n_1677),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_1726),
.B(n_1373),
.Y(n_2294)
);

OA21x2_ASAP7_75t_L g2295 ( 
.A1(n_1743),
.A2(n_1573),
.B(n_1560),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1890),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1962),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_R g2298 ( 
.A(n_1992),
.B(n_800),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1965),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1756),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1978),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_1987),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_1909),
.Y(n_2303)
);

CKINVDCx5p33_ASAP7_75t_R g2304 ( 
.A(n_2012),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1757),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1758),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_1759),
.B(n_1484),
.Y(n_2307)
);

NOR2xp33_ASAP7_75t_L g2308 ( 
.A(n_1887),
.B(n_1484),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1761),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_1674),
.Y(n_2310)
);

BUFx6f_ASAP7_75t_L g2311 ( 
.A(n_1773),
.Y(n_2311)
);

CKINVDCx20_ASAP7_75t_R g2312 ( 
.A(n_1677),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1797),
.B(n_1373),
.Y(n_2313)
);

AND2x4_ASAP7_75t_L g2314 ( 
.A(n_1800),
.B(n_1560),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1801),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1806),
.B(n_1373),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_1683),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_1811),
.B(n_1512),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1813),
.Y(n_2319)
);

BUFx6f_ASAP7_75t_L g2320 ( 
.A(n_1814),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1816),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1819),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_1821),
.B(n_1512),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_1824),
.B(n_1509),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_1833),
.Y(n_2325)
);

AND2x4_ASAP7_75t_L g2326 ( 
.A(n_1834),
.B(n_1573),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1847),
.B(n_1509),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_SL g2328 ( 
.A(n_1855),
.B(n_1509),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_1856),
.Y(n_2329)
);

BUFx6f_ASAP7_75t_L g2330 ( 
.A(n_1859),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1861),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_1862),
.Y(n_2332)
);

INVx3_ASAP7_75t_L g2333 ( 
.A(n_1864),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_1868),
.B(n_1509),
.Y(n_2334)
);

CKINVDCx5p33_ASAP7_75t_R g2335 ( 
.A(n_2022),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_1869),
.Y(n_2336)
);

AOI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_1780),
.A2(n_1379),
.B1(n_1608),
.B2(n_1558),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1874),
.B(n_1537),
.Y(n_2338)
);

OR2x2_ASAP7_75t_L g2339 ( 
.A(n_1877),
.B(n_1537),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_1879),
.Y(n_2340)
);

BUFx6f_ASAP7_75t_L g2341 ( 
.A(n_1881),
.Y(n_2341)
);

NAND2xp33_ASAP7_75t_L g2342 ( 
.A(n_1996),
.B(n_1509),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_1882),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1883),
.Y(n_2344)
);

OA21x2_ASAP7_75t_L g2345 ( 
.A1(n_1897),
.A2(n_1611),
.B(n_1576),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_1899),
.Y(n_2346)
);

CKINVDCx5p33_ASAP7_75t_R g2347 ( 
.A(n_2024),
.Y(n_2347)
);

INVx3_ASAP7_75t_L g2348 ( 
.A(n_1904),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_1908),
.B(n_1576),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1912),
.Y(n_2350)
);

NOR2xp33_ASAP7_75t_L g2351 ( 
.A(n_1780),
.B(n_1546),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_1918),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_1919),
.Y(n_2353)
);

AND2x6_ASAP7_75t_L g2354 ( 
.A(n_1924),
.B(n_779),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1931),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_1933),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_1942),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_1944),
.B(n_1546),
.Y(n_2358)
);

INVx3_ASAP7_75t_L g2359 ( 
.A(n_1949),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_1953),
.Y(n_2360)
);

NOR2xp33_ASAP7_75t_R g2361 ( 
.A(n_1957),
.B(n_802),
.Y(n_2361)
);

NOR2x1_ASAP7_75t_L g2362 ( 
.A(n_1968),
.B(n_1437),
.Y(n_2362)
);

OAI21x1_ASAP7_75t_L g2363 ( 
.A1(n_1680),
.A2(n_1654),
.B(n_1638),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1680),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_L g2365 ( 
.A(n_1976),
.B(n_1605),
.Y(n_2365)
);

INVx3_ASAP7_75t_L g2366 ( 
.A(n_1690),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1690),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_1693),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_1976),
.B(n_1509),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_1693),
.B(n_1605),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_1960),
.B(n_1509),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_1701),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_1960),
.B(n_1465),
.Y(n_2373)
);

AND3x2_ASAP7_75t_L g2374 ( 
.A(n_1701),
.B(n_845),
.C(n_779),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1938),
.B(n_1465),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_1938),
.A2(n_833),
.B1(n_941),
.B2(n_735),
.Y(n_2376)
);

OA21x2_ASAP7_75t_L g2377 ( 
.A1(n_1719),
.A2(n_1638),
.B(n_1611),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_1719),
.B(n_1652),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_1723),
.Y(n_2379)
);

OAI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_1723),
.A2(n_810),
.B1(n_813),
.B2(n_807),
.Y(n_2380)
);

INVx3_ASAP7_75t_L g2381 ( 
.A(n_1725),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1725),
.Y(n_2382)
);

OA21x2_ASAP7_75t_L g2383 ( 
.A1(n_1732),
.A2(n_1654),
.B(n_1641),
.Y(n_2383)
);

BUFx6f_ASAP7_75t_L g2384 ( 
.A(n_1732),
.Y(n_2384)
);

AND2x4_ASAP7_75t_L g2385 ( 
.A(n_1736),
.B(n_1438),
.Y(n_2385)
);

NAND2xp33_ASAP7_75t_R g2386 ( 
.A(n_1736),
.B(n_814),
.Y(n_2386)
);

CKINVDCx5p33_ASAP7_75t_R g2387 ( 
.A(n_1745),
.Y(n_2387)
);

CKINVDCx16_ASAP7_75t_R g2388 ( 
.A(n_1745),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1747),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1747),
.Y(n_2390)
);

CKINVDCx20_ASAP7_75t_R g2391 ( 
.A(n_1751),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1751),
.Y(n_2392)
);

OR2x2_ASAP7_75t_L g2393 ( 
.A(n_1755),
.B(n_1652),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_1755),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_1771),
.B(n_1393),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_1771),
.B(n_1471),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_1776),
.Y(n_2397)
);

OAI22xp5_ASAP7_75t_SL g2398 ( 
.A1(n_1776),
.A2(n_965),
.B1(n_970),
.B2(n_949),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_1782),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_1782),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1783),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1783),
.B(n_1465),
.Y(n_2402)
);

INVx3_ASAP7_75t_L g2403 ( 
.A(n_1785),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_1785),
.B(n_1511),
.Y(n_2404)
);

BUFx2_ASAP7_75t_L g2405 ( 
.A(n_1786),
.Y(n_2405)
);

AND2x6_ASAP7_75t_L g2406 ( 
.A(n_1786),
.B(n_845),
.Y(n_2406)
);

HB1xp67_ASAP7_75t_L g2407 ( 
.A(n_1790),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_1790),
.B(n_1439),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_1793),
.B(n_1465),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1793),
.Y(n_2410)
);

AND3x2_ASAP7_75t_L g2411 ( 
.A(n_1795),
.B(n_894),
.C(n_845),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_1795),
.B(n_1556),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_1802),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_1802),
.Y(n_2414)
);

CKINVDCx20_ASAP7_75t_R g2415 ( 
.A(n_1804),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1804),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_1807),
.B(n_1585),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_1807),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_1810),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_1810),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1812),
.B(n_1585),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_1812),
.Y(n_2422)
);

CKINVDCx5p33_ASAP7_75t_R g2423 ( 
.A(n_1827),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1827),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_1828),
.B(n_1443),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1828),
.Y(n_2426)
);

CKINVDCx5p33_ASAP7_75t_R g2427 ( 
.A(n_1830),
.Y(n_2427)
);

OA21x2_ASAP7_75t_L g2428 ( 
.A1(n_1830),
.A2(n_1636),
.B(n_1635),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_1840),
.B(n_1587),
.Y(n_2429)
);

INVxp67_ASAP7_75t_L g2430 ( 
.A(n_1840),
.Y(n_2430)
);

XNOR2xp5_ASAP7_75t_L g2431 ( 
.A(n_1845),
.B(n_978),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_1845),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_1848),
.B(n_1444),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_1848),
.Y(n_2434)
);

AND2x4_ASAP7_75t_L g2435 ( 
.A(n_1851),
.B(n_1448),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_1851),
.Y(n_2436)
);

HB1xp67_ASAP7_75t_L g2437 ( 
.A(n_2032),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2043),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2132),
.B(n_1585),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2043),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_2229),
.B(n_1612),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_2035),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2043),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2046),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2046),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2046),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2112),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2195),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_2075),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_2195),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2195),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2307),
.B(n_1621),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_2063),
.B(n_2131),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2149),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2063),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2149),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2063),
.Y(n_2457)
);

NAND2xp33_ASAP7_75t_SL g2458 ( 
.A(n_2060),
.B(n_1084),
.Y(n_2458)
);

OAI22xp5_ASAP7_75t_SL g2459 ( 
.A1(n_2146),
.A2(n_1865),
.B1(n_1871),
.B2(n_1857),
.Y(n_2459)
);

INVx3_ASAP7_75t_L g2460 ( 
.A(n_2149),
.Y(n_2460)
);

AND2x4_ASAP7_75t_L g2461 ( 
.A(n_2131),
.B(n_1449),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2159),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2164),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2318),
.B(n_1633),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_2172),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2112),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2165),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2166),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2170),
.Y(n_2469)
);

BUFx6f_ASAP7_75t_L g2470 ( 
.A(n_2172),
.Y(n_2470)
);

INVx1_ASAP7_75t_SL g2471 ( 
.A(n_2323),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2186),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2188),
.Y(n_2473)
);

NAND2x1_ASAP7_75t_L g2474 ( 
.A(n_2039),
.B(n_1004),
.Y(n_2474)
);

AND2x2_ASAP7_75t_L g2475 ( 
.A(n_2338),
.B(n_1451),
.Y(n_2475)
);

AND2x4_ASAP7_75t_L g2476 ( 
.A(n_2131),
.B(n_1452),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2190),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2191),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2192),
.Y(n_2479)
);

HB1xp67_ASAP7_75t_L g2480 ( 
.A(n_2370),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2127),
.Y(n_2481)
);

OAI22xp5_ASAP7_75t_SL g2482 ( 
.A1(n_2282),
.A2(n_1865),
.B1(n_1871),
.B2(n_1857),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2193),
.Y(n_2483)
);

BUFx6f_ASAP7_75t_L g2484 ( 
.A(n_2172),
.Y(n_2484)
);

INVx2_ASAP7_75t_L g2485 ( 
.A(n_2127),
.Y(n_2485)
);

INVx3_ASAP7_75t_L g2486 ( 
.A(n_2295),
.Y(n_2486)
);

BUFx2_ASAP7_75t_L g2487 ( 
.A(n_2378),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2155),
.B(n_1585),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2027),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2197),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2205),
.Y(n_2491)
);

BUFx3_ASAP7_75t_L g2492 ( 
.A(n_2205),
.Y(n_2492)
);

INVx1_ASAP7_75t_SL g2493 ( 
.A(n_2358),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2201),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2204),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2027),
.Y(n_2496)
);

OAI22xp5_ASAP7_75t_SL g2497 ( 
.A1(n_2291),
.A2(n_1878),
.B1(n_1884),
.B2(n_1876),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2172),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2029),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_SL g2500 ( 
.A(n_2168),
.B(n_1876),
.Y(n_2500)
);

HB1xp67_ASAP7_75t_L g2501 ( 
.A(n_2373),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2034),
.Y(n_2502)
);

BUFx6f_ASAP7_75t_L g2503 ( 
.A(n_2189),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2031),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_2189),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2189),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2037),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2036),
.B(n_1455),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_SL g2509 ( 
.A(n_2406),
.Y(n_2509)
);

BUFx2_ASAP7_75t_L g2510 ( 
.A(n_2385),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2034),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2042),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2044),
.Y(n_2513)
);

INVxp67_ASAP7_75t_L g2514 ( 
.A(n_2308),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2351),
.B(n_1456),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2295),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2042),
.Y(n_2517)
);

AND2x4_ASAP7_75t_L g2518 ( 
.A(n_2155),
.B(n_1457),
.Y(n_2518)
);

BUFx2_ASAP7_75t_L g2519 ( 
.A(n_2385),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2061),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2045),
.Y(n_2521)
);

AND2x6_ASAP7_75t_L g2522 ( 
.A(n_2259),
.B(n_894),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2295),
.Y(n_2523)
);

BUFx6f_ASAP7_75t_SL g2524 ( 
.A(n_2406),
.Y(n_2524)
);

CKINVDCx20_ASAP7_75t_R g2525 ( 
.A(n_2033),
.Y(n_2525)
);

OAI22xp5_ASAP7_75t_SL g2526 ( 
.A1(n_2398),
.A2(n_1884),
.B1(n_1885),
.B2(n_1878),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2061),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2073),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_2132),
.B(n_1274),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2157),
.B(n_1066),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2049),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2073),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2051),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_2189),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2057),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2099),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2058),
.Y(n_2537)
);

NAND2xp5_ASAP7_75t_SL g2538 ( 
.A(n_2313),
.B(n_2316),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2059),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_2211),
.Y(n_2540)
);

INVxp67_ASAP7_75t_L g2541 ( 
.A(n_2308),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_SL g2542 ( 
.A(n_2406),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2324),
.B(n_1153),
.Y(n_2543)
);

BUFx6f_ASAP7_75t_L g2544 ( 
.A(n_2345),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2099),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2103),
.Y(n_2546)
);

CKINVDCx16_ASAP7_75t_R g2547 ( 
.A(n_2107),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2103),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2064),
.Y(n_2549)
);

BUFx2_ASAP7_75t_L g2550 ( 
.A(n_2385),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2067),
.Y(n_2551)
);

BUFx8_ASAP7_75t_L g2552 ( 
.A(n_2174),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2039),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_L g2554 ( 
.A(n_2110),
.B(n_815),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2076),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2079),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2080),
.Y(n_2557)
);

INVx3_ASAP7_75t_L g2558 ( 
.A(n_2039),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2081),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2085),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2408),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2104),
.Y(n_2562)
);

AND2x2_ASAP7_75t_L g2563 ( 
.A(n_2351),
.B(n_1458),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2155),
.B(n_1137),
.Y(n_2564)
);

AOI22xp5_ASAP7_75t_L g2565 ( 
.A1(n_2097),
.A2(n_1461),
.B1(n_1463),
.B2(n_1459),
.Y(n_2565)
);

INVx3_ASAP7_75t_L g2566 ( 
.A(n_2053),
.Y(n_2566)
);

INVx2_ASAP7_75t_L g2567 ( 
.A(n_2104),
.Y(n_2567)
);

HB1xp67_ASAP7_75t_L g2568 ( 
.A(n_2375),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2092),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2053),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2100),
.Y(n_2571)
);

INVxp67_ASAP7_75t_L g2572 ( 
.A(n_2339),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2053),
.Y(n_2573)
);

XNOR2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2431),
.B(n_1885),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2184),
.B(n_1137),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2184),
.B(n_1139),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2345),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2345),
.Y(n_2578)
);

AND2x4_ASAP7_75t_L g2579 ( 
.A(n_2184),
.B(n_1466),
.Y(n_2579)
);

INVx3_ASAP7_75t_L g2580 ( 
.A(n_2169),
.Y(n_2580)
);

INVx3_ASAP7_75t_L g2581 ( 
.A(n_2169),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2094),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2207),
.B(n_2327),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2094),
.Y(n_2584)
);

BUFx6f_ASAP7_75t_L g2585 ( 
.A(n_2211),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2334),
.B(n_894),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2105),
.Y(n_2587)
);

OAI22xp5_ASAP7_75t_SL g2588 ( 
.A1(n_2388),
.A2(n_1893),
.B1(n_1896),
.B2(n_1889),
.Y(n_2588)
);

OR2x2_ASAP7_75t_L g2589 ( 
.A(n_2393),
.B(n_1468),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2111),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2094),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2120),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2078),
.Y(n_2593)
);

BUFx3_ASAP7_75t_L g2594 ( 
.A(n_2205),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2121),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2371),
.B(n_931),
.Y(n_2596)
);

INVxp67_ASAP7_75t_L g2597 ( 
.A(n_2185),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2124),
.Y(n_2598)
);

OAI22xp5_ASAP7_75t_SL g2599 ( 
.A1(n_2033),
.A2(n_1893),
.B1(n_1896),
.B2(n_1889),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2211),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2125),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2402),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2128),
.Y(n_2603)
);

INVxp67_ASAP7_75t_L g2604 ( 
.A(n_2202),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2133),
.Y(n_2605)
);

BUFx2_ASAP7_75t_L g2606 ( 
.A(n_2408),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2136),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2314),
.B(n_1469),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2169),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_2138),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2141),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2144),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2208),
.Y(n_2613)
);

BUFx2_ASAP7_75t_L g2614 ( 
.A(n_2408),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2078),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2314),
.B(n_1472),
.Y(n_2616)
);

BUFx6f_ASAP7_75t_L g2617 ( 
.A(n_2363),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2116),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2147),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2150),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2153),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2116),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2425),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2154),
.Y(n_2624)
);

HB1xp67_ASAP7_75t_L g2625 ( 
.A(n_2409),
.Y(n_2625)
);

INVx3_ASAP7_75t_L g2626 ( 
.A(n_2208),
.Y(n_2626)
);

INVx3_ASAP7_75t_L g2627 ( 
.A(n_2209),
.Y(n_2627)
);

AND2x4_ASAP7_75t_L g2628 ( 
.A(n_2207),
.B(n_1477),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2158),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2417),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2130),
.Y(n_2631)
);

INVx2_ASAP7_75t_L g2632 ( 
.A(n_2130),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2230),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2207),
.B(n_1139),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2126),
.A2(n_817),
.B1(n_818),
.B2(n_816),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2065),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2065),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2065),
.Y(n_2638)
);

AND2x2_ASAP7_75t_L g2639 ( 
.A(n_2314),
.B(n_1478),
.Y(n_2639)
);

AND2x4_ASAP7_75t_L g2640 ( 
.A(n_2074),
.B(n_1480),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2074),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2326),
.B(n_1481),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2074),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_SL g2644 ( 
.A1(n_2048),
.A2(n_1910),
.B1(n_1927),
.B2(n_1900),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2115),
.B(n_1142),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_SL g2646 ( 
.A(n_2283),
.B(n_2286),
.Y(n_2646)
);

BUFx6f_ASAP7_75t_L g2647 ( 
.A(n_2211),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_SL g2648 ( 
.A(n_2406),
.Y(n_2648)
);

NAND2xp33_ASAP7_75t_SL g2649 ( 
.A(n_2238),
.B(n_1142),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2097),
.A2(n_1486),
.B1(n_1487),
.B2(n_1483),
.Y(n_2650)
);

BUFx3_ASAP7_75t_L g2651 ( 
.A(n_2086),
.Y(n_2651)
);

INVx3_ASAP7_75t_L g2652 ( 
.A(n_2209),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2160),
.Y(n_2653)
);

BUFx2_ASAP7_75t_L g2654 ( 
.A(n_2425),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2223),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2115),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2160),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2163),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2163),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2425),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2115),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_2214),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2173),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2173),
.Y(n_2664)
);

HB1xp67_ASAP7_75t_L g2665 ( 
.A(n_2421),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2214),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2199),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2199),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2200),
.Y(n_2669)
);

HB1xp67_ASAP7_75t_L g2670 ( 
.A(n_2082),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2289),
.B(n_1167),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2200),
.Y(n_2672)
);

BUFx2_ASAP7_75t_L g2673 ( 
.A(n_2433),
.Y(n_2673)
);

BUFx6f_ASAP7_75t_SL g2674 ( 
.A(n_2406),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2206),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2206),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2216),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2218),
.B(n_1167),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2216),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2217),
.Y(n_2680)
);

AND2x4_ASAP7_75t_L g2681 ( 
.A(n_2026),
.B(n_1491),
.Y(n_2681)
);

INVx3_ASAP7_75t_L g2682 ( 
.A(n_2223),
.Y(n_2682)
);

BUFx2_ASAP7_75t_L g2683 ( 
.A(n_2433),
.Y(n_2683)
);

NOR2xp33_ASAP7_75t_L g2684 ( 
.A(n_2156),
.B(n_819),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2217),
.Y(n_2685)
);

OAI22xp5_ASAP7_75t_SL g2686 ( 
.A1(n_2048),
.A2(n_1910),
.B1(n_1927),
.B2(n_1900),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2228),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2026),
.B(n_1492),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2228),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2232),
.Y(n_2690)
);

XOR2xp5_ASAP7_75t_L g2691 ( 
.A(n_2069),
.B(n_1928),
.Y(n_2691)
);

BUFx6f_ASAP7_75t_L g2692 ( 
.A(n_2214),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_2214),
.B(n_931),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2232),
.Y(n_2694)
);

CKINVDCx20_ASAP7_75t_R g2695 ( 
.A(n_2069),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2235),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2235),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2225),
.B(n_1169),
.Y(n_2698)
);

BUFx6f_ASAP7_75t_SL g2699 ( 
.A(n_2300),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2227),
.B(n_2097),
.Y(n_2700)
);

AND2x2_ASAP7_75t_L g2701 ( 
.A(n_2326),
.B(n_1493),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2241),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2433),
.Y(n_2703)
);

AND2x6_ASAP7_75t_L g2704 ( 
.A(n_2259),
.B(n_931),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2097),
.B(n_1169),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2241),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2242),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2242),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2244),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2244),
.Y(n_2710)
);

INVx3_ASAP7_75t_L g2711 ( 
.A(n_2239),
.Y(n_2711)
);

INVxp67_ASAP7_75t_L g2712 ( 
.A(n_2404),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2245),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2245),
.Y(n_2714)
);

AOI22xp5_ASAP7_75t_L g2715 ( 
.A1(n_2097),
.A2(n_1496),
.B1(n_1497),
.B2(n_1495),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2210),
.Y(n_2716)
);

INVx3_ASAP7_75t_L g2717 ( 
.A(n_2239),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2252),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2252),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2231),
.Y(n_2720)
);

AND2x4_ASAP7_75t_L g2721 ( 
.A(n_2026),
.B(n_1498),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2117),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2326),
.B(n_1501),
.Y(n_2723)
);

INVx1_ASAP7_75t_SL g2724 ( 
.A(n_2395),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2117),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2233),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2234),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2237),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2260),
.B(n_1502),
.Y(n_2729)
);

INVxp67_ASAP7_75t_L g2730 ( 
.A(n_2404),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2246),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2262),
.B(n_1503),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2247),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2122),
.Y(n_2734)
);

AND2x2_ASAP7_75t_L g2735 ( 
.A(n_2349),
.B(n_1504),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2122),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_SL g2737 ( 
.A(n_2349),
.B(n_935),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2248),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2249),
.Y(n_2739)
);

INVx2_ASAP7_75t_L g2740 ( 
.A(n_2123),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2251),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2210),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2253),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2254),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2255),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2256),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2349),
.B(n_1505),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2257),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2377),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2377),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2377),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2123),
.Y(n_2752)
);

AND2x4_ASAP7_75t_L g2753 ( 
.A(n_2363),
.B(n_1506),
.Y(n_2753)
);

INVxp67_ASAP7_75t_L g2754 ( 
.A(n_2429),
.Y(n_2754)
);

BUFx6f_ASAP7_75t_L g2755 ( 
.A(n_2054),
.Y(n_2755)
);

AND2x4_ASAP7_75t_L g2756 ( 
.A(n_2086),
.B(n_1507),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2062),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2088),
.B(n_1508),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2087),
.Y(n_2759)
);

NAND2xp33_ASAP7_75t_SL g2760 ( 
.A(n_2328),
.B(n_935),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2101),
.Y(n_2761)
);

BUFx6f_ASAP7_75t_L g2762 ( 
.A(n_2054),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2139),
.Y(n_2763)
);

INVx2_ASAP7_75t_L g2764 ( 
.A(n_2151),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2143),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2161),
.Y(n_2766)
);

NOR2xp33_ASAP7_75t_L g2767 ( 
.A(n_2038),
.B(n_820),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2215),
.Y(n_2768)
);

INVx3_ASAP7_75t_L g2769 ( 
.A(n_2056),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2151),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2056),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2109),
.Y(n_2772)
);

OA21x2_ASAP7_75t_L g2773 ( 
.A1(n_2109),
.A2(n_2240),
.B(n_2224),
.Y(n_2773)
);

OAI22xp5_ASAP7_75t_SL g2774 ( 
.A1(n_2114),
.A2(n_1928),
.B1(n_827),
.B2(n_828),
.Y(n_2774)
);

INVx3_ASAP7_75t_L g2775 ( 
.A(n_2056),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2383),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2056),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2383),
.Y(n_2778)
);

AND2x4_ASAP7_75t_L g2779 ( 
.A(n_2091),
.B(n_2294),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2068),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2054),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2068),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2068),
.Y(n_2783)
);

BUFx2_ASAP7_75t_L g2784 ( 
.A(n_2435),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2263),
.B(n_1515),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2383),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2068),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2176),
.Y(n_2788)
);

NAND2xp5_ASAP7_75t_L g2789 ( 
.A(n_2294),
.B(n_1516),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2091),
.B(n_1517),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2071),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2071),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2071),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2176),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2194),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2071),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2428),
.Y(n_2797)
);

AOI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2084),
.A2(n_1520),
.B1(n_1521),
.B2(n_1518),
.Y(n_2798)
);

BUFx6f_ASAP7_75t_L g2799 ( 
.A(n_2054),
.Y(n_2799)
);

INVx3_ASAP7_75t_L g2800 ( 
.A(n_2090),
.Y(n_2800)
);

INVx1_ASAP7_75t_SL g2801 ( 
.A(n_2396),
.Y(n_2801)
);

BUFx6f_ASAP7_75t_L g2802 ( 
.A(n_2055),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2328),
.B(n_2198),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2090),
.Y(n_2804)
);

BUFx2_ASAP7_75t_L g2805 ( 
.A(n_2435),
.Y(n_2805)
);

AND2x4_ASAP7_75t_L g2806 ( 
.A(n_2162),
.B(n_1522),
.Y(n_2806)
);

AND3x1_ASAP7_75t_L g2807 ( 
.A(n_2429),
.B(n_1058),
.C(n_1053),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2428),
.Y(n_2808)
);

OAI22xp5_ASAP7_75t_SL g2809 ( 
.A1(n_2114),
.A2(n_829),
.B1(n_834),
.B2(n_824),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2428),
.Y(n_2810)
);

INVx3_ASAP7_75t_L g2811 ( 
.A(n_2090),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2090),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_2093),
.Y(n_2813)
);

NAND2xp5_ASAP7_75t_SL g2814 ( 
.A(n_2038),
.B(n_935),
.Y(n_2814)
);

BUFx2_ASAP7_75t_L g2815 ( 
.A(n_2435),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2181),
.B(n_2220),
.Y(n_2816)
);

HB1xp67_ASAP7_75t_L g2817 ( 
.A(n_2368),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2093),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2250),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2250),
.Y(n_2820)
);

AOI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2084),
.A2(n_1525),
.B1(n_1527),
.B2(n_1524),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2093),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2102),
.B(n_996),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2250),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2250),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2093),
.Y(n_2826)
);

INVx1_ASAP7_75t_SL g2827 ( 
.A(n_2135),
.Y(n_2827)
);

CKINVDCx11_ASAP7_75t_R g2828 ( 
.A(n_2135),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2212),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2119),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2142),
.Y(n_2831)
);

INVxp67_ASAP7_75t_L g2832 ( 
.A(n_2183),
.Y(n_2832)
);

BUFx6f_ASAP7_75t_L g2833 ( 
.A(n_2055),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2055),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_SL g2835 ( 
.A(n_2369),
.B(n_996),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2119),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2119),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2119),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2142),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2142),
.Y(n_2840)
);

BUFx6f_ASAP7_75t_L g2841 ( 
.A(n_2055),
.Y(n_2841)
);

BUFx6f_ASAP7_75t_L g2842 ( 
.A(n_2142),
.Y(n_2842)
);

OAI22xp5_ASAP7_75t_L g2843 ( 
.A1(n_2041),
.A2(n_838),
.B1(n_839),
.B2(n_835),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2119),
.Y(n_2844)
);

OAI22xp5_ASAP7_75t_L g2845 ( 
.A1(n_2181),
.A2(n_2220),
.B1(n_2118),
.B2(n_2337),
.Y(n_2845)
);

INVxp67_ASAP7_75t_L g2846 ( 
.A(n_2213),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2364),
.Y(n_2847)
);

BUFx6f_ASAP7_75t_L g2848 ( 
.A(n_2167),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_SL g2849 ( 
.A(n_2152),
.B(n_2134),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2296),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2167),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2342),
.B(n_1528),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2118),
.A2(n_842),
.B1(n_843),
.B2(n_840),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2175),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2296),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2177),
.B(n_1531),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2182),
.B(n_1533),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2354),
.A2(n_1539),
.B1(n_1541),
.B2(n_1536),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2167),
.Y(n_2859)
);

OAI22xp5_ASAP7_75t_SL g2860 ( 
.A1(n_2175),
.A2(n_848),
.B1(n_850),
.B2(n_846),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2438),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2788),
.B(n_2354),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2453),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2489),
.Y(n_2864)
);

BUFx3_ASAP7_75t_L g2865 ( 
.A(n_2847),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2440),
.Y(n_2866)
);

INVxp67_ASAP7_75t_SL g2867 ( 
.A(n_2448),
.Y(n_2867)
);

XOR2xp5_ASAP7_75t_L g2868 ( 
.A(n_2574),
.B(n_2293),
.Y(n_2868)
);

INVx4_ASAP7_75t_L g2869 ( 
.A(n_2716),
.Y(n_2869)
);

OR2x2_ASAP7_75t_L g2870 ( 
.A(n_2724),
.B(n_2412),
.Y(n_2870)
);

INVx6_ASAP7_75t_L g2871 ( 
.A(n_2552),
.Y(n_2871)
);

NOR2xp33_ASAP7_75t_L g2872 ( 
.A(n_2514),
.B(n_2274),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2443),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2441),
.B(n_2333),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2794),
.B(n_2354),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2757),
.B(n_2354),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2444),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2445),
.Y(n_2878)
);

NOR2xp33_ASAP7_75t_L g2879 ( 
.A(n_2541),
.B(n_2816),
.Y(n_2879)
);

NAND2xp33_ASAP7_75t_L g2880 ( 
.A(n_2465),
.B(n_2354),
.Y(n_2880)
);

CKINVDCx20_ASAP7_75t_R g2881 ( 
.A(n_2547),
.Y(n_2881)
);

AND2x4_ASAP7_75t_L g2882 ( 
.A(n_2491),
.B(n_2492),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2446),
.Y(n_2883)
);

INVx3_ASAP7_75t_L g2884 ( 
.A(n_2453),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2491),
.B(n_2261),
.Y(n_2885)
);

AND2x4_ASAP7_75t_L g2886 ( 
.A(n_2492),
.B(n_2261),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_2816),
.A2(n_1003),
.B1(n_1027),
.B2(n_996),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2759),
.B(n_2342),
.Y(n_2888)
);

INVxp67_ASAP7_75t_SL g2889 ( 
.A(n_2448),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2814),
.A2(n_1003),
.B1(n_1033),
.B2(n_1027),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2455),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2515),
.B(n_2563),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2457),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2814),
.A2(n_1003),
.B1(n_1033),
.B2(n_1027),
.Y(n_2894)
);

CKINVDCx20_ASAP7_75t_R g2895 ( 
.A(n_2525),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2489),
.Y(n_2896)
);

AND2x6_ASAP7_75t_L g2897 ( 
.A(n_2544),
.B(n_2266),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2515),
.B(n_2187),
.Y(n_2898)
);

BUFx6f_ASAP7_75t_L g2899 ( 
.A(n_2594),
.Y(n_2899)
);

INVxp67_ASAP7_75t_SL g2900 ( 
.A(n_2450),
.Y(n_2900)
);

INVx1_ASAP7_75t_L g2901 ( 
.A(n_2636),
.Y(n_2901)
);

AO22x2_ASAP7_75t_L g2902 ( 
.A1(n_2845),
.A2(n_2364),
.B1(n_2382),
.B2(n_2372),
.Y(n_2902)
);

INVxp67_ASAP7_75t_SL g2903 ( 
.A(n_2450),
.Y(n_2903)
);

BUFx3_ASAP7_75t_L g2904 ( 
.A(n_2847),
.Y(n_2904)
);

INVx4_ASAP7_75t_L g2905 ( 
.A(n_2716),
.Y(n_2905)
);

OR2x6_ASAP7_75t_L g2906 ( 
.A(n_2510),
.B(n_2368),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2496),
.Y(n_2907)
);

BUFx3_ASAP7_75t_L g2908 ( 
.A(n_2552),
.Y(n_2908)
);

INVxp67_ASAP7_75t_SL g2909 ( 
.A(n_2451),
.Y(n_2909)
);

INVx2_ASAP7_75t_L g2910 ( 
.A(n_2496),
.Y(n_2910)
);

CKINVDCx5p33_ASAP7_75t_R g2911 ( 
.A(n_2828),
.Y(n_2911)
);

AND2x4_ASAP7_75t_L g2912 ( 
.A(n_2594),
.B(n_2264),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2712),
.B(n_2281),
.Y(n_2913)
);

BUFx2_ASAP7_75t_L g2914 ( 
.A(n_2437),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2637),
.Y(n_2915)
);

NOR2x1p5_ASAP7_75t_L g2916 ( 
.A(n_2651),
.B(n_2310),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2638),
.Y(n_2917)
);

INVx1_ASAP7_75t_SL g2918 ( 
.A(n_2442),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2641),
.Y(n_2919)
);

AOI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2779),
.A2(n_2767),
.B1(n_2439),
.B2(n_2529),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2730),
.B(n_2281),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2643),
.Y(n_2922)
);

BUFx6f_ASAP7_75t_L g2923 ( 
.A(n_2716),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2656),
.Y(n_2924)
);

BUFx6f_ASAP7_75t_L g2925 ( 
.A(n_2716),
.Y(n_2925)
);

HB1xp67_ASAP7_75t_L g2926 ( 
.A(n_2449),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_SL g2927 ( 
.A(n_2742),
.B(n_2300),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2661),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2441),
.B(n_2333),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2452),
.B(n_2336),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_2502),
.Y(n_2931)
);

NAND3xp33_ASAP7_75t_L g2932 ( 
.A(n_2767),
.B(n_2380),
.C(n_2106),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2502),
.Y(n_2933)
);

BUFx3_ASAP7_75t_L g2934 ( 
.A(n_2552),
.Y(n_2934)
);

INVx2_ASAP7_75t_L g2935 ( 
.A(n_2511),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2452),
.B(n_2336),
.Y(n_2936)
);

INVx5_ASAP7_75t_L g2937 ( 
.A(n_2544),
.Y(n_2937)
);

INVx1_ASAP7_75t_SL g2938 ( 
.A(n_2801),
.Y(n_2938)
);

AND2x4_ASAP7_75t_L g2939 ( 
.A(n_2651),
.B(n_2264),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2453),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2618),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2563),
.B(n_2761),
.Y(n_2942)
);

OR2x6_ASAP7_75t_L g2943 ( 
.A(n_2510),
.B(n_2368),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2742),
.B(n_2300),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2511),
.Y(n_2945)
);

INVxp67_ASAP7_75t_L g2946 ( 
.A(n_2464),
.Y(n_2946)
);

AOI22xp5_ASAP7_75t_L g2947 ( 
.A1(n_2779),
.A2(n_2309),
.B1(n_2322),
.B2(n_2306),
.Y(n_2947)
);

CKINVDCx5p33_ASAP7_75t_R g2948 ( 
.A(n_2828),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2512),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_2589),
.Y(n_2950)
);

NOR2xp33_ASAP7_75t_L g2951 ( 
.A(n_2754),
.B(n_2348),
.Y(n_2951)
);

INVx3_ASAP7_75t_L g2952 ( 
.A(n_2580),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2618),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_SL g2954 ( 
.A(n_2742),
.B(n_2300),
.Y(n_2954)
);

OR2x2_ASAP7_75t_L g2955 ( 
.A(n_2589),
.B(n_2471),
.Y(n_2955)
);

INVx3_ASAP7_75t_L g2956 ( 
.A(n_2580),
.Y(n_2956)
);

HB1xp67_ASAP7_75t_L g2957 ( 
.A(n_2703),
.Y(n_2957)
);

BUFx3_ASAP7_75t_L g2958 ( 
.A(n_2817),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2763),
.B(n_2187),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2622),
.Y(n_2960)
);

CKINVDCx5p33_ASAP7_75t_R g2961 ( 
.A(n_2699),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2765),
.B(n_2134),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2622),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2631),
.Y(n_2964)
);

AOI22xp5_ASAP7_75t_L g2965 ( 
.A1(n_2779),
.A2(n_2309),
.B1(n_2322),
.B2(n_2306),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2631),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_L g2967 ( 
.A1(n_2749),
.A2(n_1033),
.B1(n_1135),
.B2(n_1047),
.Y(n_2967)
);

INVx1_ASAP7_75t_SL g2968 ( 
.A(n_2493),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2512),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2517),
.Y(n_2970)
);

AND2x2_ASAP7_75t_SL g2971 ( 
.A(n_2753),
.B(n_2368),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2766),
.B(n_2272),
.Y(n_2972)
);

INVx3_ASAP7_75t_L g2973 ( 
.A(n_2580),
.Y(n_2973)
);

NOR2x1p5_ASAP7_75t_L g2974 ( 
.A(n_2850),
.B(n_2310),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_SL g2975 ( 
.A(n_2742),
.B(n_2311),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_2829),
.B(n_2272),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2581),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2632),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_SL g2979 ( 
.A(n_2832),
.B(n_2311),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2583),
.B(n_2273),
.Y(n_2980)
);

NOR2xp33_ASAP7_75t_L g2981 ( 
.A(n_2597),
.B(n_2348),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2758),
.B(n_2273),
.Y(n_2982)
);

NOR2xp33_ASAP7_75t_L g2983 ( 
.A(n_2604),
.B(n_2359),
.Y(n_2983)
);

CKINVDCx8_ASAP7_75t_R g2984 ( 
.A(n_2519),
.Y(n_2984)
);

INVx3_ASAP7_75t_L g2985 ( 
.A(n_2581),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2758),
.B(n_2276),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2464),
.B(n_2359),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2632),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2461),
.B(n_2311),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2653),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2653),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2657),
.Y(n_2992)
);

INVxp33_ASAP7_75t_L g2993 ( 
.A(n_2670),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_SL g2994 ( 
.A(n_2461),
.B(n_2311),
.Y(n_2994)
);

NAND2xp5_ASAP7_75t_SL g2995 ( 
.A(n_2461),
.B(n_2320),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2657),
.Y(n_2996)
);

CKINVDCx5p33_ASAP7_75t_R g2997 ( 
.A(n_2699),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2501),
.B(n_2360),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_SL g2999 ( 
.A(n_2476),
.B(n_2320),
.Y(n_2999)
);

INVx4_ASAP7_75t_L g3000 ( 
.A(n_2465),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2565),
.A2(n_2376),
.B1(n_2332),
.B2(n_2352),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2517),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2658),
.Y(n_3003)
);

NOR2xp33_ASAP7_75t_L g3004 ( 
.A(n_2568),
.B(n_2360),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2476),
.B(n_2320),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2520),
.Y(n_3006)
);

AOI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2439),
.A2(n_2332),
.B1(n_2352),
.B2(n_2331),
.Y(n_3007)
);

AND2x6_ASAP7_75t_L g3008 ( 
.A(n_2544),
.B(n_2266),
.Y(n_3008)
);

OR2x2_ASAP7_75t_L g3009 ( 
.A(n_2487),
.B(n_2419),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2795),
.B(n_2276),
.Y(n_3010)
);

INVxp67_ASAP7_75t_L g3011 ( 
.A(n_2475),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2658),
.Y(n_3012)
);

INVx3_ASAP7_75t_L g3013 ( 
.A(n_2581),
.Y(n_3013)
);

AND2x6_ASAP7_75t_L g3014 ( 
.A(n_2544),
.B(n_2267),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2659),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2520),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2659),
.Y(n_3017)
);

INVx1_ASAP7_75t_SL g3018 ( 
.A(n_2487),
.Y(n_3018)
);

INVx1_ASAP7_75t_SL g3019 ( 
.A(n_2827),
.Y(n_3019)
);

CKINVDCx20_ASAP7_75t_R g3020 ( 
.A(n_2525),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2663),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2781),
.Y(n_3022)
);

NOR2xp33_ASAP7_75t_L g3023 ( 
.A(n_2602),
.B(n_2258),
.Y(n_3023)
);

INVx4_ASAP7_75t_L g3024 ( 
.A(n_2465),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2527),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2663),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2527),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2625),
.B(n_2331),
.Y(n_3028)
);

INVx1_ASAP7_75t_SL g3029 ( 
.A(n_2480),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2577),
.B(n_2280),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2630),
.B(n_2356),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2577),
.B(n_2280),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2676),
.Y(n_3033)
);

HB1xp67_ASAP7_75t_L g3034 ( 
.A(n_2519),
.Y(n_3034)
);

BUFx2_ASAP7_75t_L g3035 ( 
.A(n_2550),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2528),
.Y(n_3036)
);

INVx4_ASAP7_75t_L g3037 ( 
.A(n_2465),
.Y(n_3037)
);

NAND2x1p5_ASAP7_75t_L g3038 ( 
.A(n_2470),
.B(n_2320),
.Y(n_3038)
);

AND2x4_ASAP7_75t_L g3039 ( 
.A(n_2756),
.B(n_2790),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2475),
.B(n_2329),
.Y(n_3040)
);

BUFx3_ASAP7_75t_L g3041 ( 
.A(n_2855),
.Y(n_3041)
);

NOR2xp33_ASAP7_75t_L g3042 ( 
.A(n_2665),
.B(n_2356),
.Y(n_3042)
);

NOR2xp33_ASAP7_75t_SL g3043 ( 
.A(n_2500),
.B(n_2243),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2528),
.Y(n_3044)
);

BUFx6f_ASAP7_75t_L g3045 ( 
.A(n_2781),
.Y(n_3045)
);

BUFx6f_ASAP7_75t_L g3046 ( 
.A(n_2781),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2676),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2508),
.B(n_2329),
.Y(n_3048)
);

BUFx6f_ASAP7_75t_L g3049 ( 
.A(n_2781),
.Y(n_3049)
);

BUFx3_ASAP7_75t_L g3050 ( 
.A(n_2695),
.Y(n_3050)
);

AO22x2_ASAP7_75t_L g3051 ( 
.A1(n_2797),
.A2(n_2382),
.B1(n_2397),
.B2(n_2372),
.Y(n_3051)
);

OAI21xp33_ASAP7_75t_L g3052 ( 
.A1(n_2554),
.A2(n_2361),
.B(n_2298),
.Y(n_3052)
);

NOR2xp33_ASAP7_75t_L g3053 ( 
.A(n_2554),
.B(n_2684),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2679),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2578),
.B(n_2040),
.Y(n_3055)
);

BUFx6f_ASAP7_75t_L g3056 ( 
.A(n_2781),
.Y(n_3056)
);

INVx4_ASAP7_75t_L g3057 ( 
.A(n_2470),
.Y(n_3057)
);

AOI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2529),
.A2(n_2270),
.B1(n_2271),
.B2(n_2269),
.Y(n_3058)
);

BUFx4f_ASAP7_75t_L g3059 ( 
.A(n_2522),
.Y(n_3059)
);

AND2x6_ASAP7_75t_L g3060 ( 
.A(n_2544),
.B(n_2267),
.Y(n_3060)
);

BUFx6f_ASAP7_75t_L g3061 ( 
.A(n_2799),
.Y(n_3061)
);

NAND3x1_ASAP7_75t_L g3062 ( 
.A(n_2684),
.B(n_2366),
.C(n_2381),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_L g3063 ( 
.A(n_2578),
.B(n_2040),
.Y(n_3063)
);

BUFx2_ASAP7_75t_L g3064 ( 
.A(n_2550),
.Y(n_3064)
);

INVxp33_ASAP7_75t_SL g3065 ( 
.A(n_2691),
.Y(n_3065)
);

NOR2xp33_ASAP7_75t_L g3066 ( 
.A(n_2572),
.B(n_2305),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2679),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2530),
.B(n_2315),
.Y(n_3068)
);

INVx2_ASAP7_75t_L g3069 ( 
.A(n_2532),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2532),
.Y(n_3070)
);

INVxp33_ASAP7_75t_L g3071 ( 
.A(n_2691),
.Y(n_3071)
);

AND2x6_ASAP7_75t_L g3072 ( 
.A(n_2570),
.B(n_2329),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_2695),
.Y(n_3073)
);

AND2x6_ASAP7_75t_L g3074 ( 
.A(n_2570),
.B(n_2329),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2486),
.B(n_2152),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2799),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2536),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2694),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_2530),
.B(n_2319),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2536),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_2699),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2486),
.B(n_2152),
.Y(n_3082)
);

BUFx2_ASAP7_75t_L g3083 ( 
.A(n_2561),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2545),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2545),
.Y(n_3085)
);

NOR2xp33_ASAP7_75t_L g3086 ( 
.A(n_2543),
.B(n_2321),
.Y(n_3086)
);

INVx1_ASAP7_75t_SL g3087 ( 
.A(n_2854),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2694),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_2486),
.B(n_2152),
.Y(n_3089)
);

AND2x4_ASAP7_75t_L g3090 ( 
.A(n_2756),
.B(n_2330),
.Y(n_3090)
);

AND2x4_ASAP7_75t_L g3091 ( 
.A(n_2756),
.B(n_2330),
.Y(n_3091)
);

INVx3_ASAP7_75t_L g3092 ( 
.A(n_2609),
.Y(n_3092)
);

INVx2_ASAP7_75t_L g3093 ( 
.A(n_2546),
.Y(n_3093)
);

BUFx6f_ASAP7_75t_SL g3094 ( 
.A(n_2790),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_2543),
.B(n_2325),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2708),
.Y(n_3096)
);

NAND2xp5_ASAP7_75t_L g3097 ( 
.A(n_2516),
.B(n_2275),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2516),
.B(n_2299),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2708),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2714),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2714),
.Y(n_3101)
);

NOR2xp33_ASAP7_75t_L g3102 ( 
.A(n_2846),
.B(n_2343),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2546),
.Y(n_3103)
);

BUFx6f_ASAP7_75t_L g3104 ( 
.A(n_2799),
.Y(n_3104)
);

BUFx10_ASAP7_75t_L g3105 ( 
.A(n_2790),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2516),
.B(n_2299),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2722),
.Y(n_3107)
);

AND3x2_ASAP7_75t_L g3108 ( 
.A(n_2561),
.B(n_2365),
.C(n_2317),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2722),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2725),
.Y(n_3110)
);

BUFx3_ASAP7_75t_L g3111 ( 
.A(n_2854),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2523),
.B(n_2167),
.Y(n_3112)
);

AO21x2_ASAP7_75t_L g3113 ( 
.A1(n_2705),
.A2(n_2361),
.B(n_2298),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2523),
.B(n_2344),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2476),
.B(n_2330),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2523),
.B(n_2346),
.Y(n_3116)
);

HB1xp67_ASAP7_75t_L g3117 ( 
.A(n_2606),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2609),
.B(n_2350),
.Y(n_3118)
);

INVx3_ASAP7_75t_L g3119 ( 
.A(n_2609),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_2508),
.B(n_2355),
.Y(n_3120)
);

BUFx10_ASAP7_75t_L g3121 ( 
.A(n_2806),
.Y(n_3121)
);

INVx4_ASAP7_75t_L g3122 ( 
.A(n_2470),
.Y(n_3122)
);

CKINVDCx20_ASAP7_75t_R g3123 ( 
.A(n_2574),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2803),
.B(n_2168),
.Y(n_3124)
);

AOI22xp33_ASAP7_75t_L g3125 ( 
.A1(n_2750),
.A2(n_2751),
.B1(n_2760),
.B2(n_2776),
.Y(n_3125)
);

AOI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2835),
.A2(n_2277),
.B1(n_2290),
.B2(n_2279),
.Y(n_3126)
);

BUFx10_ASAP7_75t_L g3127 ( 
.A(n_2806),
.Y(n_3127)
);

NOR2xp33_ASAP7_75t_L g3128 ( 
.A(n_2606),
.B(n_2614),
.Y(n_3128)
);

BUFx4f_ASAP7_75t_L g3129 ( 
.A(n_2522),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_2518),
.B(n_2330),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2725),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2856),
.B(n_2292),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2856),
.B(n_2340),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_SL g3134 ( 
.A(n_2518),
.B(n_2340),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2734),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2760),
.A2(n_1135),
.B1(n_1140),
.B2(n_1047),
.Y(n_3136)
);

BUFx2_ASAP7_75t_L g3137 ( 
.A(n_2614),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2734),
.Y(n_3138)
);

INVx2_ASAP7_75t_L g3139 ( 
.A(n_2548),
.Y(n_3139)
);

NOR2xp33_ASAP7_75t_L g3140 ( 
.A(n_2623),
.B(n_2340),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_2623),
.B(n_2340),
.Y(n_3141)
);

AND2x6_ASAP7_75t_L g3142 ( 
.A(n_2573),
.B(n_2454),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_2778),
.A2(n_1135),
.B1(n_1140),
.B2(n_1047),
.Y(n_3143)
);

OR2x2_ASAP7_75t_L g3144 ( 
.A(n_2654),
.B(n_2397),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2736),
.Y(n_3145)
);

CKINVDCx5p33_ASAP7_75t_R g3146 ( 
.A(n_2599),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2654),
.B(n_2341),
.Y(n_3147)
);

INVx3_ASAP7_75t_L g3148 ( 
.A(n_2613),
.Y(n_3148)
);

BUFx3_ASAP7_75t_L g3149 ( 
.A(n_2660),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_SL g3150 ( 
.A(n_2518),
.B(n_2341),
.Y(n_3150)
);

CKINVDCx20_ASAP7_75t_R g3151 ( 
.A(n_2644),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_2736),
.Y(n_3152)
);

INVx3_ASAP7_75t_L g3153 ( 
.A(n_2613),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2857),
.B(n_2052),
.Y(n_3154)
);

INVx4_ASAP7_75t_L g3155 ( 
.A(n_2470),
.Y(n_3155)
);

AND2x4_ASAP7_75t_L g3156 ( 
.A(n_2681),
.B(n_2341),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2740),
.Y(n_3157)
);

CKINVDCx5p33_ASAP7_75t_R g3158 ( 
.A(n_2686),
.Y(n_3158)
);

CKINVDCx5p33_ASAP7_75t_R g3159 ( 
.A(n_2588),
.Y(n_3159)
);

HB1xp67_ASAP7_75t_L g3160 ( 
.A(n_2660),
.Y(n_3160)
);

AND2x4_ASAP7_75t_L g3161 ( 
.A(n_2681),
.B(n_2341),
.Y(n_3161)
);

INVx2_ASAP7_75t_SL g3162 ( 
.A(n_2608),
.Y(n_3162)
);

INVx2_ASAP7_75t_L g3163 ( 
.A(n_2548),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2740),
.Y(n_3164)
);

NAND2xp33_ASAP7_75t_L g3165 ( 
.A(n_2484),
.B(n_2498),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2752),
.Y(n_3166)
);

AND2x2_ASAP7_75t_L g3167 ( 
.A(n_2857),
.B(n_2608),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2752),
.Y(n_3168)
);

INVx5_ASAP7_75t_L g3169 ( 
.A(n_2617),
.Y(n_3169)
);

INVx4_ASAP7_75t_L g3170 ( 
.A(n_2484),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2764),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_SL g3172 ( 
.A(n_2579),
.B(n_2357),
.Y(n_3172)
);

INVx5_ASAP7_75t_L g3173 ( 
.A(n_2617),
.Y(n_3173)
);

INVx4_ASAP7_75t_L g3174 ( 
.A(n_2484),
.Y(n_3174)
);

NOR2xp33_ASAP7_75t_L g3175 ( 
.A(n_2673),
.B(n_2357),
.Y(n_3175)
);

AND2x6_ASAP7_75t_L g3176 ( 
.A(n_2573),
.B(n_2357),
.Y(n_3176)
);

NOR2xp33_ASAP7_75t_L g3177 ( 
.A(n_2673),
.B(n_2357),
.Y(n_3177)
);

INVx4_ASAP7_75t_L g3178 ( 
.A(n_2484),
.Y(n_3178)
);

NOR2xp33_ASAP7_75t_L g3179 ( 
.A(n_2683),
.B(n_2258),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2616),
.B(n_2140),
.Y(n_3180)
);

INVx2_ASAP7_75t_SL g3181 ( 
.A(n_2616),
.Y(n_3181)
);

AND2x4_ASAP7_75t_L g3182 ( 
.A(n_2681),
.B(n_2265),
.Y(n_3182)
);

BUFx6f_ASAP7_75t_L g3183 ( 
.A(n_2799),
.Y(n_3183)
);

INVx2_ASAP7_75t_L g3184 ( 
.A(n_2562),
.Y(n_3184)
);

INVx4_ASAP7_75t_L g3185 ( 
.A(n_2498),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2764),
.Y(n_3186)
);

AND2x2_ASAP7_75t_SL g3187 ( 
.A(n_2753),
.B(n_2384),
.Y(n_3187)
);

AND2x2_ASAP7_75t_L g3188 ( 
.A(n_2639),
.B(n_2278),
.Y(n_3188)
);

AND2x4_ASAP7_75t_L g3189 ( 
.A(n_2688),
.B(n_2265),
.Y(n_3189)
);

BUFx6f_ASAP7_75t_L g3190 ( 
.A(n_2799),
.Y(n_3190)
);

BUFx3_ASAP7_75t_L g3191 ( 
.A(n_2683),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2639),
.B(n_2642),
.Y(n_3192)
);

NOR2xp33_ASAP7_75t_L g3193 ( 
.A(n_2784),
.B(n_2297),
.Y(n_3193)
);

BUFx4f_ASAP7_75t_L g3194 ( 
.A(n_2522),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2770),
.Y(n_3195)
);

AND2x4_ASAP7_75t_L g3196 ( 
.A(n_2688),
.B(n_2265),
.Y(n_3196)
);

INVx3_ASAP7_75t_L g3197 ( 
.A(n_2613),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_2770),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_2562),
.Y(n_3199)
);

INVx4_ASAP7_75t_L g3200 ( 
.A(n_2498),
.Y(n_3200)
);

NAND2xp33_ASAP7_75t_L g3201 ( 
.A(n_2498),
.B(n_2196),
.Y(n_3201)
);

INVxp67_ASAP7_75t_SL g3202 ( 
.A(n_2451),
.Y(n_3202)
);

INVx3_ASAP7_75t_L g3203 ( 
.A(n_2626),
.Y(n_3203)
);

BUFx6f_ASAP7_75t_L g3204 ( 
.A(n_2755),
.Y(n_3204)
);

INVx3_ASAP7_75t_L g3205 ( 
.A(n_2626),
.Y(n_3205)
);

BUFx6f_ASAP7_75t_L g3206 ( 
.A(n_2755),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_2784),
.Y(n_3207)
);

NAND2xp5_ASAP7_75t_L g3208 ( 
.A(n_2626),
.B(n_2627),
.Y(n_3208)
);

BUFx2_ASAP7_75t_L g3209 ( 
.A(n_2805),
.Y(n_3209)
);

INVx1_ASAP7_75t_SL g3210 ( 
.A(n_2805),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2664),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2667),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_2627),
.B(n_2052),
.Y(n_3213)
);

NOR2xp33_ASAP7_75t_L g3214 ( 
.A(n_2815),
.B(n_2301),
.Y(n_3214)
);

INVx4_ASAP7_75t_SL g3215 ( 
.A(n_2509),
.Y(n_3215)
);

AND2x4_ASAP7_75t_L g3216 ( 
.A(n_2688),
.B(n_2721),
.Y(n_3216)
);

BUFx3_ASAP7_75t_L g3217 ( 
.A(n_2815),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_2567),
.Y(n_3218)
);

AND2x6_ASAP7_75t_L g3219 ( 
.A(n_2454),
.B(n_2047),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2627),
.B(n_2302),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_2721),
.B(n_2050),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_2642),
.B(n_2226),
.Y(n_3222)
);

INVx4_ASAP7_75t_L g3223 ( 
.A(n_2503),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2567),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2668),
.Y(n_3225)
);

BUFx6f_ASAP7_75t_L g3226 ( 
.A(n_2755),
.Y(n_3226)
);

INVx1_ASAP7_75t_L g3227 ( 
.A(n_2669),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2672),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_SL g3229 ( 
.A(n_2579),
.B(n_2196),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2675),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2677),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_2718),
.Y(n_3232)
);

INVx1_ASAP7_75t_SL g3233 ( 
.A(n_2701),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_2652),
.B(n_2374),
.Y(n_3234)
);

BUFx6f_ASAP7_75t_L g3235 ( 
.A(n_2755),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_2680),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2718),
.Y(n_3237)
);

INVx4_ASAP7_75t_L g3238 ( 
.A(n_2503),
.Y(n_3238)
);

BUFx4f_ASAP7_75t_L g3239 ( 
.A(n_2522),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2652),
.B(n_2411),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2685),
.Y(n_3241)
);

NAND2xp5_ASAP7_75t_SL g3242 ( 
.A(n_2579),
.B(n_2203),
.Y(n_3242)
);

OR2x6_ASAP7_75t_L g3243 ( 
.A(n_2459),
.B(n_2384),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2687),
.Y(n_3244)
);

INVx3_ASAP7_75t_L g3245 ( 
.A(n_2652),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_2701),
.B(n_2226),
.Y(n_3246)
);

INVx2_ASAP7_75t_L g3247 ( 
.A(n_2719),
.Y(n_3247)
);

AND2x4_ASAP7_75t_L g3248 ( 
.A(n_2721),
.B(n_2628),
.Y(n_3248)
);

INVx2_ASAP7_75t_L g3249 ( 
.A(n_2719),
.Y(n_3249)
);

INVx2_ASAP7_75t_L g3250 ( 
.A(n_2582),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2582),
.Y(n_3251)
);

INVx1_ASAP7_75t_SL g3252 ( 
.A(n_2723),
.Y(n_3252)
);

AND2x4_ASAP7_75t_L g3253 ( 
.A(n_2628),
.B(n_2640),
.Y(n_3253)
);

NOR2xp33_ASAP7_75t_L g3254 ( 
.A(n_2768),
.B(n_2203),
.Y(n_3254)
);

CKINVDCx20_ASAP7_75t_R g3255 ( 
.A(n_2497),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2655),
.B(n_2028),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2689),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2723),
.B(n_2226),
.Y(n_3258)
);

CKINVDCx16_ASAP7_75t_R g3259 ( 
.A(n_2482),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2655),
.B(n_2028),
.Y(n_3260)
);

BUFx3_ASAP7_75t_L g3261 ( 
.A(n_2806),
.Y(n_3261)
);

BUFx6f_ASAP7_75t_L g3262 ( 
.A(n_2762),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2584),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_L g3264 ( 
.A1(n_2786),
.A2(n_1145),
.B1(n_1218),
.B2(n_1140),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_SL g3265 ( 
.A(n_2628),
.B(n_2221),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_2735),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2690),
.Y(n_3267)
);

INVx4_ASAP7_75t_L g3268 ( 
.A(n_2503),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_2640),
.B(n_2384),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_2735),
.B(n_2284),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_2640),
.B(n_2221),
.Y(n_3271)
);

AO22x2_ASAP7_75t_L g3272 ( 
.A1(n_2808),
.A2(n_2413),
.B1(n_2419),
.B2(n_2400),
.Y(n_3272)
);

INVx3_ASAP7_75t_L g3273 ( 
.A(n_2655),
.Y(n_3273)
);

BUFx6f_ASAP7_75t_L g3274 ( 
.A(n_2762),
.Y(n_3274)
);

HB1xp67_ASAP7_75t_L g3275 ( 
.A(n_2747),
.Y(n_3275)
);

BUFx6f_ASAP7_75t_L g3276 ( 
.A(n_2762),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2696),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2584),
.Y(n_3278)
);

INVx5_ASAP7_75t_L g3279 ( 
.A(n_2617),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2682),
.B(n_2028),
.Y(n_3280)
);

INVx2_ASAP7_75t_L g3281 ( 
.A(n_2591),
.Y(n_3281)
);

CKINVDCx5p33_ASAP7_75t_R g3282 ( 
.A(n_2895),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_2901),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_2915),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2917),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_3090),
.B(n_2747),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2864),
.Y(n_3287)
);

AND2x6_ASAP7_75t_SL g3288 ( 
.A(n_3243),
.B(n_2365),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3053),
.B(n_2810),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3053),
.B(n_2564),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_2892),
.B(n_2575),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_2892),
.B(n_2576),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3040),
.A2(n_2649),
.B1(n_2524),
.B2(n_2542),
.Y(n_3293)
);

AND2x4_ASAP7_75t_L g3294 ( 
.A(n_3090),
.B(n_2462),
.Y(n_3294)
);

AOI22xp5_ASAP7_75t_L g3295 ( 
.A1(n_2874),
.A2(n_2649),
.B1(n_2524),
.B2(n_2542),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2942),
.B(n_2634),
.Y(n_3296)
);

BUFx6f_ASAP7_75t_L g3297 ( 
.A(n_3022),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_2896),
.Y(n_3298)
);

NOR2xp33_ASAP7_75t_L g3299 ( 
.A(n_2879),
.B(n_2222),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2942),
.B(n_2645),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_2879),
.B(n_2463),
.Y(n_3301)
);

AO221x1_ASAP7_75t_L g3302 ( 
.A1(n_3001),
.A2(n_2366),
.B1(n_2860),
.B2(n_2809),
.C(n_2853),
.Y(n_3302)
);

BUFx3_ASAP7_75t_L g3303 ( 
.A(n_2914),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3167),
.B(n_2467),
.Y(n_3304)
);

AOI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_2929),
.A2(n_2524),
.B1(n_2542),
.B2(n_2509),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_2980),
.B(n_2468),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2919),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_2980),
.B(n_2469),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2907),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_2910),
.Y(n_3310)
);

INVx2_ASAP7_75t_L g3311 ( 
.A(n_2931),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_2920),
.B(n_3124),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_3048),
.B(n_3124),
.Y(n_3313)
);

INVx2_ASAP7_75t_SL g3314 ( 
.A(n_2865),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_2982),
.B(n_2472),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_2872),
.B(n_2222),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2982),
.B(n_2986),
.Y(n_3317)
);

NAND2xp33_ASAP7_75t_L g3318 ( 
.A(n_3072),
.B(n_2236),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_2937),
.A2(n_2700),
.B(n_2646),
.Y(n_3319)
);

NOR2xp33_ASAP7_75t_L g3320 ( 
.A(n_2872),
.B(n_2946),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2922),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_2986),
.B(n_2976),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_2976),
.B(n_2473),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2930),
.B(n_2236),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2972),
.B(n_2477),
.Y(n_3325)
);

OAI22xp33_ASAP7_75t_L g3326 ( 
.A1(n_2898),
.A2(n_2715),
.B1(n_2650),
.B2(n_2798),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2933),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2972),
.B(n_2478),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3010),
.B(n_2479),
.Y(n_3329)
);

INVx2_ASAP7_75t_SL g3330 ( 
.A(n_2904),
.Y(n_3330)
);

NOR3xp33_ASAP7_75t_L g3331 ( 
.A(n_3254),
.B(n_2379),
.C(n_2367),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_2906),
.Y(n_3332)
);

INVx2_ASAP7_75t_SL g3333 ( 
.A(n_2918),
.Y(n_3333)
);

AOI221xp5_ASAP7_75t_L g3334 ( 
.A1(n_2946),
.A2(n_2458),
.B1(n_2807),
.B2(n_2635),
.C(n_2774),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_3010),
.B(n_2483),
.Y(n_3335)
);

O2A1O1Ixp5_ASAP7_75t_L g3336 ( 
.A1(n_2862),
.A2(n_2538),
.B(n_2646),
.C(n_2596),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_3011),
.B(n_2243),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_3011),
.B(n_2268),
.Y(n_3338)
);

OAI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_2898),
.A2(n_2852),
.B1(n_2711),
.B2(n_2717),
.Y(n_3339)
);

BUFx3_ASAP7_75t_L g3340 ( 
.A(n_2881),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3192),
.B(n_2490),
.Y(n_3341)
);

AOI22xp5_ASAP7_75t_L g3342 ( 
.A1(n_3188),
.A2(n_2648),
.B1(n_2674),
.B2(n_2509),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_2935),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_2955),
.B(n_2400),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_2937),
.B(n_2617),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_3233),
.B(n_2268),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3120),
.B(n_2494),
.Y(n_3347)
);

AO221x1_ASAP7_75t_L g3348 ( 
.A1(n_3001),
.A2(n_2902),
.B1(n_2366),
.B2(n_3272),
.C(n_3051),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3120),
.B(n_2495),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_2945),
.Y(n_3350)
);

AO221x1_ASAP7_75t_L g3351 ( 
.A1(n_2902),
.A2(n_3272),
.B1(n_3051),
.B2(n_2394),
.C(n_2401),
.Y(n_3351)
);

O2A1O1Ixp33_ASAP7_75t_L g3352 ( 
.A1(n_3068),
.A2(n_2823),
.B(n_2835),
.C(n_2843),
.Y(n_3352)
);

OAI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3132),
.A2(n_2821),
.B1(n_2504),
.B2(n_2507),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2924),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3133),
.B(n_2499),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_L g3356 ( 
.A1(n_2887),
.A2(n_2458),
.B1(n_2596),
.B2(n_2648),
.Y(n_3356)
);

OAI22xp5_ASAP7_75t_L g3357 ( 
.A1(n_2888),
.A2(n_2959),
.B1(n_2867),
.B2(n_2900),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_2928),
.Y(n_3358)
);

INVx1_ASAP7_75t_SL g3359 ( 
.A(n_2938),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_2936),
.B(n_2285),
.Y(n_3360)
);

NOR3xp33_ASAP7_75t_L g3361 ( 
.A(n_3254),
.B(n_2390),
.C(n_2389),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_2987),
.B(n_2285),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3028),
.B(n_2513),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_2949),
.Y(n_3364)
);

AOI22xp33_ASAP7_75t_L g3365 ( 
.A1(n_2887),
.A2(n_2648),
.B1(n_2674),
.B2(n_2753),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3028),
.B(n_2521),
.Y(n_3366)
);

O2A1O1Ixp5_ASAP7_75t_L g3367 ( 
.A1(n_2862),
.A2(n_2538),
.B(n_2586),
.C(n_2474),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_SL g3368 ( 
.A(n_3052),
.B(n_2287),
.Y(n_3368)
);

INVx3_ASAP7_75t_L g3369 ( 
.A(n_2923),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_L g3370 ( 
.A(n_3252),
.B(n_2287),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2950),
.B(n_2353),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_SL g3372 ( 
.A(n_3043),
.B(n_2353),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_SL g3373 ( 
.A(n_3253),
.B(n_3091),
.Y(n_3373)
);

NOR2xp33_ASAP7_75t_L g3374 ( 
.A(n_3018),
.B(n_2413),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3031),
.B(n_2531),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3031),
.B(n_3042),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3042),
.B(n_2533),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2913),
.B(n_2535),
.Y(n_3378)
);

O2A1O1Ixp5_ASAP7_75t_L g3379 ( 
.A1(n_2875),
.A2(n_2586),
.B(n_2474),
.C(n_2772),
.Y(n_3379)
);

AOI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_3068),
.A2(n_2674),
.B1(n_2539),
.B2(n_2549),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2941),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_2913),
.B(n_2537),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_2937),
.B(n_2617),
.Y(n_3383)
);

BUFx6f_ASAP7_75t_SL g3384 ( 
.A(n_2908),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_2921),
.B(n_2551),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_SL g3386 ( 
.A(n_2937),
.B(n_2682),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2969),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2921),
.B(n_2555),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_L g3389 ( 
.A(n_2968),
.B(n_2420),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_2970),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_2867),
.A2(n_2505),
.B(n_2503),
.Y(n_3391)
);

AND2x2_ASAP7_75t_SL g3392 ( 
.A(n_2971),
.B(n_2858),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2953),
.Y(n_3393)
);

NOR2xp33_ASAP7_75t_L g3394 ( 
.A(n_2951),
.B(n_3266),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_L g3395 ( 
.A(n_2889),
.B(n_2556),
.Y(n_3395)
);

AOI22xp5_ASAP7_75t_L g3396 ( 
.A1(n_3079),
.A2(n_2559),
.B1(n_2560),
.B2(n_2557),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2889),
.B(n_2569),
.Y(n_3397)
);

OAI221xp5_ASAP7_75t_L g3398 ( 
.A1(n_2932),
.A2(n_3162),
.B1(n_3181),
.B2(n_3132),
.C(n_3266),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_SL g3399 ( 
.A(n_3253),
.B(n_2384),
.Y(n_3399)
);

AOI21xp5_ASAP7_75t_L g3400 ( 
.A1(n_2900),
.A2(n_2506),
.B(n_2505),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3180),
.B(n_2288),
.Y(n_3401)
);

AOI22xp33_ASAP7_75t_L g3402 ( 
.A1(n_2902),
.A2(n_2737),
.B1(n_2789),
.B2(n_2704),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2903),
.B(n_2909),
.Y(n_3403)
);

AOI21xp5_ASAP7_75t_L g3404 ( 
.A1(n_2903),
.A2(n_2506),
.B(n_2505),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2960),
.Y(n_3405)
);

AOI22x1_ASAP7_75t_L g3406 ( 
.A1(n_3232),
.A2(n_2836),
.B1(n_2837),
.B2(n_2830),
.Y(n_3406)
);

NOR2xp33_ASAP7_75t_L g3407 ( 
.A(n_2951),
.B(n_2420),
.Y(n_3407)
);

NAND2xp33_ASAP7_75t_SL g3408 ( 
.A(n_2961),
.B(n_2394),
.Y(n_3408)
);

BUFx12f_ASAP7_75t_L g3409 ( 
.A(n_2871),
.Y(n_3409)
);

INVxp67_ASAP7_75t_L g3410 ( 
.A(n_2926),
.Y(n_3410)
);

AOI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_3079),
.A2(n_2571),
.B1(n_2590),
.B2(n_2587),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_2909),
.B(n_2592),
.Y(n_3412)
);

INVx2_ASAP7_75t_L g3413 ( 
.A(n_3002),
.Y(n_3413)
);

OAI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_2947),
.A2(n_2595),
.B1(n_2601),
.B2(n_2598),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3202),
.B(n_2603),
.Y(n_3415)
);

AOI22xp33_ASAP7_75t_L g3416 ( 
.A1(n_3136),
.A2(n_2737),
.B1(n_2704),
.B2(n_2522),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_3091),
.B(n_2394),
.Y(n_3417)
);

NAND3xp33_ASAP7_75t_L g3418 ( 
.A(n_3102),
.B(n_3023),
.C(n_3066),
.Y(n_3418)
);

INVx2_ASAP7_75t_L g3419 ( 
.A(n_3006),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2963),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3016),
.Y(n_3421)
);

AOI21xp5_ASAP7_75t_L g3422 ( 
.A1(n_3202),
.A2(n_2506),
.B(n_2505),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3086),
.B(n_2605),
.Y(n_3423)
);

INVxp67_ASAP7_75t_L g3424 ( 
.A(n_2926),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_SL g3425 ( 
.A(n_3169),
.B(n_2682),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3025),
.Y(n_3426)
);

AOI21xp5_ASAP7_75t_L g3427 ( 
.A1(n_2959),
.A2(n_2534),
.B(n_2506),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3027),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3036),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_3044),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3275),
.B(n_2422),
.Y(n_3431)
);

AND2x4_ASAP7_75t_L g3432 ( 
.A(n_3156),
.B(n_2607),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_3086),
.B(n_2610),
.Y(n_3433)
);

INVx4_ASAP7_75t_L g3434 ( 
.A(n_2923),
.Y(n_3434)
);

AOI22xp5_ASAP7_75t_L g3435 ( 
.A1(n_3095),
.A2(n_2611),
.B1(n_2619),
.B2(n_2612),
.Y(n_3435)
);

OR2x6_ASAP7_75t_L g3436 ( 
.A(n_2871),
.B(n_2394),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2964),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3095),
.B(n_2620),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_2966),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3098),
.B(n_2621),
.Y(n_3440)
);

NOR2xp67_ASAP7_75t_SL g3441 ( 
.A(n_3169),
.B(n_2534),
.Y(n_3441)
);

INVx1_ASAP7_75t_L g3442 ( 
.A(n_2978),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2988),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_2888),
.A2(n_2540),
.B(n_2534),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_SL g3445 ( 
.A(n_3169),
.B(n_2711),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3275),
.B(n_2422),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3069),
.Y(n_3447)
);

NAND2xp5_ASAP7_75t_L g3448 ( 
.A(n_3098),
.B(n_3106),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3106),
.B(n_2624),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_2998),
.B(n_2629),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3009),
.B(n_2392),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_2990),
.Y(n_3452)
);

AND2x2_ASAP7_75t_L g3453 ( 
.A(n_3270),
.B(n_2303),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3136),
.A2(n_3264),
.B1(n_3143),
.B2(n_2890),
.Y(n_3454)
);

INVxp67_ASAP7_75t_SL g3455 ( 
.A(n_3165),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_3070),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_2998),
.B(n_2633),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_2870),
.B(n_2399),
.Y(n_3458)
);

NAND3xp33_ASAP7_75t_L g3459 ( 
.A(n_3102),
.B(n_2423),
.C(n_2387),
.Y(n_3459)
);

INVx3_ASAP7_75t_L g3460 ( 
.A(n_2923),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3004),
.B(n_2720),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_3156),
.B(n_3161),
.Y(n_3462)
);

AOI22xp33_ASAP7_75t_L g3463 ( 
.A1(n_3143),
.A2(n_2704),
.B1(n_2522),
.B2(n_2702),
.Y(n_3463)
);

NAND2xp33_ASAP7_75t_L g3464 ( 
.A(n_3072),
.B(n_2534),
.Y(n_3464)
);

O2A1O1Ixp5_ASAP7_75t_L g3465 ( 
.A1(n_2875),
.A2(n_2876),
.B(n_2772),
.C(n_3114),
.Y(n_3465)
);

OAI221xp5_ASAP7_75t_L g3466 ( 
.A1(n_3193),
.A2(n_2410),
.B1(n_2418),
.B2(n_2416),
.C(n_2414),
.Y(n_3466)
);

AOI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3004),
.A2(n_3248),
.B1(n_2981),
.B2(n_2983),
.Y(n_3467)
);

OAI22x1_ASAP7_75t_L g3468 ( 
.A1(n_2868),
.A2(n_2387),
.B1(n_2427),
.B2(n_2423),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_SL g3469 ( 
.A(n_3169),
.B(n_2711),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3118),
.B(n_2726),
.Y(n_3470)
);

A2O1A1Ixp33_ASAP7_75t_L g3471 ( 
.A1(n_3007),
.A2(n_2728),
.B(n_2731),
.C(n_2727),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_SL g3472 ( 
.A(n_3161),
.B(n_2401),
.Y(n_3472)
);

INVx2_ASAP7_75t_L g3473 ( 
.A(n_3077),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3118),
.B(n_2733),
.Y(n_3474)
);

NAND2xp5_ASAP7_75t_SL g3475 ( 
.A(n_2965),
.B(n_2401),
.Y(n_3475)
);

OR2x2_ASAP7_75t_L g3476 ( 
.A(n_3019),
.B(n_2424),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3080),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2991),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_L g3479 ( 
.A(n_3030),
.B(n_2738),
.Y(n_3479)
);

OR2x2_ASAP7_75t_L g3480 ( 
.A(n_3087),
.B(n_2426),
.Y(n_3480)
);

NAND2xp33_ASAP7_75t_L g3481 ( 
.A(n_3072),
.B(n_2540),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3030),
.B(n_2739),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_2992),
.Y(n_3483)
);

AND2x6_ASAP7_75t_SL g3484 ( 
.A(n_3243),
.B(n_2432),
.Y(n_3484)
);

OAI22x1_ASAP7_75t_R g3485 ( 
.A1(n_3123),
.A2(n_2312),
.B1(n_2391),
.B2(n_2293),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3032),
.B(n_3220),
.Y(n_3486)
);

INVx2_ASAP7_75t_SL g3487 ( 
.A(n_3029),
.Y(n_3487)
);

INVx2_ASAP7_75t_L g3488 ( 
.A(n_3084),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_SL g3489 ( 
.A(n_3248),
.B(n_2401),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3222),
.B(n_2098),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3264),
.A2(n_2704),
.B1(n_2706),
.B2(n_2697),
.Y(n_3491)
);

BUFx3_ASAP7_75t_L g3492 ( 
.A(n_3020),
.Y(n_3492)
);

INVx2_ASAP7_75t_SL g3493 ( 
.A(n_2958),
.Y(n_3493)
);

NOR2xp33_ASAP7_75t_L g3494 ( 
.A(n_3066),
.B(n_2436),
.Y(n_3494)
);

INVx2_ASAP7_75t_SL g3495 ( 
.A(n_2974),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_3039),
.B(n_2540),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3032),
.B(n_2741),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2996),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3003),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3220),
.B(n_2743),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_2981),
.B(n_2744),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3085),
.Y(n_3502)
);

INVx2_ASAP7_75t_L g3503 ( 
.A(n_3093),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3039),
.B(n_2540),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_SL g3505 ( 
.A(n_3269),
.B(n_2585),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_2983),
.B(n_2745),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_SL g3507 ( 
.A(n_3269),
.B(n_2585),
.Y(n_3507)
);

INVx2_ASAP7_75t_L g3508 ( 
.A(n_3103),
.Y(n_3508)
);

INVx2_ASAP7_75t_SL g3509 ( 
.A(n_3144),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3114),
.B(n_2746),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3116),
.B(n_3154),
.Y(n_3511)
);

INVx2_ASAP7_75t_SL g3512 ( 
.A(n_3246),
.Y(n_3512)
);

NOR2xp33_ASAP7_75t_L g3513 ( 
.A(n_3128),
.B(n_2748),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_3116),
.B(n_2717),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3012),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3015),
.Y(n_3516)
);

NOR2xp33_ASAP7_75t_L g3517 ( 
.A(n_3128),
.B(n_2179),
.Y(n_3517)
);

OAI22xp5_ASAP7_75t_L g3518 ( 
.A1(n_2962),
.A2(n_2717),
.B1(n_2844),
.B2(n_2838),
.Y(n_3518)
);

AOI21xp5_ASAP7_75t_L g3519 ( 
.A1(n_3097),
.A2(n_2600),
.B(n_2585),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_3258),
.B(n_2098),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3017),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3154),
.B(n_2671),
.Y(n_3522)
);

OAI22xp5_ASAP7_75t_L g3523 ( 
.A1(n_2962),
.A2(n_2585),
.B1(n_2647),
.B2(n_2600),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3021),
.Y(n_3524)
);

AND2x4_ASAP7_75t_L g3525 ( 
.A(n_2882),
.B(n_3216),
.Y(n_3525)
);

OR2x2_ASAP7_75t_L g3526 ( 
.A(n_3210),
.B(n_2405),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_2861),
.B(n_2866),
.Y(n_3527)
);

O2A1O1Ixp33_ASAP7_75t_L g3528 ( 
.A1(n_3234),
.A2(n_2823),
.B(n_2698),
.C(n_2678),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_2873),
.B(n_2729),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3139),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_2877),
.B(n_2732),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3026),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3163),
.Y(n_3533)
);

INVx2_ASAP7_75t_L g3534 ( 
.A(n_3184),
.Y(n_3534)
);

NAND2xp33_ASAP7_75t_L g3535 ( 
.A(n_3072),
.B(n_3074),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_2878),
.B(n_2785),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_2971),
.B(n_3187),
.Y(n_3537)
);

INVx2_ASAP7_75t_SL g3538 ( 
.A(n_3050),
.Y(n_3538)
);

NAND3xp33_ASAP7_75t_L g3539 ( 
.A(n_3193),
.B(n_2434),
.C(n_2427),
.Y(n_3539)
);

AOI221xp5_ASAP7_75t_L g3540 ( 
.A1(n_3214),
.A2(n_2526),
.B1(n_855),
.B2(n_856),
.C(n_853),
.Y(n_3540)
);

AO21x2_ASAP7_75t_L g3541 ( 
.A1(n_2876),
.A2(n_2849),
.B(n_2488),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_2883),
.B(n_2707),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_SL g3543 ( 
.A(n_3065),
.B(n_2179),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3199),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_2891),
.B(n_2709),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3218),
.Y(n_3546)
);

INVx2_ASAP7_75t_L g3547 ( 
.A(n_3224),
.Y(n_3547)
);

INVx8_ASAP7_75t_L g3548 ( 
.A(n_2906),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_2893),
.B(n_2710),
.Y(n_3549)
);

AND2x2_ASAP7_75t_L g3550 ( 
.A(n_3214),
.B(n_2098),
.Y(n_3550)
);

AOI22xp33_ASAP7_75t_L g3551 ( 
.A1(n_2890),
.A2(n_2704),
.B1(n_2713),
.B2(n_2693),
.Y(n_3551)
);

A2O1A1Ixp33_ASAP7_75t_L g3552 ( 
.A1(n_3140),
.A2(n_2820),
.B(n_2819),
.C(n_2824),
.Y(n_3552)
);

INVx2_ASAP7_75t_L g3553 ( 
.A(n_3250),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_L g3554 ( 
.A(n_3179),
.B(n_3034),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_2863),
.B(n_2553),
.Y(n_3555)
);

INVx2_ASAP7_75t_L g3556 ( 
.A(n_3251),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_2863),
.B(n_2553),
.Y(n_3557)
);

NOR2xp33_ASAP7_75t_L g3558 ( 
.A(n_3179),
.B(n_2430),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3263),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_SL g3560 ( 
.A(n_3173),
.B(n_2600),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_SL g3561 ( 
.A(n_3173),
.B(n_2600),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3033),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_SL g3563 ( 
.A(n_2911),
.B(n_2304),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_2884),
.B(n_2553),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_2884),
.B(n_2558),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3047),
.Y(n_3566)
);

BUFx3_ASAP7_75t_L g3567 ( 
.A(n_3073),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3140),
.B(n_2558),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3141),
.B(n_2558),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_L g3570 ( 
.A(n_3034),
.B(n_3117),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3141),
.B(n_2566),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3278),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3147),
.B(n_2566),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3281),
.Y(n_3574)
);

AOI22xp33_ASAP7_75t_L g3575 ( 
.A1(n_2894),
.A2(n_2704),
.B1(n_2693),
.B2(n_1218),
.Y(n_3575)
);

AND2x2_ASAP7_75t_L g3576 ( 
.A(n_3117),
.B(n_2362),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_L g3577 ( 
.A(n_3160),
.B(n_2381),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3187),
.B(n_3147),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_L g3579 ( 
.A(n_3160),
.B(n_2403),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_3207),
.B(n_2403),
.Y(n_3580)
);

INVxp67_ASAP7_75t_L g3581 ( 
.A(n_3207),
.Y(n_3581)
);

AOI22xp33_ASAP7_75t_L g3582 ( 
.A1(n_2894),
.A2(n_1218),
.B1(n_1145),
.B2(n_1058),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3054),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3175),
.B(n_2566),
.Y(n_3584)
);

NAND2xp5_ASAP7_75t_L g3585 ( 
.A(n_3175),
.B(n_2825),
.Y(n_3585)
);

OAI22xp5_ASAP7_75t_L g3586 ( 
.A1(n_3173),
.A2(n_3279),
.B1(n_3125),
.B2(n_3208),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_3177),
.A2(n_2386),
.B1(n_2335),
.B2(n_2347),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3067),
.Y(n_3588)
);

OAI22xp33_ASAP7_75t_L g3589 ( 
.A1(n_3243),
.A2(n_2386),
.B1(n_1145),
.B2(n_2434),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3177),
.B(n_2647),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3035),
.B(n_2304),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_L g3592 ( 
.A(n_2993),
.B(n_3064),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_2940),
.B(n_3211),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3078),
.Y(n_3594)
);

INVx4_ASAP7_75t_L g3595 ( 
.A(n_2925),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3083),
.B(n_2335),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3212),
.B(n_2647),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3088),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_L g3599 ( 
.A(n_3225),
.B(n_2647),
.Y(n_3599)
);

NOR2xp33_ASAP7_75t_L g3600 ( 
.A(n_3137),
.B(n_2347),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3096),
.Y(n_3601)
);

NAND2xp5_ASAP7_75t_SL g3602 ( 
.A(n_3216),
.B(n_2662),
.Y(n_3602)
);

INVxp33_ASAP7_75t_L g3603 ( 
.A(n_3111),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_SL g3604 ( 
.A(n_3121),
.B(n_2662),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3099),
.Y(n_3605)
);

OR2x6_ASAP7_75t_L g3606 ( 
.A(n_2871),
.B(n_2070),
.Y(n_3606)
);

INVx2_ASAP7_75t_SL g3607 ( 
.A(n_2916),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3227),
.B(n_2662),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3228),
.B(n_2662),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3230),
.B(n_2666),
.Y(n_3610)
);

NOR2xp67_ASAP7_75t_L g3611 ( 
.A(n_3058),
.B(n_2178),
.Y(n_3611)
);

AND2x4_ASAP7_75t_L g3612 ( 
.A(n_2882),
.B(n_2804),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3231),
.B(n_3236),
.Y(n_3613)
);

AOI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_2989),
.A2(n_2849),
.B1(n_2180),
.B2(n_2178),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3241),
.B(n_2666),
.Y(n_3615)
);

NAND2xp5_ASAP7_75t_L g3616 ( 
.A(n_3244),
.B(n_2666),
.Y(n_3616)
);

NAND2xp5_ASAP7_75t_SL g3617 ( 
.A(n_3121),
.B(n_2666),
.Y(n_3617)
);

NOR2xp33_ASAP7_75t_L g3618 ( 
.A(n_3209),
.B(n_2180),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3100),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3257),
.B(n_2692),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3267),
.B(n_2692),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_SL g3622 ( 
.A(n_3127),
.B(n_2692),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3277),
.B(n_2692),
.Y(n_3623)
);

OR2x2_ASAP7_75t_L g3624 ( 
.A(n_2957),
.B(n_2407),
.Y(n_3624)
);

AOI221xp5_ASAP7_75t_SL g3625 ( 
.A1(n_3234),
.A2(n_1062),
.B1(n_1073),
.B2(n_1063),
.C(n_1053),
.Y(n_3625)
);

INVx3_ASAP7_75t_L g3626 ( 
.A(n_2925),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_L g3627 ( 
.A(n_2957),
.B(n_2096),
.Y(n_3627)
);

BUFx2_ASAP7_75t_L g3628 ( 
.A(n_2906),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3101),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3237),
.Y(n_3630)
);

AND2x4_ASAP7_75t_L g3631 ( 
.A(n_3261),
.B(n_2804),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3247),
.Y(n_3632)
);

INVx2_ASAP7_75t_SL g3633 ( 
.A(n_3149),
.Y(n_3633)
);

INVxp67_ASAP7_75t_L g3634 ( 
.A(n_3191),
.Y(n_3634)
);

BUFx2_ASAP7_75t_R g3635 ( 
.A(n_2948),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3097),
.A2(n_2460),
.B(n_2841),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_3127),
.B(n_2171),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3041),
.B(n_2593),
.Y(n_3638)
);

BUFx3_ASAP7_75t_L g3639 ( 
.A(n_3217),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_3148),
.B(n_2593),
.Y(n_3640)
);

CKINVDCx5p33_ASAP7_75t_R g3641 ( 
.A(n_2997),
.Y(n_3641)
);

NOR2xp33_ASAP7_75t_L g3642 ( 
.A(n_2984),
.B(n_2108),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3148),
.B(n_2615),
.Y(n_3643)
);

AND2x4_ASAP7_75t_L g3644 ( 
.A(n_2939),
.B(n_2812),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3153),
.B(n_2615),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3153),
.B(n_2851),
.Y(n_3646)
);

NOR2xp33_ASAP7_75t_L g3647 ( 
.A(n_3240),
.B(n_2145),
.Y(n_3647)
);

OR2x2_ASAP7_75t_L g3648 ( 
.A(n_3071),
.B(n_2030),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_3197),
.B(n_2859),
.Y(n_3649)
);

A2O1A1Ixp33_ASAP7_75t_L g3650 ( 
.A1(n_3126),
.A2(n_2591),
.B(n_2818),
.C(n_2812),
.Y(n_3650)
);

AOI22xp5_ASAP7_75t_L g3651 ( 
.A1(n_2994),
.A2(n_2391),
.B1(n_2415),
.B2(n_2312),
.Y(n_3651)
);

AO22x1_ASAP7_75t_L g3652 ( 
.A1(n_3146),
.A2(n_2072),
.B1(n_2077),
.B2(n_2030),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3249),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_L g3654 ( 
.A(n_3240),
.B(n_2072),
.Y(n_3654)
);

INVx2_ASAP7_75t_L g3655 ( 
.A(n_3107),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3197),
.B(n_2826),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3109),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3110),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3203),
.B(n_2826),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3203),
.B(n_2851),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_L g3661 ( 
.A(n_3229),
.B(n_2077),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3131),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3205),
.B(n_2818),
.Y(n_3663)
);

INVx3_ASAP7_75t_L g3664 ( 
.A(n_3612),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3283),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3284),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3605),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3376),
.B(n_2995),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3290),
.B(n_2999),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3655),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3658),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3322),
.B(n_3142),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3403),
.A2(n_3279),
.B(n_3173),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_SL g3674 ( 
.A(n_3372),
.B(n_3182),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3285),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_R g3676 ( 
.A(n_3282),
.B(n_2415),
.Y(n_3676)
);

AO22x1_ASAP7_75t_L g3677 ( 
.A1(n_3316),
.A2(n_3517),
.B1(n_3299),
.B2(n_3370),
.Y(n_3677)
);

BUFx2_ASAP7_75t_L g3678 ( 
.A(n_3303),
.Y(n_3678)
);

INVxp67_ASAP7_75t_L g3679 ( 
.A(n_3389),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3320),
.B(n_3005),
.Y(n_3680)
);

INVx5_ASAP7_75t_L g3681 ( 
.A(n_3297),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3287),
.Y(n_3682)
);

BUFx4f_ASAP7_75t_L g3683 ( 
.A(n_3409),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3302),
.A2(n_3182),
.B1(n_3196),
.B2(n_3189),
.Y(n_3684)
);

BUFx6f_ASAP7_75t_L g3685 ( 
.A(n_3297),
.Y(n_3685)
);

AOI22xp5_ASAP7_75t_L g3686 ( 
.A1(n_3299),
.A2(n_3265),
.B1(n_3271),
.B2(n_3242),
.Y(n_3686)
);

INVx4_ASAP7_75t_L g3687 ( 
.A(n_3548),
.Y(n_3687)
);

INVx1_ASAP7_75t_L g3688 ( 
.A(n_3307),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3317),
.B(n_3142),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3401),
.B(n_2943),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3320),
.B(n_3115),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3298),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_3347),
.B(n_3130),
.Y(n_3693)
);

INVx3_ASAP7_75t_L g3694 ( 
.A(n_3612),
.Y(n_3694)
);

NAND2x1p5_ASAP7_75t_L g3695 ( 
.A(n_3441),
.B(n_2869),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3309),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3321),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_SL g3698 ( 
.A(n_3418),
.B(n_3189),
.Y(n_3698)
);

INVxp67_ASAP7_75t_L g3699 ( 
.A(n_3389),
.Y(n_3699)
);

AND2x4_ASAP7_75t_L g3700 ( 
.A(n_3525),
.B(n_2899),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_L g3701 ( 
.A(n_3349),
.B(n_3134),
.Y(n_3701)
);

OAI22xp5_ASAP7_75t_SL g3702 ( 
.A1(n_3494),
.A2(n_3151),
.B1(n_3255),
.B2(n_3259),
.Y(n_3702)
);

INVx2_ASAP7_75t_L g3703 ( 
.A(n_3310),
.Y(n_3703)
);

BUFx6f_ASAP7_75t_L g3704 ( 
.A(n_3297),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3311),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3327),
.Y(n_3706)
);

CKINVDCx5p33_ASAP7_75t_R g3707 ( 
.A(n_3641),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3343),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3350),
.Y(n_3709)
);

BUFx2_ASAP7_75t_SL g3710 ( 
.A(n_3333),
.Y(n_3710)
);

OR2x6_ASAP7_75t_L g3711 ( 
.A(n_3548),
.B(n_2943),
.Y(n_3711)
);

NOR2xp33_ASAP7_75t_L g3712 ( 
.A(n_3316),
.B(n_2083),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3354),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3358),
.Y(n_3714)
);

OAI221xp5_ASAP7_75t_L g3715 ( 
.A1(n_3334),
.A2(n_2979),
.B1(n_2095),
.B2(n_2113),
.C(n_2089),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3364),
.Y(n_3716)
);

AO21x2_ASAP7_75t_L g3717 ( 
.A1(n_3312),
.A2(n_3082),
.B(n_3075),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3387),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3390),
.Y(n_3719)
);

AOI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3589),
.A2(n_3196),
.B1(n_3094),
.B2(n_2943),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3296),
.B(n_3150),
.Y(n_3721)
);

BUFx6f_ASAP7_75t_L g3722 ( 
.A(n_3297),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3527),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3346),
.B(n_3081),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3300),
.B(n_3172),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3413),
.Y(n_3726)
);

INVx1_ASAP7_75t_L g3727 ( 
.A(n_3613),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3419),
.Y(n_3728)
);

NAND2xp5_ASAP7_75t_SL g3729 ( 
.A(n_3346),
.B(n_3105),
.Y(n_3729)
);

INVxp67_ASAP7_75t_L g3730 ( 
.A(n_3592),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_SL g3731 ( 
.A(n_3370),
.B(n_3105),
.Y(n_3731)
);

HB1xp67_ASAP7_75t_L g3732 ( 
.A(n_3359),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3363),
.B(n_2885),
.Y(n_3733)
);

INVx3_ASAP7_75t_SL g3734 ( 
.A(n_3436),
.Y(n_3734)
);

INVx1_ASAP7_75t_L g3735 ( 
.A(n_3381),
.Y(n_3735)
);

NAND2x1p5_ASAP7_75t_L g3736 ( 
.A(n_3639),
.B(n_2869),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3291),
.B(n_3142),
.Y(n_3737)
);

INVx3_ASAP7_75t_L g3738 ( 
.A(n_3644),
.Y(n_3738)
);

NAND2x1p5_ASAP7_75t_L g3739 ( 
.A(n_3487),
.B(n_2905),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3393),
.Y(n_3740)
);

OAI22xp5_ASAP7_75t_SL g3741 ( 
.A1(n_3494),
.A2(n_3158),
.B1(n_3159),
.B2(n_2089),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3405),
.Y(n_3742)
);

INVx2_ASAP7_75t_SL g3743 ( 
.A(n_3493),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3420),
.Y(n_3744)
);

O2A1O1Ixp5_ASAP7_75t_L g3745 ( 
.A1(n_3312),
.A2(n_2927),
.B(n_2954),
.C(n_2944),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_L g3746 ( 
.A(n_3517),
.B(n_2083),
.Y(n_3746)
);

INVx3_ASAP7_75t_L g3747 ( 
.A(n_3644),
.Y(n_3747)
);

AOI22xp5_ASAP7_75t_L g3748 ( 
.A1(n_3313),
.A2(n_3094),
.B1(n_3062),
.B2(n_3201),
.Y(n_3748)
);

CKINVDCx5p33_ASAP7_75t_R g3749 ( 
.A(n_3635),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3437),
.Y(n_3750)
);

INVx1_ASAP7_75t_L g3751 ( 
.A(n_3439),
.Y(n_3751)
);

INVx2_ASAP7_75t_SL g3752 ( 
.A(n_3567),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3366),
.B(n_2885),
.Y(n_3753)
);

AOI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3513),
.A2(n_2975),
.B1(n_3272),
.B2(n_3051),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3442),
.Y(n_3755)
);

INVxp67_ASAP7_75t_L g3756 ( 
.A(n_3592),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3443),
.Y(n_3757)
);

INVx2_ASAP7_75t_L g3758 ( 
.A(n_3421),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3292),
.B(n_3142),
.Y(n_3759)
);

NAND2xp5_ASAP7_75t_L g3760 ( 
.A(n_3375),
.B(n_2886),
.Y(n_3760)
);

AND2x6_ASAP7_75t_L g3761 ( 
.A(n_3305),
.B(n_2952),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_3306),
.B(n_3142),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_3344),
.B(n_3526),
.Y(n_3763)
);

INVx3_ASAP7_75t_L g3764 ( 
.A(n_3434),
.Y(n_3764)
);

BUFx4f_ASAP7_75t_L g3765 ( 
.A(n_3436),
.Y(n_3765)
);

AOI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3513),
.A2(n_2939),
.B1(n_3221),
.B2(n_2886),
.Y(n_3766)
);

NAND2xp5_ASAP7_75t_L g3767 ( 
.A(n_3377),
.B(n_2912),
.Y(n_3767)
);

AND2x4_ASAP7_75t_L g3768 ( 
.A(n_3525),
.B(n_2899),
.Y(n_3768)
);

A2O1A1Ixp33_ASAP7_75t_SL g3769 ( 
.A1(n_3558),
.A2(n_2880),
.B(n_3125),
.C(n_3205),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3323),
.B(n_2912),
.Y(n_3770)
);

CKINVDCx5p33_ASAP7_75t_R g3771 ( 
.A(n_3492),
.Y(n_3771)
);

INVx5_ASAP7_75t_L g3772 ( 
.A(n_3548),
.Y(n_3772)
);

NOR3xp33_ASAP7_75t_SL g3773 ( 
.A(n_3589),
.B(n_2113),
.C(n_2095),
.Y(n_3773)
);

INVx3_ASAP7_75t_L g3774 ( 
.A(n_3434),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3308),
.B(n_3245),
.Y(n_3775)
);

OR2x2_ASAP7_75t_SL g3776 ( 
.A(n_3648),
.B(n_2899),
.Y(n_3776)
);

INVxp67_ASAP7_75t_L g3777 ( 
.A(n_3624),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3464),
.A2(n_3279),
.B(n_3063),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3452),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_SL g3780 ( 
.A(n_3587),
.B(n_2925),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3478),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3426),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3483),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_3325),
.B(n_3221),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3558),
.B(n_2137),
.Y(n_3785)
);

AOI22xp33_ASAP7_75t_SL g3786 ( 
.A1(n_3661),
.A2(n_2137),
.B1(n_2934),
.B2(n_2066),
.Y(n_3786)
);

INVx3_ASAP7_75t_L g3787 ( 
.A(n_3595),
.Y(n_3787)
);

INVx2_ASAP7_75t_L g3788 ( 
.A(n_3428),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3498),
.Y(n_3789)
);

INVx3_ASAP7_75t_L g3790 ( 
.A(n_3595),
.Y(n_3790)
);

AND2x2_ASAP7_75t_SL g3791 ( 
.A(n_3318),
.B(n_3239),
.Y(n_3791)
);

BUFx2_ASAP7_75t_L g3792 ( 
.A(n_3591),
.Y(n_3792)
);

NAND2xp5_ASAP7_75t_L g3793 ( 
.A(n_3328),
.B(n_3245),
.Y(n_3793)
);

AND2x4_ASAP7_75t_L g3794 ( 
.A(n_3286),
.B(n_3512),
.Y(n_3794)
);

NOR2xp33_ASAP7_75t_L g3795 ( 
.A(n_3337),
.B(n_3108),
.Y(n_3795)
);

CKINVDCx5p33_ASAP7_75t_R g3796 ( 
.A(n_3340),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_SL g3797 ( 
.A(n_3337),
.B(n_3038),
.Y(n_3797)
);

INVx4_ASAP7_75t_L g3798 ( 
.A(n_3436),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_3338),
.B(n_3038),
.Y(n_3799)
);

INVx2_ASAP7_75t_L g3800 ( 
.A(n_3429),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3499),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3515),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3516),
.Y(n_3803)
);

BUFx3_ASAP7_75t_L g3804 ( 
.A(n_3314),
.Y(n_3804)
);

AOI22xp5_ASAP7_75t_L g3805 ( 
.A1(n_3654),
.A2(n_3219),
.B1(n_3113),
.B2(n_3138),
.Y(n_3805)
);

INVx4_ASAP7_75t_L g3806 ( 
.A(n_3369),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3521),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3329),
.B(n_3273),
.Y(n_3808)
);

INVx2_ASAP7_75t_SL g3809 ( 
.A(n_3330),
.Y(n_3809)
);

BUFx6f_ASAP7_75t_L g3810 ( 
.A(n_3332),
.Y(n_3810)
);

BUFx6f_ASAP7_75t_L g3811 ( 
.A(n_3628),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3335),
.B(n_3273),
.Y(n_3812)
);

AND2x4_ASAP7_75t_L g3813 ( 
.A(n_3286),
.B(n_3215),
.Y(n_3813)
);

BUFx8_ASAP7_75t_L g3814 ( 
.A(n_3384),
.Y(n_3814)
);

BUFx6f_ASAP7_75t_L g3815 ( 
.A(n_3607),
.Y(n_3815)
);

INVx2_ASAP7_75t_SL g3816 ( 
.A(n_3633),
.Y(n_3816)
);

AND2x4_ASAP7_75t_L g3817 ( 
.A(n_3432),
.B(n_3215),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3430),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3423),
.B(n_3208),
.Y(n_3819)
);

OAI22xp5_ASAP7_75t_SL g3820 ( 
.A1(n_3466),
.A2(n_2967),
.B1(n_2219),
.B2(n_857),
.Y(n_3820)
);

AND2x2_ASAP7_75t_L g3821 ( 
.A(n_3453),
.B(n_3550),
.Y(n_3821)
);

HB1xp67_ASAP7_75t_L g3822 ( 
.A(n_3410),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3524),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3433),
.B(n_2905),
.Y(n_3824)
);

AND2x4_ASAP7_75t_L g3825 ( 
.A(n_3432),
.B(n_3215),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3447),
.Y(n_3826)
);

BUFx6f_ASAP7_75t_L g3827 ( 
.A(n_3369),
.Y(n_3827)
);

OAI22xp5_ASAP7_75t_SL g3828 ( 
.A1(n_3654),
.A2(n_2967),
.B1(n_860),
.B2(n_861),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3438),
.B(n_2952),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_3301),
.B(n_3315),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3394),
.B(n_2956),
.Y(n_3831)
);

NAND2xp5_ASAP7_75t_SL g3832 ( 
.A(n_3338),
.B(n_3279),
.Y(n_3832)
);

OR2x6_ASAP7_75t_L g3833 ( 
.A(n_3606),
.B(n_3204),
.Y(n_3833)
);

BUFx12f_ASAP7_75t_L g3834 ( 
.A(n_3606),
.Y(n_3834)
);

BUFx6f_ASAP7_75t_L g3835 ( 
.A(n_3460),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_SL g3836 ( 
.A(n_3371),
.B(n_2066),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3532),
.Y(n_3837)
);

AND2x4_ASAP7_75t_L g3838 ( 
.A(n_3294),
.B(n_3462),
.Y(n_3838)
);

NOR2xp33_ASAP7_75t_L g3839 ( 
.A(n_3554),
.B(n_3108),
.Y(n_3839)
);

AO22x1_ASAP7_75t_L g3840 ( 
.A1(n_3371),
.A2(n_2066),
.B1(n_3074),
.B2(n_3072),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_3394),
.B(n_2956),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3562),
.Y(n_3842)
);

NAND2x1p5_ASAP7_75t_L g3843 ( 
.A(n_3509),
.B(n_3024),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3566),
.Y(n_3844)
);

BUFx3_ASAP7_75t_L g3845 ( 
.A(n_3538),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3410),
.Y(n_3846)
);

CKINVDCx20_ASAP7_75t_R g3847 ( 
.A(n_3485),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_SL g3848 ( 
.A(n_3467),
.B(n_3611),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3456),
.Y(n_3849)
);

INVx2_ASAP7_75t_SL g3850 ( 
.A(n_3476),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3583),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3588),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3594),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3596),
.B(n_2171),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_3554),
.B(n_2148),
.Y(n_3855)
);

INVx2_ASAP7_75t_L g3856 ( 
.A(n_3473),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_SL g3857 ( 
.A(n_3596),
.B(n_3600),
.Y(n_3857)
);

BUFx2_ASAP7_75t_L g3858 ( 
.A(n_3634),
.Y(n_3858)
);

NAND2x1p5_ASAP7_75t_L g3859 ( 
.A(n_3460),
.B(n_3000),
.Y(n_3859)
);

AOI22xp33_ASAP7_75t_L g3860 ( 
.A1(n_3331),
.A2(n_3113),
.B1(n_3219),
.B2(n_3145),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_SL g3861 ( 
.A(n_3600),
.B(n_3262),
.Y(n_3861)
);

INVxp67_ASAP7_75t_L g3862 ( 
.A(n_3374),
.Y(n_3862)
);

OAI22xp5_ASAP7_75t_SL g3863 ( 
.A1(n_3661),
.A2(n_864),
.B1(n_866),
.B2(n_851),
.Y(n_3863)
);

HB1xp67_ASAP7_75t_L g3864 ( 
.A(n_3424),
.Y(n_3864)
);

NOR2xp33_ASAP7_75t_SL g3865 ( 
.A(n_3543),
.B(n_3074),
.Y(n_3865)
);

BUFx2_ASAP7_75t_L g3866 ( 
.A(n_3634),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3598),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3601),
.Y(n_3868)
);

OR2x2_ASAP7_75t_L g3869 ( 
.A(n_3480),
.B(n_3135),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3618),
.B(n_3276),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3618),
.B(n_3276),
.Y(n_3871)
);

OAI22xp5_ASAP7_75t_SL g3872 ( 
.A1(n_3539),
.A2(n_868),
.B1(n_870),
.B2(n_867),
.Y(n_3872)
);

HB1xp67_ASAP7_75t_L g3873 ( 
.A(n_3424),
.Y(n_3873)
);

NOR2xp33_ASAP7_75t_L g3874 ( 
.A(n_3450),
.B(n_3152),
.Y(n_3874)
);

INVx2_ASAP7_75t_SL g3875 ( 
.A(n_3606),
.Y(n_3875)
);

INVxp67_ASAP7_75t_L g3876 ( 
.A(n_3374),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3619),
.Y(n_3877)
);

INVx3_ASAP7_75t_L g3878 ( 
.A(n_3626),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_SL g3879 ( 
.A(n_3458),
.B(n_3226),
.Y(n_3879)
);

BUFx2_ASAP7_75t_L g3880 ( 
.A(n_3581),
.Y(n_3880)
);

AOI22xp33_ASAP7_75t_L g3881 ( 
.A1(n_3331),
.A2(n_3219),
.B1(n_3157),
.B2(n_3166),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3576),
.B(n_3164),
.Y(n_3882)
);

INVx2_ASAP7_75t_L g3883 ( 
.A(n_3477),
.Y(n_3883)
);

AND2x6_ASAP7_75t_SL g3884 ( 
.A(n_3642),
.B(n_1062),
.Y(n_3884)
);

NOR2xp33_ASAP7_75t_L g3885 ( 
.A(n_3457),
.B(n_3168),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3488),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_3626),
.Y(n_3887)
);

INVxp67_ASAP7_75t_SL g3888 ( 
.A(n_3455),
.Y(n_3888)
);

AO22x1_ASAP7_75t_L g3889 ( 
.A1(n_3642),
.A2(n_3176),
.B1(n_3074),
.B2(n_3008),
.Y(n_3889)
);

BUFx12f_ASAP7_75t_L g3890 ( 
.A(n_3484),
.Y(n_3890)
);

INVxp67_ASAP7_75t_L g3891 ( 
.A(n_3627),
.Y(n_3891)
);

AOI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3407),
.A2(n_3219),
.B1(n_3171),
.B2(n_3195),
.Y(n_3892)
);

INVx2_ASAP7_75t_L g3893 ( 
.A(n_3502),
.Y(n_3893)
);

AND2x4_ASAP7_75t_L g3894 ( 
.A(n_3294),
.B(n_3186),
.Y(n_3894)
);

AOI22xp33_ASAP7_75t_L g3895 ( 
.A1(n_3361),
.A2(n_3219),
.B1(n_3198),
.B2(n_3176),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3629),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_3461),
.B(n_2973),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3407),
.B(n_2973),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3657),
.Y(n_3899)
);

NAND2xp5_ASAP7_75t_L g3900 ( 
.A(n_3289),
.B(n_2977),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3662),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3490),
.B(n_1542),
.Y(n_3902)
);

AND2x4_ASAP7_75t_L g3903 ( 
.A(n_3373),
.B(n_2977),
.Y(n_3903)
);

INVxp67_ASAP7_75t_L g3904 ( 
.A(n_3627),
.Y(n_3904)
);

AOI22xp33_ASAP7_75t_L g3905 ( 
.A1(n_3361),
.A2(n_3176),
.B1(n_3074),
.B2(n_2985),
.Y(n_3905)
);

INVx3_ASAP7_75t_L g3906 ( 
.A(n_3631),
.Y(n_3906)
);

AOI22xp5_ASAP7_75t_L g3907 ( 
.A1(n_3647),
.A2(n_3176),
.B1(n_2985),
.B2(n_3092),
.Y(n_3907)
);

AOI22x1_ASAP7_75t_L g3908 ( 
.A1(n_3455),
.A2(n_3092),
.B1(n_3119),
.B2(n_3013),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3503),
.Y(n_3909)
);

AND2x6_ASAP7_75t_SL g3910 ( 
.A(n_3458),
.B(n_1063),
.Y(n_3910)
);

BUFx12f_ASAP7_75t_L g3911 ( 
.A(n_3495),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3508),
.Y(n_3912)
);

INVx2_ASAP7_75t_L g3913 ( 
.A(n_3530),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_SL g3914 ( 
.A(n_3647),
.B(n_3226),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3533),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3534),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3614),
.B(n_3451),
.Y(n_3917)
);

INVx3_ASAP7_75t_L g3918 ( 
.A(n_3631),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3544),
.Y(n_3919)
);

OAI22xp5_ASAP7_75t_L g3920 ( 
.A1(n_3454),
.A2(n_3055),
.B1(n_3063),
.B2(n_3013),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3378),
.B(n_3119),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3546),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3547),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3593),
.Y(n_3924)
);

BUFx2_ASAP7_75t_L g3925 ( 
.A(n_3581),
.Y(n_3925)
);

BUFx3_ASAP7_75t_L g3926 ( 
.A(n_3570),
.Y(n_3926)
);

AOI22x1_ASAP7_75t_L g3927 ( 
.A1(n_3444),
.A2(n_2839),
.B1(n_2840),
.B2(n_2822),
.Y(n_3927)
);

AOI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3392),
.A2(n_3176),
.B1(n_3008),
.B2(n_3014),
.Y(n_3928)
);

BUFx6f_ASAP7_75t_SL g3929 ( 
.A(n_3392),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3382),
.B(n_3055),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3542),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3385),
.B(n_2897),
.Y(n_3932)
);

BUFx6f_ASAP7_75t_L g3933 ( 
.A(n_3417),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_SL g3934 ( 
.A(n_3451),
.B(n_3262),
.Y(n_3934)
);

INVxp67_ASAP7_75t_L g3935 ( 
.A(n_3570),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3545),
.Y(n_3936)
);

CKINVDCx5p33_ASAP7_75t_R g3937 ( 
.A(n_3384),
.Y(n_3937)
);

INVx2_ASAP7_75t_L g3938 ( 
.A(n_3553),
.Y(n_3938)
);

AND2x4_ASAP7_75t_L g3939 ( 
.A(n_3399),
.B(n_3000),
.Y(n_3939)
);

CKINVDCx5p33_ASAP7_75t_R g3940 ( 
.A(n_3288),
.Y(n_3940)
);

AOI22xp5_ASAP7_75t_L g3941 ( 
.A1(n_3431),
.A2(n_3008),
.B1(n_3014),
.B2(n_2897),
.Y(n_3941)
);

INVx2_ASAP7_75t_SL g3942 ( 
.A(n_3520),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_SL g3943 ( 
.A(n_3651),
.B(n_3262),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3549),
.Y(n_3944)
);

AND2x4_ASAP7_75t_L g3945 ( 
.A(n_3489),
.B(n_3024),
.Y(n_3945)
);

NAND2xp33_ASAP7_75t_SL g3946 ( 
.A(n_3928),
.B(n_3454),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_SL g3947 ( 
.A(n_3686),
.B(n_3459),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_SL g3948 ( 
.A(n_3686),
.B(n_3355),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3857),
.B(n_3324),
.Y(n_3949)
);

NAND2xp33_ASAP7_75t_SL g3950 ( 
.A(n_3929),
.B(n_3365),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3712),
.B(n_3360),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_SL g3952 ( 
.A(n_3785),
.B(n_3362),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3830),
.B(n_3388),
.Y(n_3953)
);

NAND2xp33_ASAP7_75t_SL g3954 ( 
.A(n_3929),
.B(n_3365),
.Y(n_3954)
);

NOR2xp33_ASAP7_75t_L g3955 ( 
.A(n_3677),
.B(n_3603),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_SL g3956 ( 
.A(n_3746),
.B(n_3396),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_SL g3957 ( 
.A(n_3784),
.B(n_3411),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_SL g3958 ( 
.A(n_3679),
.B(n_3435),
.Y(n_3958)
);

AND2x4_ASAP7_75t_L g3959 ( 
.A(n_3772),
.B(n_3537),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_L g3960 ( 
.A(n_3924),
.B(n_3304),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3723),
.B(n_3501),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3699),
.B(n_3506),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3862),
.B(n_3500),
.Y(n_3963)
);

NAND2xp33_ASAP7_75t_SL g3964 ( 
.A(n_3702),
.B(n_3468),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3876),
.B(n_3368),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_SL g3966 ( 
.A(n_3766),
.B(n_3470),
.Y(n_3966)
);

NAND2xp33_ASAP7_75t_SL g3967 ( 
.A(n_3702),
.B(n_3637),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3766),
.B(n_3474),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3917),
.B(n_3380),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_SL g3970 ( 
.A(n_3891),
.B(n_3577),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3904),
.B(n_3727),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_SL g3972 ( 
.A(n_3850),
.B(n_3931),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_SL g3973 ( 
.A(n_3936),
.B(n_3577),
.Y(n_3973)
);

NAND2xp33_ASAP7_75t_SL g3974 ( 
.A(n_3676),
.B(n_3341),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3944),
.B(n_3579),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3680),
.B(n_3579),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3691),
.B(n_3580),
.Y(n_3977)
);

NAND2xp33_ASAP7_75t_SL g3978 ( 
.A(n_3741),
.B(n_3578),
.Y(n_3978)
);

NAND2xp33_ASAP7_75t_SL g3979 ( 
.A(n_3741),
.B(n_3395),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_3821),
.B(n_3431),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_SL g3981 ( 
.A(n_3733),
.B(n_3580),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3753),
.B(n_3414),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_3760),
.B(n_3414),
.Y(n_3983)
);

NAND2xp33_ASAP7_75t_SL g3984 ( 
.A(n_3707),
.B(n_3397),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_SL g3985 ( 
.A(n_3767),
.B(n_3730),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_SL g3986 ( 
.A(n_3756),
.B(n_3353),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_L g3987 ( 
.A(n_3763),
.B(n_3446),
.Y(n_3987)
);

NAND2xp5_ASAP7_75t_L g3988 ( 
.A(n_3874),
.B(n_3446),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_SL g3989 ( 
.A(n_3854),
.B(n_3353),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_SL g3990 ( 
.A(n_3865),
.B(n_3293),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3865),
.B(n_3295),
.Y(n_3991)
);

NAND2xp33_ASAP7_75t_SL g3992 ( 
.A(n_3773),
.B(n_3412),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3770),
.B(n_3563),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3855),
.B(n_3529),
.Y(n_3994)
);

NAND2xp33_ASAP7_75t_SL g3995 ( 
.A(n_3847),
.B(n_3415),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_SL g3996 ( 
.A(n_3669),
.B(n_3531),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3885),
.B(n_3536),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_SL g3998 ( 
.A(n_3926),
.B(n_3510),
.Y(n_3998)
);

NAND2xp33_ASAP7_75t_SL g3999 ( 
.A(n_3749),
.B(n_3472),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3839),
.B(n_3342),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3721),
.B(n_3479),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_SL g4002 ( 
.A(n_3725),
.B(n_3482),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3848),
.B(n_3497),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_SL g4004 ( 
.A(n_3935),
.B(n_3724),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3668),
.B(n_3638),
.Y(n_4005)
);

NAND2xp33_ASAP7_75t_SL g4006 ( 
.A(n_3734),
.B(n_3356),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3882),
.B(n_3522),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3693),
.B(n_3356),
.Y(n_4008)
);

NAND2xp33_ASAP7_75t_SL g4009 ( 
.A(n_3820),
.B(n_3491),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_SL g4010 ( 
.A(n_3701),
.B(n_3440),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_SL g4011 ( 
.A(n_3838),
.B(n_3449),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_SL g4012 ( 
.A(n_3838),
.B(n_3408),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_SL g4013 ( 
.A(n_3795),
.B(n_3475),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_SL g4014 ( 
.A(n_3869),
.B(n_3486),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3792),
.B(n_3585),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_3894),
.B(n_3590),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3894),
.B(n_3540),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3674),
.B(n_3471),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_SL g4019 ( 
.A(n_3765),
.B(n_3698),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_SL g4020 ( 
.A(n_3765),
.B(n_3786),
.Y(n_4020)
);

NAND2xp33_ASAP7_75t_SL g4021 ( 
.A(n_3820),
.B(n_3491),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3777),
.B(n_3326),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_SL g4023 ( 
.A(n_3748),
.B(n_3326),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3902),
.B(n_3398),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3748),
.B(n_3528),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3729),
.B(n_3352),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_SL g4027 ( 
.A(n_3731),
.B(n_3511),
.Y(n_4027)
);

NAND2xp5_ASAP7_75t_L g4028 ( 
.A(n_3690),
.B(n_3652),
.Y(n_4028)
);

NAND2xp33_ASAP7_75t_SL g4029 ( 
.A(n_3687),
.B(n_3463),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_SL g4030 ( 
.A(n_3738),
.B(n_3597),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_SL g4031 ( 
.A(n_3738),
.B(n_3747),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_SL g4032 ( 
.A(n_3747),
.B(n_3599),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_SL g4033 ( 
.A(n_3772),
.B(n_3608),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_SL g4034 ( 
.A(n_3772),
.B(n_3609),
.Y(n_4034)
);

NAND2xp5_ASAP7_75t_SL g4035 ( 
.A(n_3933),
.B(n_3610),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3930),
.B(n_3653),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3933),
.B(n_3615),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_SL g4038 ( 
.A(n_3933),
.B(n_3903),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3903),
.B(n_3664),
.Y(n_4039)
);

NAND2xp33_ASAP7_75t_SL g4040 ( 
.A(n_3687),
.B(n_3463),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3732),
.B(n_3630),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_3664),
.B(n_3616),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_SL g4043 ( 
.A(n_3694),
.B(n_3620),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3694),
.B(n_3621),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_SL g4045 ( 
.A(n_3861),
.B(n_3870),
.Y(n_4045)
);

NAND2xp5_ASAP7_75t_SL g4046 ( 
.A(n_3871),
.B(n_3623),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3831),
.B(n_3632),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_SL g4048 ( 
.A(n_3940),
.B(n_3906),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_3906),
.B(n_3357),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3841),
.B(n_3625),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_SL g4051 ( 
.A(n_3918),
.B(n_3568),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_3819),
.B(n_3556),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_SL g4053 ( 
.A(n_3918),
.B(n_3569),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3794),
.B(n_3559),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_3794),
.B(n_3572),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3797),
.B(n_3571),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_SL g4057 ( 
.A(n_3799),
.B(n_3573),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_SL g4058 ( 
.A(n_3942),
.B(n_3584),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_3720),
.B(n_3574),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_3828),
.B(n_3496),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_SL g4061 ( 
.A(n_3828),
.B(n_3504),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_3914),
.B(n_3586),
.Y(n_4062)
);

NAND2xp33_ASAP7_75t_SL g4063 ( 
.A(n_3905),
.B(n_3345),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_SL g4064 ( 
.A(n_3810),
.B(n_3514),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_SL g4065 ( 
.A(n_3810),
.B(n_3602),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3822),
.B(n_3448),
.Y(n_4066)
);

NAND2xp33_ASAP7_75t_SL g4067 ( 
.A(n_3798),
.B(n_3345),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3810),
.B(n_3604),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_SL g4069 ( 
.A(n_3811),
.B(n_3617),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_SL g4070 ( 
.A(n_3811),
.B(n_3622),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3811),
.B(n_3402),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_SL g4072 ( 
.A(n_3824),
.B(n_3402),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_SL g4073 ( 
.A(n_3684),
.B(n_3523),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_SL g4074 ( 
.A(n_3880),
.B(n_3319),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_3925),
.B(n_3391),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_3872),
.B(n_3400),
.Y(n_4076)
);

NAND2xp33_ASAP7_75t_SL g4077 ( 
.A(n_3798),
.B(n_3383),
.Y(n_4077)
);

AND2x4_ASAP7_75t_L g4078 ( 
.A(n_3711),
.B(n_3505),
.Y(n_4078)
);

NAND2xp33_ASAP7_75t_SL g4079 ( 
.A(n_3817),
.B(n_3383),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3872),
.B(n_3404),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3683),
.B(n_3422),
.Y(n_4081)
);

NAND2xp33_ASAP7_75t_SL g4082 ( 
.A(n_3815),
.B(n_3022),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3683),
.B(n_3339),
.Y(n_4083)
);

NAND2xp33_ASAP7_75t_SL g4084 ( 
.A(n_3815),
.B(n_3022),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_SL g4085 ( 
.A(n_3771),
.B(n_3640),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3667),
.B(n_3643),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3846),
.B(n_3348),
.Y(n_4087)
);

NAND2xp33_ASAP7_75t_SL g4088 ( 
.A(n_3815),
.B(n_3045),
.Y(n_4088)
);

NAND2xp5_ASAP7_75t_SL g4089 ( 
.A(n_3670),
.B(n_3645),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_SL g4090 ( 
.A(n_3671),
.B(n_3507),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3864),
.B(n_3582),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_3879),
.B(n_3552),
.Y(n_4092)
);

NAND2xp33_ASAP7_75t_SL g4093 ( 
.A(n_3752),
.B(n_3045),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_SL g4094 ( 
.A(n_3875),
.B(n_3037),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_SL g4095 ( 
.A(n_3873),
.B(n_3037),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_SL g4096 ( 
.A(n_3836),
.B(n_3057),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_SL g4097 ( 
.A(n_3796),
.B(n_3881),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3907),
.B(n_3057),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_3700),
.B(n_3768),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_3907),
.B(n_3122),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_3775),
.B(n_3582),
.Y(n_4101)
);

NAND2xp33_ASAP7_75t_SL g4102 ( 
.A(n_3743),
.B(n_3045),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_SL g4103 ( 
.A(n_3858),
.B(n_3122),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_SL g4104 ( 
.A(n_3866),
.B(n_3155),
.Y(n_4104)
);

NAND2xp33_ASAP7_75t_SL g4105 ( 
.A(n_3809),
.B(n_3046),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_SL g4106 ( 
.A(n_3888),
.B(n_3155),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3775),
.B(n_3351),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_3943),
.B(n_3170),
.Y(n_4108)
);

NAND2xp5_ASAP7_75t_SL g4109 ( 
.A(n_3678),
.B(n_3170),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_SL g4110 ( 
.A(n_3805),
.B(n_3174),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3805),
.B(n_3174),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_3934),
.B(n_3178),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_SL g4113 ( 
.A(n_3898),
.B(n_3178),
.Y(n_4113)
);

NAND2xp33_ASAP7_75t_SL g4114 ( 
.A(n_3816),
.B(n_3046),
.Y(n_4114)
);

NAND2xp33_ASAP7_75t_SL g4115 ( 
.A(n_3937),
.B(n_3046),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_SL g4116 ( 
.A(n_3793),
.B(n_3185),
.Y(n_4116)
);

XNOR2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3863),
.B(n_6),
.Y(n_4117)
);

NAND2xp33_ASAP7_75t_SL g4118 ( 
.A(n_3817),
.B(n_3049),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_3808),
.B(n_3185),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3812),
.B(n_3200),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_SL g4121 ( 
.A(n_3932),
.B(n_3200),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_SL g4122 ( 
.A(n_3863),
.B(n_3223),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_SL g4123 ( 
.A(n_3897),
.B(n_3223),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_3700),
.B(n_1544),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_SL g4125 ( 
.A(n_3912),
.B(n_3238),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_SL g4126 ( 
.A(n_3916),
.B(n_3238),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_SL g4127 ( 
.A(n_3919),
.B(n_3268),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_3829),
.B(n_3555),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_SL g4129 ( 
.A(n_3923),
.B(n_3268),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_3768),
.B(n_3921),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_SL g4131 ( 
.A(n_3939),
.B(n_3427),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_SL g4132 ( 
.A(n_3939),
.B(n_3659),
.Y(n_4132)
);

NAND2xp33_ASAP7_75t_SL g4133 ( 
.A(n_3825),
.B(n_3049),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3945),
.B(n_3660),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_3945),
.B(n_3663),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3739),
.B(n_3646),
.Y(n_4136)
);

NAND2xp33_ASAP7_75t_SL g4137 ( 
.A(n_3825),
.B(n_3049),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_SL g4138 ( 
.A(n_3941),
.B(n_3762),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3665),
.B(n_3557),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_SL g4140 ( 
.A(n_3941),
.B(n_3649),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_SL g4141 ( 
.A(n_3762),
.B(n_3656),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_SL g4142 ( 
.A(n_3737),
.B(n_3204),
.Y(n_4142)
);

NAND2xp33_ASAP7_75t_L g4143 ( 
.A(n_3761),
.B(n_3008),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_SL g4144 ( 
.A(n_3737),
.B(n_3204),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_SL g4145 ( 
.A(n_3759),
.B(n_3206),
.Y(n_4145)
);

AND2x4_ASAP7_75t_L g4146 ( 
.A(n_3711),
.B(n_3650),
.Y(n_4146)
);

AND2x2_ASAP7_75t_L g4147 ( 
.A(n_3682),
.B(n_1547),
.Y(n_4147)
);

NAND2xp33_ASAP7_75t_SL g4148 ( 
.A(n_3813),
.B(n_3056),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_SL g4149 ( 
.A(n_3759),
.B(n_3226),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_SL g4150 ( 
.A(n_3895),
.B(n_3235),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_3692),
.B(n_1548),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_SL g4152 ( 
.A(n_3780),
.B(n_3206),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_SL g4153 ( 
.A(n_3696),
.B(n_3206),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3666),
.B(n_3564),
.Y(n_4154)
);

NAND2xp5_ASAP7_75t_SL g4155 ( 
.A(n_3703),
.B(n_3274),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_SL g4156 ( 
.A(n_3705),
.B(n_3274),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_SL g4157 ( 
.A(n_3706),
.B(n_3274),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_3708),
.B(n_3709),
.Y(n_4158)
);

NAND2xp5_ASAP7_75t_SL g4159 ( 
.A(n_3716),
.B(n_3718),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_SL g4160 ( 
.A(n_3719),
.B(n_3276),
.Y(n_4160)
);

NAND2xp33_ASAP7_75t_SL g4161 ( 
.A(n_3813),
.B(n_3056),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_SL g4162 ( 
.A(n_3726),
.B(n_3235),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_SL g4163 ( 
.A(n_3728),
.B(n_3235),
.Y(n_4163)
);

NAND2xp33_ASAP7_75t_SL g4164 ( 
.A(n_3675),
.B(n_3056),
.Y(n_4164)
);

NAND2xp5_ASAP7_75t_SL g4165 ( 
.A(n_3758),
.B(n_3061),
.Y(n_4165)
);

AND2x4_ASAP7_75t_L g4166 ( 
.A(n_3711),
.B(n_3386),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_SL g4167 ( 
.A(n_3782),
.B(n_3061),
.Y(n_4167)
);

NAND2xp5_ASAP7_75t_L g4168 ( 
.A(n_3688),
.B(n_3565),
.Y(n_4168)
);

NAND2xp5_ASAP7_75t_L g4169 ( 
.A(n_3697),
.B(n_2897),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_SL g4170 ( 
.A(n_3788),
.B(n_3061),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_3713),
.B(n_2897),
.Y(n_4171)
);

XNOR2xp5_ASAP7_75t_L g4172 ( 
.A(n_3776),
.B(n_3575),
.Y(n_4172)
);

NAND2xp33_ASAP7_75t_SL g4173 ( 
.A(n_3714),
.B(n_3076),
.Y(n_4173)
);

NAND2xp33_ASAP7_75t_SL g4174 ( 
.A(n_3827),
.B(n_3076),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_SL g4175 ( 
.A(n_3800),
.B(n_3076),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3910),
.B(n_2897),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_SL g4177 ( 
.A(n_3818),
.B(n_3104),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_SL g4178 ( 
.A(n_3826),
.B(n_3104),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_SL g4179 ( 
.A(n_3849),
.B(n_3104),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3910),
.B(n_3008),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_SL g4181 ( 
.A(n_3856),
.B(n_3183),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_SL g4182 ( 
.A(n_3883),
.B(n_3183),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_SL g4183 ( 
.A(n_3886),
.B(n_3183),
.Y(n_4183)
);

NAND2xp33_ASAP7_75t_SL g4184 ( 
.A(n_3827),
.B(n_3190),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_SL g4185 ( 
.A(n_3893),
.B(n_3190),
.Y(n_4185)
);

NAND2xp33_ASAP7_75t_SL g4186 ( 
.A(n_3827),
.B(n_3190),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_L g4187 ( 
.A(n_3710),
.B(n_3014),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3909),
.B(n_3014),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_SL g4189 ( 
.A(n_3913),
.B(n_3519),
.Y(n_4189)
);

NAND2xp5_ASAP7_75t_SL g4190 ( 
.A(n_3915),
.B(n_3336),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_3922),
.B(n_3336),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_SL g4192 ( 
.A(n_3938),
.B(n_3416),
.Y(n_4192)
);

NAND2xp33_ASAP7_75t_SL g4193 ( 
.A(n_3920),
.B(n_3416),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_3845),
.B(n_3059),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_SL g4195 ( 
.A(n_3892),
.B(n_3059),
.Y(n_4195)
);

NAND2xp5_ASAP7_75t_L g4196 ( 
.A(n_3735),
.B(n_3014),
.Y(n_4196)
);

NAND2xp33_ASAP7_75t_SL g4197 ( 
.A(n_3920),
.B(n_3560),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_3740),
.B(n_3060),
.Y(n_4198)
);

NAND2xp33_ASAP7_75t_SL g4199 ( 
.A(n_3672),
.B(n_3560),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_SL g4200 ( 
.A(n_3892),
.B(n_3129),
.Y(n_4200)
);

AND2x4_ASAP7_75t_L g4201 ( 
.A(n_3833),
.B(n_3386),
.Y(n_4201)
);

NAND2xp5_ASAP7_75t_SL g4202 ( 
.A(n_3742),
.B(n_3129),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_SL g4203 ( 
.A(n_3744),
.B(n_3750),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3751),
.B(n_3060),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_SL g4205 ( 
.A(n_3755),
.B(n_3194),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_4158),
.Y(n_4206)
);

NAND2xp5_ASAP7_75t_L g4207 ( 
.A(n_3988),
.B(n_3757),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4203),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_3994),
.B(n_3715),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_4159),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_SL g4211 ( 
.A(n_3984),
.B(n_3860),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4054),
.Y(n_4212)
);

AND2x4_ASAP7_75t_L g4213 ( 
.A(n_4201),
.B(n_3833),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_4066),
.Y(n_4214)
);

INVx3_ASAP7_75t_L g4215 ( 
.A(n_3959),
.Y(n_4215)
);

INVx4_ASAP7_75t_L g4216 ( 
.A(n_4124),
.Y(n_4216)
);

INVx5_ASAP7_75t_L g4217 ( 
.A(n_3959),
.Y(n_4217)
);

INVx2_ASAP7_75t_L g4218 ( 
.A(n_4055),
.Y(n_4218)
);

OAI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_3997),
.A2(n_3833),
.B1(n_3890),
.B2(n_3754),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4007),
.B(n_3779),
.Y(n_4220)
);

BUFx2_ASAP7_75t_L g4221 ( 
.A(n_4099),
.Y(n_4221)
);

BUFx8_ASAP7_75t_L g4222 ( 
.A(n_4147),
.Y(n_4222)
);

INVx2_ASAP7_75t_L g4223 ( 
.A(n_4151),
.Y(n_4223)
);

O2A1O1Ixp33_ASAP7_75t_SL g4224 ( 
.A1(n_3956),
.A2(n_3769),
.B(n_3832),
.C(n_3672),
.Y(n_4224)
);

OAI22xp5_ASAP7_75t_L g4225 ( 
.A1(n_4172),
.A2(n_3754),
.B1(n_3843),
.B2(n_3834),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_3972),
.Y(n_4226)
);

INVx2_ASAP7_75t_SL g4227 ( 
.A(n_4041),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_3953),
.B(n_3781),
.Y(n_4228)
);

BUFx6f_ASAP7_75t_L g4229 ( 
.A(n_4201),
.Y(n_4229)
);

AND2x4_ASAP7_75t_L g4230 ( 
.A(n_4201),
.B(n_4078),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3961),
.B(n_3783),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_3987),
.B(n_3789),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_4090),
.Y(n_4233)
);

NOR2xp33_ASAP7_75t_L g4234 ( 
.A(n_4000),
.B(n_3884),
.Y(n_4234)
);

AOI21xp5_ASAP7_75t_L g4235 ( 
.A1(n_4143),
.A2(n_3481),
.B(n_3535),
.Y(n_4235)
);

INVx2_ASAP7_75t_L g4236 ( 
.A(n_4130),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_3980),
.B(n_3998),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_3960),
.Y(n_4238)
);

INVx3_ASAP7_75t_L g4239 ( 
.A(n_3959),
.Y(n_4239)
);

AND2x2_ASAP7_75t_L g4240 ( 
.A(n_3985),
.B(n_3867),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3996),
.B(n_3801),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_4023),
.A2(n_3673),
.B(n_3778),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4014),
.B(n_3802),
.Y(n_4243)
);

BUFx6f_ASAP7_75t_L g4244 ( 
.A(n_4078),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_SL g4245 ( 
.A(n_4024),
.B(n_3791),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4022),
.B(n_3803),
.Y(n_4246)
);

INVx2_ASAP7_75t_L g4247 ( 
.A(n_4086),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_SL g4248 ( 
.A(n_3995),
.B(n_3745),
.Y(n_4248)
);

INVxp67_ASAP7_75t_SL g4249 ( 
.A(n_4015),
.Y(n_4249)
);

INVx3_ASAP7_75t_L g4250 ( 
.A(n_4078),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_3976),
.B(n_3807),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_L g4252 ( 
.A(n_3977),
.B(n_3823),
.Y(n_4252)
);

INVx6_ASAP7_75t_L g4253 ( 
.A(n_4166),
.Y(n_4253)
);

INVxp67_ASAP7_75t_SL g4254 ( 
.A(n_4139),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_3971),
.Y(n_4255)
);

BUFx2_ASAP7_75t_L g4256 ( 
.A(n_4028),
.Y(n_4256)
);

CKINVDCx5p33_ASAP7_75t_R g4257 ( 
.A(n_4004),
.Y(n_4257)
);

BUFx2_ASAP7_75t_L g4258 ( 
.A(n_4082),
.Y(n_4258)
);

BUFx4f_ASAP7_75t_L g4259 ( 
.A(n_4166),
.Y(n_4259)
);

BUFx2_ASAP7_75t_L g4260 ( 
.A(n_4084),
.Y(n_4260)
);

BUFx2_ASAP7_75t_L g4261 ( 
.A(n_4088),
.Y(n_4261)
);

CKINVDCx11_ASAP7_75t_R g4262 ( 
.A(n_4166),
.Y(n_4262)
);

NAND2x1p5_ASAP7_75t_L g4263 ( 
.A(n_4033),
.B(n_3681),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4087),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_4089),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_4193),
.A2(n_3889),
.B(n_3840),
.Y(n_4266)
);

INVx4_ASAP7_75t_L g4267 ( 
.A(n_4146),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_3979),
.B(n_3837),
.Y(n_4268)
);

BUFx6f_ASAP7_75t_L g4269 ( 
.A(n_4038),
.Y(n_4269)
);

NAND2xp5_ASAP7_75t_SL g4270 ( 
.A(n_3955),
.B(n_3842),
.Y(n_4270)
);

AND2x4_ASAP7_75t_SL g4271 ( 
.A(n_4146),
.B(n_3764),
.Y(n_4271)
);

BUFx2_ASAP7_75t_L g4272 ( 
.A(n_4093),
.Y(n_4272)
);

BUFx6f_ASAP7_75t_L g4273 ( 
.A(n_4048),
.Y(n_4273)
);

INVx1_ASAP7_75t_L g4274 ( 
.A(n_4154),
.Y(n_4274)
);

INVx8_ASAP7_75t_L g4275 ( 
.A(n_4146),
.Y(n_4275)
);

CKINVDCx20_ASAP7_75t_R g4276 ( 
.A(n_3974),
.Y(n_4276)
);

AOI21xp5_ASAP7_75t_L g4277 ( 
.A1(n_4193),
.A2(n_3689),
.B(n_3900),
.Y(n_4277)
);

CKINVDCx5p33_ASAP7_75t_R g4278 ( 
.A(n_3964),
.Y(n_4278)
);

BUFx6f_ASAP7_75t_L g4279 ( 
.A(n_4194),
.Y(n_4279)
);

NOR2xp33_ASAP7_75t_L g4280 ( 
.A(n_3951),
.B(n_3884),
.Y(n_4280)
);

BUFx2_ASAP7_75t_L g4281 ( 
.A(n_4102),
.Y(n_4281)
);

OAI22xp5_ASAP7_75t_L g4282 ( 
.A1(n_4176),
.A2(n_3736),
.B1(n_3851),
.B2(n_3844),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_3965),
.B(n_3868),
.Y(n_4283)
);

HB1xp67_ASAP7_75t_L g4284 ( 
.A(n_4064),
.Y(n_4284)
);

OAI22xp5_ASAP7_75t_L g4285 ( 
.A1(n_4180),
.A2(n_3852),
.B1(n_3877),
.B2(n_3853),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_4168),
.Y(n_4286)
);

BUFx12f_ASAP7_75t_L g4287 ( 
.A(n_4117),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3963),
.B(n_3896),
.Y(n_4288)
);

OAI22xp5_ASAP7_75t_L g4289 ( 
.A1(n_4097),
.A2(n_3952),
.B1(n_4017),
.B2(n_4060),
.Y(n_4289)
);

O2A1O1Ixp33_ASAP7_75t_L g4290 ( 
.A1(n_3947),
.A2(n_3989),
.B(n_3969),
.C(n_4061),
.Y(n_4290)
);

INVx2_ASAP7_75t_L g4291 ( 
.A(n_4058),
.Y(n_4291)
);

A2O1A1Ixp33_ASAP7_75t_L g4292 ( 
.A1(n_3978),
.A2(n_3901),
.B(n_3899),
.C(n_3239),
.Y(n_4292)
);

OAI22xp33_ASAP7_75t_L g4293 ( 
.A1(n_4020),
.A2(n_3804),
.B1(n_3689),
.B2(n_3900),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_3958),
.B(n_3761),
.Y(n_4294)
);

AND2x2_ASAP7_75t_L g4295 ( 
.A(n_3970),
.B(n_3878),
.Y(n_4295)
);

INVxp67_ASAP7_75t_L g4296 ( 
.A(n_3949),
.Y(n_4296)
);

AOI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_4025),
.A2(n_3908),
.B(n_3636),
.Y(n_4297)
);

AO22x1_ASAP7_75t_L g4298 ( 
.A1(n_4050),
.A2(n_3761),
.B1(n_3814),
.B2(n_4187),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4047),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4153),
.Y(n_4300)
);

BUFx3_ASAP7_75t_L g4301 ( 
.A(n_4169),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_SL g4302 ( 
.A(n_3993),
.B(n_3835),
.Y(n_4302)
);

NOR2xp33_ASAP7_75t_L g4303 ( 
.A(n_4085),
.B(n_3911),
.Y(n_4303)
);

OAI22xp5_ASAP7_75t_L g4304 ( 
.A1(n_4019),
.A2(n_3695),
.B1(n_3774),
.B2(n_3764),
.Y(n_4304)
);

NOR2x1_ASAP7_75t_L g4305 ( 
.A(n_3962),
.B(n_3806),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4155),
.Y(n_4306)
);

BUFx6f_ASAP7_75t_L g4307 ( 
.A(n_4109),
.Y(n_4307)
);

BUFx6f_ASAP7_75t_L g4308 ( 
.A(n_4103),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4156),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_4001),
.B(n_4002),
.Y(n_4310)
);

INVx4_ASAP7_75t_L g4311 ( 
.A(n_4105),
.Y(n_4311)
);

AOI21xp5_ASAP7_75t_L g4312 ( 
.A1(n_4003),
.A2(n_3561),
.B(n_3445),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_4107),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_3986),
.B(n_4010),
.Y(n_4314)
);

O2A1O1Ixp33_ASAP7_75t_L g4315 ( 
.A1(n_4013),
.A2(n_1074),
.B(n_1075),
.C(n_1073),
.Y(n_4315)
);

OR2x6_ASAP7_75t_L g4316 ( 
.A(n_4012),
.B(n_3859),
.Y(n_4316)
);

INVxp67_ASAP7_75t_SL g4317 ( 
.A(n_4011),
.Y(n_4317)
);

AOI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_3967),
.A2(n_3761),
.B1(n_3814),
.B2(n_875),
.Y(n_4318)
);

INVx2_ASAP7_75t_L g4319 ( 
.A(n_4157),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4160),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_4190),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_3948),
.A2(n_3561),
.B(n_3445),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4191),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4016),
.B(n_3878),
.Y(n_4324)
);

A2O1A1Ixp33_ASAP7_75t_L g4325 ( 
.A1(n_4009),
.A2(n_3194),
.B(n_3367),
.C(n_3465),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_3981),
.B(n_3887),
.Y(n_4326)
);

INVx2_ASAP7_75t_L g4327 ( 
.A(n_4162),
.Y(n_4327)
);

OAI22xp5_ASAP7_75t_L g4328 ( 
.A1(n_3973),
.A2(n_3787),
.B1(n_3790),
.B2(n_3774),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_4045),
.Y(n_4329)
);

O2A1O1Ixp33_ASAP7_75t_L g4330 ( 
.A1(n_4026),
.A2(n_4076),
.B(n_4080),
.C(n_3957),
.Y(n_4330)
);

BUFx8_ASAP7_75t_L g4331 ( 
.A(n_4115),
.Y(n_4331)
);

AOI22xp33_ASAP7_75t_L g4332 ( 
.A1(n_4021),
.A2(n_1042),
.B1(n_1056),
.B2(n_1000),
.Y(n_4332)
);

AOI21x1_ASAP7_75t_L g4333 ( 
.A1(n_4018),
.A2(n_3518),
.B(n_3469),
.Y(n_4333)
);

OR2x6_ASAP7_75t_L g4334 ( 
.A(n_3990),
.B(n_3787),
.Y(n_4334)
);

NAND2xp5_ASAP7_75t_SL g4335 ( 
.A(n_4027),
.B(n_3835),
.Y(n_4335)
);

BUFx3_ASAP7_75t_L g4336 ( 
.A(n_4171),
.Y(n_4336)
);

AOI221xp5_ASAP7_75t_SL g4337 ( 
.A1(n_4083),
.A2(n_1075),
.B1(n_1078),
.B2(n_1077),
.C(n_1074),
.Y(n_4337)
);

OAI21xp5_ASAP7_75t_L g4338 ( 
.A1(n_3982),
.A2(n_3367),
.B(n_3379),
.Y(n_4338)
);

AND2x2_ASAP7_75t_L g4339 ( 
.A(n_3975),
.B(n_3887),
.Y(n_4339)
);

NAND2xp5_ASAP7_75t_L g4340 ( 
.A(n_4005),
.B(n_3835),
.Y(n_4340)
);

INVx2_ASAP7_75t_L g4341 ( 
.A(n_4163),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4036),
.B(n_3717),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4052),
.B(n_3966),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_4142),
.Y(n_4344)
);

AOI22xp33_ASAP7_75t_L g4345 ( 
.A1(n_4021),
.A2(n_1056),
.B1(n_1103),
.B2(n_1042),
.Y(n_4345)
);

NOR2xp33_ASAP7_75t_L g4346 ( 
.A(n_4096),
.B(n_3806),
.Y(n_4346)
);

AOI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_4110),
.A2(n_4111),
.B(n_3968),
.Y(n_4347)
);

INVx2_ASAP7_75t_L g4348 ( 
.A(n_4165),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4144),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4145),
.Y(n_4350)
);

O2A1O1Ixp33_ASAP7_75t_L g4351 ( 
.A1(n_4073),
.A2(n_1078),
.B(n_1081),
.C(n_1077),
.Y(n_4351)
);

INVx2_ASAP7_75t_SL g4352 ( 
.A(n_4104),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4149),
.Y(n_4353)
);

BUFx2_ASAP7_75t_L g4354 ( 
.A(n_4114),
.Y(n_4354)
);

INVx2_ASAP7_75t_L g4355 ( 
.A(n_4167),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4074),
.Y(n_4356)
);

O2A1O1Ixp33_ASAP7_75t_L g4357 ( 
.A1(n_3983),
.A2(n_1082),
.B(n_1091),
.C(n_1081),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_4141),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4152),
.Y(n_4359)
);

A2O1A1Ixp33_ASAP7_75t_SL g4360 ( 
.A1(n_4196),
.A2(n_3790),
.B(n_3575),
.C(n_1551),
.Y(n_4360)
);

AND2x4_ASAP7_75t_L g4361 ( 
.A(n_4039),
.B(n_3681),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4138),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_4031),
.B(n_3681),
.Y(n_4363)
);

NOR2xp33_ASAP7_75t_L g4364 ( 
.A(n_3999),
.B(n_3685),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_SL g4365 ( 
.A(n_3992),
.B(n_3685),
.Y(n_4365)
);

AND2x4_ASAP7_75t_L g4366 ( 
.A(n_4202),
.B(n_3685),
.Y(n_4366)
);

BUFx12f_ASAP7_75t_L g4367 ( 
.A(n_4081),
.Y(n_4367)
);

INVx5_ASAP7_75t_L g4368 ( 
.A(n_4164),
.Y(n_4368)
);

BUFx2_ASAP7_75t_L g4369 ( 
.A(n_4006),
.Y(n_4369)
);

BUFx8_ASAP7_75t_L g4370 ( 
.A(n_4118),
.Y(n_4370)
);

AOI22xp33_ASAP7_75t_L g4371 ( 
.A1(n_3950),
.A2(n_1056),
.B1(n_1103),
.B2(n_1042),
.Y(n_4371)
);

AOI22xp5_ASAP7_75t_L g4372 ( 
.A1(n_3950),
.A2(n_877),
.B1(n_882),
.B2(n_873),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4051),
.Y(n_4373)
);

INVx5_ASAP7_75t_L g4374 ( 
.A(n_4173),
.Y(n_4374)
);

BUFx2_ASAP7_75t_L g4375 ( 
.A(n_4174),
.Y(n_4375)
);

INVx2_ASAP7_75t_L g4376 ( 
.A(n_4170),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4175),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4053),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4071),
.Y(n_4379)
);

OAI22xp5_ASAP7_75t_L g4380 ( 
.A1(n_4122),
.A2(n_3551),
.B1(n_3425),
.B2(n_3469),
.Y(n_4380)
);

AOI22xp5_ASAP7_75t_L g4381 ( 
.A1(n_3954),
.A2(n_885),
.B1(n_887),
.B2(n_883),
.Y(n_4381)
);

INVx2_ASAP7_75t_L g4382 ( 
.A(n_4177),
.Y(n_4382)
);

AND2x6_ASAP7_75t_L g4383 ( 
.A(n_4198),
.B(n_3704),
.Y(n_4383)
);

BUFx3_ASAP7_75t_L g4384 ( 
.A(n_4204),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4178),
.Y(n_4385)
);

OR2x6_ASAP7_75t_L g4386 ( 
.A(n_3991),
.B(n_3704),
.Y(n_4386)
);

O2A1O1Ixp33_ASAP7_75t_L g4387 ( 
.A1(n_4008),
.A2(n_1091),
.B(n_1102),
.C(n_1082),
.Y(n_4387)
);

INVx3_ASAP7_75t_L g4388 ( 
.A(n_4188),
.Y(n_4388)
);

INVx1_ASAP7_75t_L g4389 ( 
.A(n_4062),
.Y(n_4389)
);

BUFx6f_ASAP7_75t_L g4390 ( 
.A(n_4065),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_3946),
.A2(n_3425),
.B(n_3717),
.Y(n_4391)
);

AO32x1_ASAP7_75t_L g4392 ( 
.A1(n_3954),
.A2(n_1105),
.A3(n_1111),
.B1(n_1107),
.B2(n_1102),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_4128),
.B(n_3704),
.Y(n_4393)
);

AOI22xp33_ASAP7_75t_L g4394 ( 
.A1(n_3946),
.A2(n_1056),
.B1(n_1103),
.B2(n_1042),
.Y(n_4394)
);

AOI21xp33_ASAP7_75t_L g4395 ( 
.A1(n_4092),
.A2(n_3927),
.B(n_3541),
.Y(n_4395)
);

BUFx6f_ASAP7_75t_L g4396 ( 
.A(n_4095),
.Y(n_4396)
);

AOI21xp5_ASAP7_75t_L g4397 ( 
.A1(n_4072),
.A2(n_3465),
.B(n_3379),
.Y(n_4397)
);

NOR2x1_ASAP7_75t_SL g4398 ( 
.A(n_4049),
.B(n_3541),
.Y(n_4398)
);

INVxp67_ASAP7_75t_SL g4399 ( 
.A(n_4132),
.Y(n_4399)
);

NAND2xp5_ASAP7_75t_L g4400 ( 
.A(n_4091),
.B(n_3722),
.Y(n_4400)
);

BUFx2_ASAP7_75t_SL g4401 ( 
.A(n_4068),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_SL g4402 ( 
.A(n_4079),
.B(n_4205),
.Y(n_4402)
);

AOI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_4197),
.A2(n_4200),
.B(n_4195),
.Y(n_4403)
);

A2O1A1Ixp33_ASAP7_75t_L g4404 ( 
.A1(n_4197),
.A2(n_1107),
.B(n_1111),
.C(n_1105),
.Y(n_4404)
);

BUFx2_ASAP7_75t_L g4405 ( 
.A(n_4184),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_4179),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4181),
.Y(n_4407)
);

AND2x2_ASAP7_75t_L g4408 ( 
.A(n_4059),
.B(n_3722),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_4056),
.B(n_3722),
.Y(n_4409)
);

NAND2xp5_ASAP7_75t_L g4410 ( 
.A(n_4057),
.B(n_888),
.Y(n_4410)
);

AOI21xp5_ASAP7_75t_L g4411 ( 
.A1(n_4067),
.A2(n_3112),
.B(n_3089),
.Y(n_4411)
);

OR2x2_ASAP7_75t_L g4412 ( 
.A(n_4101),
.B(n_1550),
.Y(n_4412)
);

NOR2xp33_ASAP7_75t_L g4413 ( 
.A(n_4069),
.B(n_889),
.Y(n_4413)
);

NAND2xp5_ASAP7_75t_SL g4414 ( 
.A(n_4079),
.B(n_2822),
.Y(n_4414)
);

CKINVDCx8_ASAP7_75t_R g4415 ( 
.A(n_4133),
.Y(n_4415)
);

INVx3_ASAP7_75t_L g4416 ( 
.A(n_4186),
.Y(n_4416)
);

BUFx2_ASAP7_75t_L g4417 ( 
.A(n_4137),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_4067),
.B(n_4077),
.Y(n_4418)
);

OAI21x1_ASAP7_75t_L g4419 ( 
.A1(n_4189),
.A2(n_3406),
.B(n_3213),
.Y(n_4419)
);

CKINVDCx5p33_ASAP7_75t_R g4420 ( 
.A(n_4070),
.Y(n_4420)
);

BUFx5_ASAP7_75t_L g4421 ( 
.A(n_4077),
.Y(n_4421)
);

HB1xp67_ASAP7_75t_L g4422 ( 
.A(n_4035),
.Y(n_4422)
);

BUFx2_ASAP7_75t_L g4423 ( 
.A(n_4148),
.Y(n_4423)
);

BUFx6f_ASAP7_75t_L g4424 ( 
.A(n_4034),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_4182),
.Y(n_4425)
);

INVx2_ASAP7_75t_L g4426 ( 
.A(n_4183),
.Y(n_4426)
);

NOR2xp33_ASAP7_75t_SL g4427 ( 
.A(n_4161),
.B(n_3060),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4046),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_4037),
.B(n_892),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4134),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4185),
.Y(n_4431)
);

INVx2_ASAP7_75t_L g4432 ( 
.A(n_4030),
.Y(n_4432)
);

OAI22xp5_ASAP7_75t_L g4433 ( 
.A1(n_4150),
.A2(n_3551),
.B1(n_3256),
.B2(n_3280),
.Y(n_4433)
);

BUFx3_ASAP7_75t_L g4434 ( 
.A(n_4094),
.Y(n_4434)
);

AOI22xp33_ASAP7_75t_SL g4435 ( 
.A1(n_4063),
.A2(n_1110),
.B1(n_1126),
.B2(n_1103),
.Y(n_4435)
);

INVx2_ASAP7_75t_L g4436 ( 
.A(n_4032),
.Y(n_4436)
);

OAI22xp5_ASAP7_75t_L g4437 ( 
.A1(n_4108),
.A2(n_3256),
.B1(n_3280),
.B2(n_3260),
.Y(n_4437)
);

OR2x6_ASAP7_75t_L g4438 ( 
.A(n_4135),
.B(n_3213),
.Y(n_4438)
);

A2O1A1Ixp33_ASAP7_75t_L g4439 ( 
.A1(n_4063),
.A2(n_1117),
.B(n_1119),
.C(n_1114),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4121),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_L g4441 ( 
.A(n_4042),
.B(n_895),
.Y(n_4441)
);

NAND2xp5_ASAP7_75t_SL g4442 ( 
.A(n_4075),
.B(n_2839),
.Y(n_4442)
);

NAND2xp5_ASAP7_75t_L g4443 ( 
.A(n_4043),
.B(n_899),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_SL g4444 ( 
.A(n_4136),
.B(n_2840),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4199),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4199),
.Y(n_4446)
);

NAND2xp5_ASAP7_75t_L g4447 ( 
.A(n_4044),
.B(n_902),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_SL g4448 ( 
.A(n_4113),
.B(n_2859),
.Y(n_4448)
);

OAI22xp5_ASAP7_75t_L g4449 ( 
.A1(n_4098),
.A2(n_3260),
.B1(n_905),
.B2(n_907),
.Y(n_4449)
);

BUFx3_ASAP7_75t_L g4450 ( 
.A(n_4125),
.Y(n_4450)
);

BUFx2_ASAP7_75t_L g4451 ( 
.A(n_4029),
.Y(n_4451)
);

INVx5_ASAP7_75t_L g4452 ( 
.A(n_4029),
.Y(n_4452)
);

BUFx5_ASAP7_75t_L g4453 ( 
.A(n_4131),
.Y(n_4453)
);

CKINVDCx12_ASAP7_75t_R g4454 ( 
.A(n_4295),
.Y(n_4454)
);

NAND2xp5_ASAP7_75t_SL g4455 ( 
.A(n_4290),
.B(n_4129),
.Y(n_4455)
);

AOI21xp5_ASAP7_75t_L g4456 ( 
.A1(n_4418),
.A2(n_4106),
.B(n_4040),
.Y(n_4456)
);

OAI21x1_ASAP7_75t_L g4457 ( 
.A1(n_4242),
.A2(n_4140),
.B(n_4100),
.Y(n_4457)
);

HB1xp67_ASAP7_75t_L g4458 ( 
.A(n_4284),
.Y(n_4458)
);

AO32x2_ASAP7_75t_L g4459 ( 
.A1(n_4289),
.A2(n_4192),
.A3(n_4040),
.B1(n_4123),
.B2(n_4116),
.Y(n_4459)
);

O2A1O1Ixp33_ASAP7_75t_L g4460 ( 
.A1(n_4234),
.A2(n_4112),
.B(n_1117),
.C(n_1124),
.Y(n_4460)
);

AO31x2_ASAP7_75t_L g4461 ( 
.A1(n_4398),
.A2(n_2485),
.A3(n_2481),
.B(n_2466),
.Y(n_4461)
);

OAI21x1_ASAP7_75t_L g4462 ( 
.A1(n_4297),
.A2(n_4120),
.B(n_4119),
.Y(n_4462)
);

NAND2xp33_ASAP7_75t_L g4463 ( 
.A(n_4257),
.B(n_3060),
.Y(n_4463)
);

OAI21x1_ASAP7_75t_L g4464 ( 
.A1(n_4419),
.A2(n_4127),
.B(n_4126),
.Y(n_4464)
);

AOI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_4330),
.A2(n_3112),
.B(n_3082),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_4347),
.A2(n_3089),
.B(n_3075),
.Y(n_4466)
);

OAI21xp5_ASAP7_75t_L g4467 ( 
.A1(n_4209),
.A2(n_1119),
.B(n_1114),
.Y(n_4467)
);

OAI21x1_ASAP7_75t_L g4468 ( 
.A1(n_4411),
.A2(n_2773),
.B(n_2485),
.Y(n_4468)
);

A2O1A1Ixp33_ASAP7_75t_L g4469 ( 
.A1(n_4318),
.A2(n_1127),
.B(n_1128),
.C(n_1124),
.Y(n_4469)
);

AO31x2_ASAP7_75t_L g4470 ( 
.A1(n_4398),
.A2(n_2481),
.A3(n_2466),
.B(n_2456),
.Y(n_4470)
);

INVx2_ASAP7_75t_L g4471 ( 
.A(n_4208),
.Y(n_4471)
);

O2A1O1Ixp33_ASAP7_75t_SL g4472 ( 
.A1(n_4268),
.A2(n_4439),
.B(n_4292),
.C(n_4404),
.Y(n_4472)
);

A2O1A1Ixp33_ASAP7_75t_L g4473 ( 
.A1(n_4403),
.A2(n_4435),
.B(n_4280),
.C(n_4371),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4342),
.Y(n_4474)
);

AOI21xp5_ASAP7_75t_L g4475 ( 
.A1(n_4254),
.A2(n_2773),
.B(n_2842),
.Y(n_4475)
);

NAND2xp5_ASAP7_75t_L g4476 ( 
.A(n_4236),
.B(n_903),
.Y(n_4476)
);

INVx1_ASAP7_75t_L g4477 ( 
.A(n_4358),
.Y(n_4477)
);

OAI21x1_ASAP7_75t_L g4478 ( 
.A1(n_4333),
.A2(n_2773),
.B(n_2800),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4214),
.B(n_908),
.Y(n_4479)
);

NAND2xp5_ASAP7_75t_L g4480 ( 
.A(n_4313),
.B(n_910),
.Y(n_4480)
);

AOI21xp5_ASAP7_75t_L g4481 ( 
.A1(n_4235),
.A2(n_2848),
.B(n_2842),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_SL g4482 ( 
.A(n_4314),
.B(n_1555),
.Y(n_4482)
);

NAND3xp33_ASAP7_75t_SL g4483 ( 
.A(n_4332),
.B(n_912),
.C(n_911),
.Y(n_4483)
);

AND2x2_ASAP7_75t_L g4484 ( 
.A(n_4221),
.B(n_1127),
.Y(n_4484)
);

A2O1A1Ixp33_ASAP7_75t_L g4485 ( 
.A1(n_4345),
.A2(n_1131),
.B(n_1134),
.C(n_1128),
.Y(n_4485)
);

BUFx6f_ASAP7_75t_L g4486 ( 
.A(n_4273),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_4238),
.B(n_913),
.Y(n_4487)
);

AOI22xp5_ASAP7_75t_L g4488 ( 
.A1(n_4245),
.A2(n_918),
.B1(n_922),
.B2(n_914),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_SL g4489 ( 
.A(n_4273),
.B(n_1557),
.Y(n_4489)
);

AOI21xp5_ASAP7_75t_L g4490 ( 
.A1(n_4211),
.A2(n_2848),
.B(n_2842),
.Y(n_4490)
);

AND2x2_ASAP7_75t_L g4491 ( 
.A(n_4256),
.B(n_1131),
.Y(n_4491)
);

INVx2_ASAP7_75t_L g4492 ( 
.A(n_4206),
.Y(n_4492)
);

NAND2x1p5_ASAP7_75t_L g4493 ( 
.A(n_4368),
.B(n_2800),
.Y(n_4493)
);

INVx3_ASAP7_75t_L g4494 ( 
.A(n_4216),
.Y(n_4494)
);

INVx2_ASAP7_75t_L g4495 ( 
.A(n_4291),
.Y(n_4495)
);

OAI21x1_ASAP7_75t_L g4496 ( 
.A1(n_4391),
.A2(n_2811),
.B(n_2800),
.Y(n_4496)
);

AO32x2_ASAP7_75t_L g4497 ( 
.A1(n_4285),
.A2(n_1206),
.A3(n_1126),
.B1(n_1110),
.B2(n_1138),
.Y(n_4497)
);

INVx1_ASAP7_75t_L g4498 ( 
.A(n_4356),
.Y(n_4498)
);

BUFx2_ASAP7_75t_L g4499 ( 
.A(n_4273),
.Y(n_4499)
);

OAI22xp5_ASAP7_75t_L g4500 ( 
.A1(n_4278),
.A2(n_1138),
.B1(n_1141),
.B2(n_1134),
.Y(n_4500)
);

OAI21x1_ASAP7_75t_L g4501 ( 
.A1(n_4397),
.A2(n_2813),
.B(n_2811),
.Y(n_4501)
);

AOI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_4338),
.A2(n_2848),
.B(n_2842),
.Y(n_4502)
);

AOI21xp5_ASAP7_75t_L g4503 ( 
.A1(n_4368),
.A2(n_2848),
.B(n_2813),
.Y(n_4503)
);

AND2x2_ASAP7_75t_L g4504 ( 
.A(n_4230),
.B(n_1141),
.Y(n_4504)
);

OAI22x1_ASAP7_75t_L g4505 ( 
.A1(n_4264),
.A2(n_1152),
.B1(n_1156),
.B2(n_1148),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4321),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4323),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4249),
.Y(n_4508)
);

O2A1O1Ixp33_ASAP7_75t_L g4509 ( 
.A1(n_4248),
.A2(n_1152),
.B(n_1156),
.C(n_1148),
.Y(n_4509)
);

AO31x2_ASAP7_75t_L g4510 ( 
.A1(n_4325),
.A2(n_2456),
.A3(n_1158),
.B(n_1162),
.Y(n_4510)
);

BUFx3_ASAP7_75t_L g4511 ( 
.A(n_4222),
.Y(n_4511)
);

HB1xp67_ASAP7_75t_L g4512 ( 
.A(n_4255),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_4227),
.B(n_923),
.Y(n_4513)
);

INVx1_ASAP7_75t_L g4514 ( 
.A(n_4373),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4210),
.Y(n_4515)
);

AOI21xp5_ASAP7_75t_L g4516 ( 
.A1(n_4368),
.A2(n_2813),
.B(n_2811),
.Y(n_4516)
);

AOI221xp5_ASAP7_75t_L g4517 ( 
.A1(n_4394),
.A2(n_928),
.B1(n_932),
.B2(n_927),
.C(n_924),
.Y(n_4517)
);

BUFx3_ASAP7_75t_L g4518 ( 
.A(n_4222),
.Y(n_4518)
);

OAI21xp5_ASAP7_75t_L g4519 ( 
.A1(n_4372),
.A2(n_1159),
.B(n_1158),
.Y(n_4519)
);

AOI21xp5_ASAP7_75t_L g4520 ( 
.A1(n_4374),
.A2(n_2831),
.B(n_2802),
.Y(n_4520)
);

A2O1A1Ixp33_ASAP7_75t_L g4521 ( 
.A1(n_4413),
.A2(n_1162),
.B(n_1164),
.C(n_1159),
.Y(n_4521)
);

AO31x2_ASAP7_75t_L g4522 ( 
.A1(n_4445),
.A2(n_1164),
.A3(n_1181),
.B(n_1165),
.Y(n_4522)
);

BUFx3_ASAP7_75t_L g4523 ( 
.A(n_4223),
.Y(n_4523)
);

OAI21x1_ASAP7_75t_L g4524 ( 
.A1(n_4266),
.A2(n_2831),
.B(n_2780),
.Y(n_4524)
);

AOI221xp5_ASAP7_75t_SL g4525 ( 
.A1(n_4387),
.A2(n_1181),
.B1(n_1195),
.B2(n_1188),
.C(n_1165),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_4299),
.B(n_933),
.Y(n_4526)
);

OAI21x1_ASAP7_75t_L g4527 ( 
.A1(n_4322),
.A2(n_2831),
.B(n_2780),
.Y(n_4527)
);

AO21x2_ASAP7_75t_L g4528 ( 
.A1(n_4395),
.A2(n_1562),
.B(n_1561),
.Y(n_4528)
);

OAI22xp5_ASAP7_75t_L g4529 ( 
.A1(n_4276),
.A2(n_1195),
.B1(n_1198),
.B2(n_1188),
.Y(n_4529)
);

AND2x4_ASAP7_75t_L g4530 ( 
.A(n_4230),
.B(n_1563),
.Y(n_4530)
);

OAI21xp5_ASAP7_75t_L g4531 ( 
.A1(n_4381),
.A2(n_1200),
.B(n_1198),
.Y(n_4531)
);

OAI22x1_ASAP7_75t_L g4532 ( 
.A1(n_4296),
.A2(n_1205),
.B1(n_1219),
.B2(n_1200),
.Y(n_4532)
);

AOI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4374),
.A2(n_2802),
.B(n_2762),
.Y(n_4533)
);

A2O1A1Ixp33_ASAP7_75t_L g4534 ( 
.A1(n_4357),
.A2(n_1210),
.B(n_1219),
.C(n_1205),
.Y(n_4534)
);

AOI21xp5_ASAP7_75t_L g4535 ( 
.A1(n_4374),
.A2(n_2833),
.B(n_2802),
.Y(n_4535)
);

O2A1O1Ixp33_ASAP7_75t_SL g4536 ( 
.A1(n_4302),
.A2(n_4335),
.B(n_4270),
.C(n_4365),
.Y(n_4536)
);

OR2x2_ASAP7_75t_L g4537 ( 
.A(n_4237),
.B(n_1565),
.Y(n_4537)
);

AOI21xp5_ASAP7_75t_L g4538 ( 
.A1(n_4427),
.A2(n_2833),
.B(n_2802),
.Y(n_4538)
);

OAI21x1_ASAP7_75t_L g4539 ( 
.A1(n_4277),
.A2(n_2782),
.B(n_2777),
.Y(n_4539)
);

OAI21xp5_ASAP7_75t_SL g4540 ( 
.A1(n_4225),
.A2(n_1210),
.B(n_1566),
.Y(n_4540)
);

BUFx10_ASAP7_75t_L g4541 ( 
.A(n_4303),
.Y(n_4541)
);

AO31x2_ASAP7_75t_L g4542 ( 
.A1(n_4446),
.A2(n_2782),
.A3(n_2783),
.B(n_2777),
.Y(n_4542)
);

AO31x2_ASAP7_75t_L g4543 ( 
.A1(n_4380),
.A2(n_2787),
.A3(n_2791),
.B(n_2783),
.Y(n_4543)
);

OAI22xp5_ASAP7_75t_L g4544 ( 
.A1(n_4420),
.A2(n_937),
.B1(n_938),
.B2(n_936),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4414),
.A2(n_2834),
.B(n_2833),
.Y(n_4545)
);

OAI21x1_ASAP7_75t_L g4546 ( 
.A1(n_4312),
.A2(n_2791),
.B(n_2787),
.Y(n_4546)
);

A2O1A1Ixp33_ASAP7_75t_L g4547 ( 
.A1(n_4351),
.A2(n_940),
.B(n_942),
.C(n_939),
.Y(n_4547)
);

NAND2xp33_ASAP7_75t_L g4548 ( 
.A(n_4421),
.B(n_3060),
.Y(n_4548)
);

AO31x2_ASAP7_75t_L g4549 ( 
.A1(n_4433),
.A2(n_2796),
.A3(n_2793),
.B(n_1567),
.Y(n_4549)
);

OAI21x1_ASAP7_75t_L g4550 ( 
.A1(n_4437),
.A2(n_2796),
.B(n_2793),
.Y(n_4550)
);

A2O1A1Ixp33_ASAP7_75t_L g4551 ( 
.A1(n_4369),
.A2(n_951),
.B(n_952),
.C(n_943),
.Y(n_4551)
);

AOI21xp5_ASAP7_75t_L g4552 ( 
.A1(n_4402),
.A2(n_2834),
.B(n_2833),
.Y(n_4552)
);

OAI22xp5_ASAP7_75t_L g4553 ( 
.A1(n_4216),
.A2(n_4415),
.B1(n_4294),
.B2(n_4452),
.Y(n_4553)
);

AOI21xp5_ASAP7_75t_L g4554 ( 
.A1(n_4452),
.A2(n_2841),
.B(n_2834),
.Y(n_4554)
);

INVx4_ASAP7_75t_L g4555 ( 
.A(n_4307),
.Y(n_4555)
);

INVx1_ASAP7_75t_L g4556 ( 
.A(n_4378),
.Y(n_4556)
);

OAI21xp5_ASAP7_75t_L g4557 ( 
.A1(n_4410),
.A2(n_4337),
.B(n_4412),
.Y(n_4557)
);

O2A1O1Ixp33_ASAP7_75t_L g4558 ( 
.A1(n_4219),
.A2(n_1574),
.B(n_1578),
.C(n_1569),
.Y(n_4558)
);

INVx3_ASAP7_75t_L g4559 ( 
.A(n_4269),
.Y(n_4559)
);

AOI21xp5_ASAP7_75t_L g4560 ( 
.A1(n_4452),
.A2(n_2841),
.B(n_2834),
.Y(n_4560)
);

AOI22xp33_ASAP7_75t_L g4561 ( 
.A1(n_4287),
.A2(n_1126),
.B1(n_1206),
.B2(n_1110),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4344),
.Y(n_4562)
);

AO32x2_ASAP7_75t_L g4563 ( 
.A1(n_4282),
.A2(n_4267),
.A3(n_4352),
.B1(n_4328),
.B2(n_4311),
.Y(n_4563)
);

BUFx3_ASAP7_75t_L g4564 ( 
.A(n_4279),
.Y(n_4564)
);

A2O1A1Ixp33_ASAP7_75t_L g4565 ( 
.A1(n_4315),
.A2(n_954),
.B(n_955),
.C(n_953),
.Y(n_4565)
);

OA21x2_ASAP7_75t_L g4566 ( 
.A1(n_4379),
.A2(n_1580),
.B(n_1579),
.Y(n_4566)
);

A2O1A1Ixp33_ASAP7_75t_L g4567 ( 
.A1(n_4389),
.A2(n_957),
.B(n_958),
.C(n_956),
.Y(n_4567)
);

O2A1O1Ixp33_ASAP7_75t_SL g4568 ( 
.A1(n_4310),
.A2(n_1582),
.B(n_1589),
.C(n_1586),
.Y(n_4568)
);

OAI21x1_ASAP7_75t_L g4569 ( 
.A1(n_4442),
.A2(n_2771),
.B(n_2769),
.Y(n_4569)
);

NOR2xp67_ASAP7_75t_L g4570 ( 
.A(n_4329),
.B(n_1591),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4212),
.B(n_4218),
.Y(n_4571)
);

BUFx2_ASAP7_75t_L g4572 ( 
.A(n_4213),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_4259),
.A2(n_2841),
.B(n_2447),
.Y(n_4573)
);

A2O1A1Ixp33_ASAP7_75t_L g4574 ( 
.A1(n_4451),
.A2(n_967),
.B(n_968),
.C(n_966),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4359),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4349),
.Y(n_4576)
);

NAND2x1p5_ASAP7_75t_L g4577 ( 
.A(n_4311),
.B(n_2769),
.Y(n_4577)
);

INVx3_ASAP7_75t_L g4578 ( 
.A(n_4269),
.Y(n_4578)
);

OAI22xp5_ASAP7_75t_L g4579 ( 
.A1(n_4259),
.A2(n_972),
.B1(n_973),
.B2(n_971),
.Y(n_4579)
);

AOI21xp5_ASAP7_75t_L g4580 ( 
.A1(n_4343),
.A2(n_2447),
.B(n_2769),
.Y(n_4580)
);

A2O1A1Ixp33_ASAP7_75t_L g4581 ( 
.A1(n_4362),
.A2(n_975),
.B(n_980),
.C(n_974),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_4274),
.B(n_981),
.Y(n_4582)
);

OAI21x1_ASAP7_75t_L g4583 ( 
.A1(n_4388),
.A2(n_2775),
.B(n_2771),
.Y(n_4583)
);

AOI21xp5_ASAP7_75t_L g4584 ( 
.A1(n_4224),
.A2(n_2447),
.B(n_2771),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4286),
.B(n_982),
.Y(n_4585)
);

AO31x2_ASAP7_75t_L g4586 ( 
.A1(n_4350),
.A2(n_1592),
.A3(n_1596),
.B(n_1595),
.Y(n_4586)
);

OAI21x1_ASAP7_75t_L g4587 ( 
.A1(n_4388),
.A2(n_2792),
.B(n_2775),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4317),
.B(n_983),
.Y(n_4588)
);

INVx2_ASAP7_75t_SL g4589 ( 
.A(n_4269),
.Y(n_4589)
);

CKINVDCx5p33_ASAP7_75t_R g4590 ( 
.A(n_4262),
.Y(n_4590)
);

AOI22xp33_ASAP7_75t_L g4591 ( 
.A1(n_4367),
.A2(n_1126),
.B1(n_1206),
.B2(n_1110),
.Y(n_4591)
);

OAI21x1_ASAP7_75t_L g4592 ( 
.A1(n_4246),
.A2(n_2792),
.B(n_2775),
.Y(n_4592)
);

AOI221x1_ASAP7_75t_L g4593 ( 
.A1(n_4440),
.A2(n_1598),
.B1(n_1604),
.B2(n_1603),
.C(n_1597),
.Y(n_4593)
);

NOR2xp33_ASAP7_75t_L g4594 ( 
.A(n_4226),
.B(n_984),
.Y(n_4594)
);

INVxp67_ASAP7_75t_L g4595 ( 
.A(n_4283),
.Y(n_4595)
);

NOR3xp33_ASAP7_75t_L g4596 ( 
.A(n_4298),
.B(n_1610),
.C(n_1606),
.Y(n_4596)
);

BUFx6f_ASAP7_75t_L g4597 ( 
.A(n_4279),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_SL g4598 ( 
.A(n_4293),
.B(n_1613),
.Y(n_4598)
);

INVxp67_ASAP7_75t_SL g4599 ( 
.A(n_4430),
.Y(n_4599)
);

CKINVDCx11_ASAP7_75t_R g4600 ( 
.A(n_4279),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4228),
.B(n_987),
.Y(n_4601)
);

AO31x2_ASAP7_75t_L g4602 ( 
.A1(n_4353),
.A2(n_1615),
.A3(n_1619),
.B(n_1618),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4250),
.B(n_1620),
.Y(n_4603)
);

AOI21xp5_ASAP7_75t_L g4604 ( 
.A1(n_4231),
.A2(n_2447),
.B(n_2792),
.Y(n_4604)
);

AO31x2_ASAP7_75t_L g4605 ( 
.A1(n_4267),
.A2(n_1623),
.A3(n_1628),
.B(n_1626),
.Y(n_4605)
);

OAI21x1_ASAP7_75t_L g4606 ( 
.A1(n_4247),
.A2(n_2460),
.B(n_1640),
.Y(n_4606)
);

NAND3xp33_ASAP7_75t_SL g4607 ( 
.A(n_4429),
.B(n_992),
.C(n_988),
.Y(n_4607)
);

OAI21x1_ASAP7_75t_L g4608 ( 
.A1(n_4265),
.A2(n_2460),
.B(n_1644),
.Y(n_4608)
);

NOR2xp33_ASAP7_75t_SL g4609 ( 
.A(n_4331),
.B(n_1206),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4432),
.Y(n_4610)
);

BUFx6f_ASAP7_75t_L g4611 ( 
.A(n_4308),
.Y(n_4611)
);

AND2x2_ASAP7_75t_L g4612 ( 
.A(n_4250),
.B(n_4215),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4436),
.Y(n_4613)
);

AO21x2_ASAP7_75t_L g4614 ( 
.A1(n_4448),
.A2(n_1658),
.B(n_1655),
.Y(n_4614)
);

BUFx3_ASAP7_75t_L g4615 ( 
.A(n_4390),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4215),
.B(n_1630),
.Y(n_4616)
);

INVx1_ASAP7_75t_SL g4617 ( 
.A(n_4232),
.Y(n_4617)
);

BUFx6f_ASAP7_75t_L g4618 ( 
.A(n_4308),
.Y(n_4618)
);

CKINVDCx5p33_ASAP7_75t_R g4619 ( 
.A(n_4331),
.Y(n_4619)
);

AOI21xp5_ASAP7_75t_L g4620 ( 
.A1(n_4298),
.A2(n_2447),
.B(n_2129),
.Y(n_4620)
);

BUFx2_ASAP7_75t_L g4621 ( 
.A(n_4213),
.Y(n_4621)
);

OAI22xp5_ASAP7_75t_L g4622 ( 
.A1(n_4334),
.A2(n_995),
.B1(n_998),
.B2(n_993),
.Y(n_4622)
);

AO31x2_ASAP7_75t_L g4623 ( 
.A1(n_4348),
.A2(n_1645),
.A3(n_1647),
.B(n_1646),
.Y(n_4623)
);

OAI22xp5_ASAP7_75t_L g4624 ( 
.A1(n_4334),
.A2(n_1005),
.B1(n_1006),
.B2(n_1002),
.Y(n_4624)
);

A2O1A1Ixp33_ASAP7_75t_L g4625 ( 
.A1(n_4346),
.A2(n_1007),
.B(n_1013),
.C(n_1009),
.Y(n_4625)
);

NAND3x1_ASAP7_75t_L g4626 ( 
.A(n_4305),
.B(n_1650),
.C(n_1649),
.Y(n_4626)
);

BUFx6f_ASAP7_75t_L g4627 ( 
.A(n_4308),
.Y(n_4627)
);

O2A1O1Ixp5_ASAP7_75t_SL g4628 ( 
.A1(n_4428),
.A2(n_1651),
.B(n_1660),
.C(n_1004),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4399),
.B(n_1014),
.Y(n_4629)
);

O2A1O1Ixp33_ASAP7_75t_L g4630 ( 
.A1(n_4207),
.A2(n_1019),
.B(n_1020),
.C(n_1016),
.Y(n_4630)
);

NOR2xp33_ASAP7_75t_L g4631 ( 
.A(n_4220),
.B(n_1022),
.Y(n_4631)
);

AND2x4_ASAP7_75t_L g4632 ( 
.A(n_4239),
.B(n_631),
.Y(n_4632)
);

INVx3_ASAP7_75t_SL g4633 ( 
.A(n_4366),
.Y(n_4633)
);

NOR2xp33_ASAP7_75t_L g4634 ( 
.A(n_4400),
.B(n_1024),
.Y(n_4634)
);

INVx3_ASAP7_75t_L g4635 ( 
.A(n_4390),
.Y(n_4635)
);

OAI21x1_ASAP7_75t_L g4636 ( 
.A1(n_4326),
.A2(n_633),
.B(n_632),
.Y(n_4636)
);

OAI21x1_ASAP7_75t_L g4637 ( 
.A1(n_4251),
.A2(n_640),
.B(n_637),
.Y(n_4637)
);

INVx2_ASAP7_75t_SL g4638 ( 
.A(n_4253),
.Y(n_4638)
);

AOI21xp5_ASAP7_75t_L g4639 ( 
.A1(n_4360),
.A2(n_4444),
.B(n_4316),
.Y(n_4639)
);

OAI22x1_ASAP7_75t_L g4640 ( 
.A1(n_4422),
.A2(n_1050),
.B1(n_1069),
.B2(n_1031),
.Y(n_4640)
);

BUFx3_ASAP7_75t_L g4641 ( 
.A(n_4390),
.Y(n_4641)
);

AND2x2_ASAP7_75t_L g4642 ( 
.A(n_4239),
.B(n_6),
.Y(n_4642)
);

NOR2xp33_ASAP7_75t_L g4643 ( 
.A(n_4441),
.B(n_1034),
.Y(n_4643)
);

NOR3xp33_ASAP7_75t_L g4644 ( 
.A(n_4304),
.B(n_1037),
.C(n_1035),
.Y(n_4644)
);

AO31x2_ASAP7_75t_L g4645 ( 
.A1(n_4355),
.A2(n_4377),
.A3(n_4382),
.B(n_4376),
.Y(n_4645)
);

A2O1A1Ixp33_ASAP7_75t_L g4646 ( 
.A1(n_4364),
.A2(n_1041),
.B(n_1045),
.C(n_1038),
.Y(n_4646)
);

BUFx2_ASAP7_75t_R g4647 ( 
.A(n_4401),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4316),
.A2(n_1051),
.B(n_1049),
.Y(n_4648)
);

AOI21xp5_ASAP7_75t_L g4649 ( 
.A1(n_4416),
.A2(n_1054),
.B(n_1052),
.Y(n_4649)
);

A2O1A1Ixp33_ASAP7_75t_L g4650 ( 
.A1(n_4272),
.A2(n_1060),
.B(n_1061),
.C(n_1055),
.Y(n_4650)
);

INVx2_ASAP7_75t_SL g4651 ( 
.A(n_4253),
.Y(n_4651)
);

NAND2x1p5_ASAP7_75t_L g4652 ( 
.A(n_4281),
.B(n_641),
.Y(n_4652)
);

INVx2_ASAP7_75t_L g4653 ( 
.A(n_4240),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4233),
.Y(n_4654)
);

AOI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4416),
.A2(n_1070),
.B(n_1067),
.Y(n_4655)
);

AOI221xp5_ASAP7_75t_SL g4656 ( 
.A1(n_4401),
.A2(n_1080),
.B1(n_1085),
.B2(n_1079),
.C(n_1072),
.Y(n_4656)
);

AO31x2_ASAP7_75t_L g4657 ( 
.A1(n_4385),
.A2(n_9),
.A3(n_7),
.B(n_8),
.Y(n_4657)
);

AND2x2_ASAP7_75t_L g4658 ( 
.A(n_4229),
.B(n_8),
.Y(n_4658)
);

OAI21x1_ASAP7_75t_SL g4659 ( 
.A1(n_4241),
.A2(n_9),
.B(n_10),
.Y(n_4659)
);

INVx1_ASAP7_75t_SL g4660 ( 
.A(n_4393),
.Y(n_4660)
);

AOI221xp5_ASAP7_75t_SL g4661 ( 
.A1(n_4252),
.A2(n_4447),
.B1(n_4443),
.B2(n_4354),
.C(n_4424),
.Y(n_4661)
);

A2O1A1Ixp33_ASAP7_75t_L g4662 ( 
.A1(n_4417),
.A2(n_1087),
.B(n_1088),
.C(n_1086),
.Y(n_4662)
);

OAI21x1_ASAP7_75t_L g4663 ( 
.A1(n_4406),
.A2(n_643),
.B(n_642),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4300),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4243),
.Y(n_4665)
);

AOI21xp5_ASAP7_75t_L g4666 ( 
.A1(n_4438),
.A2(n_4386),
.B(n_4217),
.Y(n_4666)
);

OAI21x1_ASAP7_75t_SL g4667 ( 
.A1(n_4288),
.A2(n_4409),
.B(n_4340),
.Y(n_4667)
);

AOI22xp33_ASAP7_75t_L g4668 ( 
.A1(n_4275),
.A2(n_1092),
.B1(n_1095),
.B2(n_1090),
.Y(n_4668)
);

INVx2_ASAP7_75t_SL g4669 ( 
.A(n_4424),
.Y(n_4669)
);

AND2x4_ASAP7_75t_L g4670 ( 
.A(n_4229),
.B(n_645),
.Y(n_4670)
);

A2O1A1Ixp33_ASAP7_75t_L g4671 ( 
.A1(n_4423),
.A2(n_4434),
.B(n_4258),
.C(n_4261),
.Y(n_4671)
);

O2A1O1Ixp33_ASAP7_75t_SL g4672 ( 
.A1(n_4370),
.A2(n_4306),
.B(n_4319),
.C(n_4309),
.Y(n_4672)
);

BUFx3_ASAP7_75t_L g4673 ( 
.A(n_4424),
.Y(n_4673)
);

INVx1_ASAP7_75t_SL g4674 ( 
.A(n_4324),
.Y(n_4674)
);

AOI21xp5_ASAP7_75t_SL g4675 ( 
.A1(n_4449),
.A2(n_1097),
.B(n_1096),
.Y(n_4675)
);

AOI21xp5_ASAP7_75t_L g4676 ( 
.A1(n_4438),
.A2(n_1101),
.B(n_1098),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_4339),
.B(n_1104),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4229),
.B(n_11),
.Y(n_4678)
);

O2A1O1Ixp33_ASAP7_75t_L g4679 ( 
.A1(n_4386),
.A2(n_1109),
.B(n_1112),
.C(n_1106),
.Y(n_4679)
);

NAND2x1p5_ASAP7_75t_L g4680 ( 
.A(n_4260),
.B(n_647),
.Y(n_4680)
);

OR2x6_ASAP7_75t_L g4681 ( 
.A(n_4275),
.B(n_648),
.Y(n_4681)
);

AO32x2_ASAP7_75t_L g4682 ( 
.A1(n_4453),
.A2(n_13),
.A3(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_4682)
);

OA21x2_ASAP7_75t_L g4683 ( 
.A1(n_4407),
.A2(n_1116),
.B(n_1115),
.Y(n_4683)
);

A2O1A1Ixp33_ASAP7_75t_L g4684 ( 
.A1(n_4450),
.A2(n_1125),
.B(n_1129),
.C(n_1123),
.Y(n_4684)
);

AO21x2_ASAP7_75t_L g4685 ( 
.A1(n_4425),
.A2(n_1133),
.B(n_1132),
.Y(n_4685)
);

AO31x2_ASAP7_75t_L g4686 ( 
.A1(n_4426),
.A2(n_15),
.A3(n_12),
.B(n_13),
.Y(n_4686)
);

OAI21x1_ASAP7_75t_L g4687 ( 
.A1(n_4431),
.A2(n_651),
.B(n_649),
.Y(n_4687)
);

INVx1_ASAP7_75t_L g4688 ( 
.A(n_4453),
.Y(n_4688)
);

INVx2_ASAP7_75t_SL g4689 ( 
.A(n_4307),
.Y(n_4689)
);

OAI21x1_ASAP7_75t_L g4690 ( 
.A1(n_4320),
.A2(n_654),
.B(n_652),
.Y(n_4690)
);

AOI21xp5_ASAP7_75t_L g4691 ( 
.A1(n_4217),
.A2(n_1146),
.B(n_1144),
.Y(n_4691)
);

A2O1A1Ixp33_ASAP7_75t_L g4692 ( 
.A1(n_4375),
.A2(n_4405),
.B(n_4271),
.C(n_4384),
.Y(n_4692)
);

OAI21x1_ASAP7_75t_L g4693 ( 
.A1(n_4327),
.A2(n_657),
.B(n_656),
.Y(n_4693)
);

AO31x2_ASAP7_75t_L g4694 ( 
.A1(n_4341),
.A2(n_19),
.A3(n_16),
.B(n_18),
.Y(n_4694)
);

OAI21x1_ASAP7_75t_L g4695 ( 
.A1(n_4263),
.A2(n_660),
.B(n_658),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4301),
.B(n_4336),
.Y(n_4696)
);

O2A1O1Ixp5_ASAP7_75t_L g4697 ( 
.A1(n_4361),
.A2(n_1150),
.B(n_1154),
.C(n_1147),
.Y(n_4697)
);

NOR2xp33_ASAP7_75t_L g4698 ( 
.A(n_4396),
.B(n_1155),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4562),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4498),
.Y(n_4700)
);

AOI221xp5_ASAP7_75t_L g4701 ( 
.A1(n_4467),
.A2(n_1166),
.B1(n_1168),
.B2(n_1163),
.C(n_1161),
.Y(n_4701)
);

OAI21x1_ASAP7_75t_L g4702 ( 
.A1(n_4475),
.A2(n_4408),
.B(n_4421),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4575),
.Y(n_4703)
);

INVx4_ASAP7_75t_SL g4704 ( 
.A(n_4511),
.Y(n_4704)
);

OAI21x1_ASAP7_75t_L g4705 ( 
.A1(n_4502),
.A2(n_4421),
.B(n_4453),
.Y(n_4705)
);

OAI21x1_ASAP7_75t_L g4706 ( 
.A1(n_4501),
.A2(n_4421),
.B(n_4453),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4506),
.Y(n_4707)
);

OAI21x1_ASAP7_75t_L g4708 ( 
.A1(n_4496),
.A2(n_4453),
.B(n_4217),
.Y(n_4708)
);

INVx2_ASAP7_75t_L g4709 ( 
.A(n_4477),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4617),
.B(n_4244),
.Y(n_4710)
);

INVx1_ASAP7_75t_L g4711 ( 
.A(n_4507),
.Y(n_4711)
);

NAND2x1p5_ASAP7_75t_L g4712 ( 
.A(n_4494),
.B(n_4307),
.Y(n_4712)
);

BUFx6f_ASAP7_75t_L g4713 ( 
.A(n_4600),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4514),
.Y(n_4714)
);

BUFx6f_ASAP7_75t_L g4715 ( 
.A(n_4611),
.Y(n_4715)
);

INVx1_ASAP7_75t_L g4716 ( 
.A(n_4576),
.Y(n_4716)
);

OA21x2_ASAP7_75t_L g4717 ( 
.A1(n_4661),
.A2(n_4366),
.B(n_4363),
.Y(n_4717)
);

INVx2_ASAP7_75t_SL g4718 ( 
.A(n_4523),
.Y(n_4718)
);

OAI21xp5_ASAP7_75t_L g4719 ( 
.A1(n_4473),
.A2(n_4361),
.B(n_4363),
.Y(n_4719)
);

BUFx2_ASAP7_75t_SL g4720 ( 
.A(n_4518),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4572),
.B(n_4621),
.Y(n_4721)
);

OAI21x1_ASAP7_75t_L g4722 ( 
.A1(n_4580),
.A2(n_4392),
.B(n_4383),
.Y(n_4722)
);

OAI21x1_ASAP7_75t_L g4723 ( 
.A1(n_4481),
.A2(n_4392),
.B(n_4383),
.Y(n_4723)
);

BUFx4f_ASAP7_75t_SL g4724 ( 
.A(n_4564),
.Y(n_4724)
);

AND2x4_ASAP7_75t_L g4725 ( 
.A(n_4612),
.B(n_4244),
.Y(n_4725)
);

BUFx8_ASAP7_75t_SL g4726 ( 
.A(n_4619),
.Y(n_4726)
);

CKINVDCx20_ASAP7_75t_R g4727 ( 
.A(n_4590),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4556),
.Y(n_4728)
);

OAI21x1_ASAP7_75t_SL g4729 ( 
.A1(n_4667),
.A2(n_4370),
.B(n_4244),
.Y(n_4729)
);

OAI21x1_ASAP7_75t_L g4730 ( 
.A1(n_4604),
.A2(n_4383),
.B(n_4396),
.Y(n_4730)
);

OR2x2_ASAP7_75t_L g4731 ( 
.A(n_4474),
.B(n_4396),
.Y(n_4731)
);

OAI21x1_ASAP7_75t_L g4732 ( 
.A1(n_4592),
.A2(n_4383),
.B(n_666),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4512),
.Y(n_4733)
);

NAND2x1p5_ASAP7_75t_L g4734 ( 
.A(n_4555),
.B(n_663),
.Y(n_4734)
);

NAND2xp5_ASAP7_75t_L g4735 ( 
.A(n_4508),
.B(n_1170),
.Y(n_4735)
);

AO21x2_ASAP7_75t_L g4736 ( 
.A1(n_4596),
.A2(n_16),
.B(n_18),
.Y(n_4736)
);

AO31x2_ASAP7_75t_L g4737 ( 
.A1(n_4593),
.A2(n_4688),
.A3(n_4666),
.B(n_4490),
.Y(n_4737)
);

CKINVDCx20_ASAP7_75t_R g4738 ( 
.A(n_4454),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4458),
.Y(n_4739)
);

INVx3_ASAP7_75t_L g4740 ( 
.A(n_4673),
.Y(n_4740)
);

AO31x2_ASAP7_75t_L g4741 ( 
.A1(n_4639),
.A2(n_22),
.A3(n_20),
.B(n_21),
.Y(n_4741)
);

HB1xp67_ASAP7_75t_L g4742 ( 
.A(n_4645),
.Y(n_4742)
);

OA21x2_ASAP7_75t_L g4743 ( 
.A1(n_4671),
.A2(n_1173),
.B(n_1171),
.Y(n_4743)
);

CKINVDCx5p33_ASAP7_75t_R g4744 ( 
.A(n_4541),
.Y(n_4744)
);

OAI22xp5_ASAP7_75t_L g4745 ( 
.A1(n_4647),
.A2(n_1178),
.B1(n_1180),
.B2(n_1175),
.Y(n_4745)
);

INVx1_ASAP7_75t_L g4746 ( 
.A(n_4471),
.Y(n_4746)
);

INVx2_ASAP7_75t_L g4747 ( 
.A(n_4645),
.Y(n_4747)
);

AND2x4_ASAP7_75t_L g4748 ( 
.A(n_4599),
.B(n_4653),
.Y(n_4748)
);

AO31x2_ASAP7_75t_L g4749 ( 
.A1(n_4584),
.A2(n_22),
.A3(n_20),
.B(n_21),
.Y(n_4749)
);

AO221x1_ASAP7_75t_L g4750 ( 
.A1(n_4553),
.A2(n_4659),
.B1(n_4486),
.B2(n_4505),
.C(n_4682),
.Y(n_4750)
);

AOI21xp5_ASAP7_75t_L g4751 ( 
.A1(n_4548),
.A2(n_1186),
.B(n_1185),
.Y(n_4751)
);

OAI21x1_ASAP7_75t_L g4752 ( 
.A1(n_4457),
.A2(n_672),
.B(n_668),
.Y(n_4752)
);

OAI21xp5_ASAP7_75t_L g4753 ( 
.A1(n_4697),
.A2(n_1190),
.B(n_1187),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4674),
.B(n_23),
.Y(n_4754)
);

HB1xp67_ASAP7_75t_L g4755 ( 
.A(n_4645),
.Y(n_4755)
);

A2O1A1Ixp33_ASAP7_75t_L g4756 ( 
.A1(n_4679),
.A2(n_1220),
.B(n_1194),
.C(n_1196),
.Y(n_4756)
);

NOR2xp33_ASAP7_75t_SL g4757 ( 
.A(n_4652),
.B(n_1192),
.Y(n_4757)
);

OA21x2_ASAP7_75t_L g4758 ( 
.A1(n_4552),
.A2(n_1201),
.B(n_1197),
.Y(n_4758)
);

BUFx2_ASAP7_75t_L g4759 ( 
.A(n_4499),
.Y(n_4759)
);

CKINVDCx8_ASAP7_75t_R g4760 ( 
.A(n_4486),
.Y(n_4760)
);

AOI22xp33_ASAP7_75t_L g4761 ( 
.A1(n_4644),
.A2(n_1203),
.B1(n_1209),
.B2(n_1202),
.Y(n_4761)
);

INVx1_ASAP7_75t_SL g4762 ( 
.A(n_4696),
.Y(n_4762)
);

OAI21x1_ASAP7_75t_L g4763 ( 
.A1(n_4524),
.A2(n_676),
.B(n_674),
.Y(n_4763)
);

BUFx3_ASAP7_75t_L g4764 ( 
.A(n_4615),
.Y(n_4764)
);

INVx1_ASAP7_75t_SL g4765 ( 
.A(n_4660),
.Y(n_4765)
);

AND2x2_ASAP7_75t_L g4766 ( 
.A(n_4595),
.B(n_23),
.Y(n_4766)
);

NAND3xp33_ASAP7_75t_L g4767 ( 
.A(n_4656),
.B(n_4469),
.C(n_4630),
.Y(n_4767)
);

AOI21xp5_ASAP7_75t_L g4768 ( 
.A1(n_4573),
.A2(n_1213),
.B(n_1211),
.Y(n_4768)
);

OAI21x1_ASAP7_75t_L g4769 ( 
.A1(n_4478),
.A2(n_679),
.B(n_678),
.Y(n_4769)
);

OAI22xp5_ASAP7_75t_L g4770 ( 
.A1(n_4692),
.A2(n_1214),
.B1(n_1217),
.B2(n_26),
.Y(n_4770)
);

OA21x2_ASAP7_75t_L g4771 ( 
.A1(n_4462),
.A2(n_24),
.B(n_25),
.Y(n_4771)
);

CKINVDCx5p33_ASAP7_75t_R g4772 ( 
.A(n_4641),
.Y(n_4772)
);

AO31x2_ASAP7_75t_L g4773 ( 
.A1(n_4545),
.A2(n_28),
.A3(n_24),
.B(n_27),
.Y(n_4773)
);

INVx3_ASAP7_75t_L g4774 ( 
.A(n_4654),
.Y(n_4774)
);

HB1xp67_ASAP7_75t_L g4775 ( 
.A(n_4610),
.Y(n_4775)
);

OR2x6_ASAP7_75t_L g4776 ( 
.A(n_4456),
.B(n_682),
.Y(n_4776)
);

CKINVDCx11_ASAP7_75t_R g4777 ( 
.A(n_4597),
.Y(n_4777)
);

AOI22xp33_ASAP7_75t_SL g4778 ( 
.A1(n_4683),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_4778)
);

NOR2xp67_ASAP7_75t_L g4779 ( 
.A(n_4537),
.B(n_29),
.Y(n_4779)
);

NOR2xp33_ASAP7_75t_L g4780 ( 
.A(n_4677),
.B(n_31),
.Y(n_4780)
);

O2A1O1Ixp33_ASAP7_75t_L g4781 ( 
.A1(n_4472),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4664),
.Y(n_4782)
);

OAI21x1_ASAP7_75t_L g4783 ( 
.A1(n_4464),
.A2(n_685),
.B(n_683),
.Y(n_4783)
);

INVx2_ASAP7_75t_L g4784 ( 
.A(n_4515),
.Y(n_4784)
);

AO31x2_ASAP7_75t_L g4785 ( 
.A1(n_4620),
.A2(n_4554),
.A3(n_4560),
.B(n_4535),
.Y(n_4785)
);

OAI21x1_ASAP7_75t_L g4786 ( 
.A1(n_4468),
.A2(n_689),
.B(n_686),
.Y(n_4786)
);

OAI21x1_ASAP7_75t_L g4787 ( 
.A1(n_4539),
.A2(n_693),
.B(n_690),
.Y(n_4787)
);

OAI21x1_ASAP7_75t_L g4788 ( 
.A1(n_4527),
.A2(n_696),
.B(n_694),
.Y(n_4788)
);

AO21x1_ASAP7_75t_L g4789 ( 
.A1(n_4682),
.A2(n_33),
.B(n_35),
.Y(n_4789)
);

BUFx2_ASAP7_75t_L g4790 ( 
.A(n_4633),
.Y(n_4790)
);

AND2x2_ASAP7_75t_L g4791 ( 
.A(n_4635),
.B(n_35),
.Y(n_4791)
);

INVxp67_ASAP7_75t_L g4792 ( 
.A(n_4491),
.Y(n_4792)
);

OAI21x1_ASAP7_75t_L g4793 ( 
.A1(n_4569),
.A2(n_36),
.B(n_39),
.Y(n_4793)
);

OAI21x1_ASAP7_75t_L g4794 ( 
.A1(n_4550),
.A2(n_36),
.B(n_39),
.Y(n_4794)
);

INVx1_ASAP7_75t_L g4795 ( 
.A(n_4665),
.Y(n_4795)
);

OAI21x1_ASAP7_75t_L g4796 ( 
.A1(n_4466),
.A2(n_40),
.B(n_41),
.Y(n_4796)
);

NOR2xp33_ASAP7_75t_L g4797 ( 
.A(n_4634),
.B(n_42),
.Y(n_4797)
);

AO21x1_ASAP7_75t_L g4798 ( 
.A1(n_4682),
.A2(n_44),
.B(n_45),
.Y(n_4798)
);

AND2x4_ASAP7_75t_L g4799 ( 
.A(n_4669),
.B(n_44),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4492),
.Y(n_4800)
);

OAI21xp5_ASAP7_75t_L g4801 ( 
.A1(n_4676),
.A2(n_45),
.B(n_46),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4613),
.B(n_46),
.Y(n_4802)
);

NOR2xp33_ASAP7_75t_L g4803 ( 
.A(n_4631),
.B(n_47),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4495),
.Y(n_4804)
);

CKINVDCx11_ASAP7_75t_R g4805 ( 
.A(n_4597),
.Y(n_4805)
);

AO21x2_ASAP7_75t_L g4806 ( 
.A1(n_4570),
.A2(n_47),
.B(n_49),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_4463),
.A2(n_50),
.B(n_51),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_4522),
.Y(n_4808)
);

OAI21x1_ASAP7_75t_L g4809 ( 
.A1(n_4583),
.A2(n_50),
.B(n_51),
.Y(n_4809)
);

OAI21x1_ASAP7_75t_L g4810 ( 
.A1(n_4587),
.A2(n_52),
.B(n_53),
.Y(n_4810)
);

AOI21xp33_ASAP7_75t_SL g4811 ( 
.A1(n_4640),
.A2(n_52),
.B(n_53),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4522),
.Y(n_4812)
);

AND2x4_ASAP7_75t_L g4813 ( 
.A(n_4638),
.B(n_56),
.Y(n_4813)
);

INVx2_ASAP7_75t_SL g4814 ( 
.A(n_4611),
.Y(n_4814)
);

OAI21x1_ASAP7_75t_L g4815 ( 
.A1(n_4628),
.A2(n_56),
.B(n_57),
.Y(n_4815)
);

OAI21x1_ASAP7_75t_L g4816 ( 
.A1(n_4546),
.A2(n_57),
.B(n_58),
.Y(n_4816)
);

NAND2xp5_ASAP7_75t_L g4817 ( 
.A(n_4571),
.B(n_60),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4651),
.B(n_4504),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4522),
.Y(n_4819)
);

AND2x4_ASAP7_75t_L g4820 ( 
.A(n_4689),
.B(n_61),
.Y(n_4820)
);

AOI22xp5_ASAP7_75t_L g4821 ( 
.A1(n_4525),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4657),
.Y(n_4822)
);

AOI21xp5_ASAP7_75t_L g4823 ( 
.A1(n_4538),
.A2(n_4465),
.B(n_4455),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_L g4824 ( 
.A(n_4484),
.B(n_63),
.Y(n_4824)
);

OAI22xp5_ASAP7_75t_L g4825 ( 
.A1(n_4591),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_4825)
);

AOI221xp5_ASAP7_75t_L g4826 ( 
.A1(n_4540),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.C(n_68),
.Y(n_4826)
);

A2O1A1Ixp33_ASAP7_75t_L g4827 ( 
.A1(n_4557),
.A2(n_4509),
.B(n_4648),
.C(n_4643),
.Y(n_4827)
);

INVxp33_ASAP7_75t_L g4828 ( 
.A(n_4698),
.Y(n_4828)
);

NOR2xp33_ASAP7_75t_L g4829 ( 
.A(n_4588),
.B(n_67),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4559),
.B(n_68),
.Y(n_4830)
);

NAND3xp33_ASAP7_75t_L g4831 ( 
.A(n_4519),
.B(n_71),
.C(n_72),
.Y(n_4831)
);

INVx5_ASAP7_75t_L g4832 ( 
.A(n_4681),
.Y(n_4832)
);

OR2x6_ASAP7_75t_L g4833 ( 
.A(n_4681),
.B(n_73),
.Y(n_4833)
);

OAI21xp5_ASAP7_75t_L g4834 ( 
.A1(n_4625),
.A2(n_73),
.B(n_74),
.Y(n_4834)
);

OAI21x1_ASAP7_75t_L g4835 ( 
.A1(n_4637),
.A2(n_75),
.B(n_76),
.Y(n_4835)
);

AOI21xp33_ASAP7_75t_L g4836 ( 
.A1(n_4683),
.A2(n_77),
.B(n_78),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4542),
.Y(n_4837)
);

OAI21x1_ASAP7_75t_L g4838 ( 
.A1(n_4566),
.A2(n_4636),
.B(n_4608),
.Y(n_4838)
);

OA21x2_ASAP7_75t_L g4839 ( 
.A1(n_4533),
.A2(n_77),
.B(n_79),
.Y(n_4839)
);

INVx3_ASAP7_75t_L g4840 ( 
.A(n_4618),
.Y(n_4840)
);

NOR2xp33_ASAP7_75t_SL g4841 ( 
.A(n_4680),
.B(n_80),
.Y(n_4841)
);

INVx1_ASAP7_75t_SL g4842 ( 
.A(n_4618),
.Y(n_4842)
);

OA21x2_ASAP7_75t_L g4843 ( 
.A1(n_4663),
.A2(n_80),
.B(n_81),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_4483),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_4844)
);

OAI21x1_ASAP7_75t_L g4845 ( 
.A1(n_4566),
.A2(n_83),
.B(n_84),
.Y(n_4845)
);

AND2x2_ASAP7_75t_L g4846 ( 
.A(n_4578),
.B(n_85),
.Y(n_4846)
);

AND2x4_ASAP7_75t_L g4847 ( 
.A(n_4589),
.B(n_86),
.Y(n_4847)
);

OAI21xp5_ASAP7_75t_L g4848 ( 
.A1(n_4646),
.A2(n_86),
.B(n_87),
.Y(n_4848)
);

OAI21x1_ASAP7_75t_L g4849 ( 
.A1(n_4606),
.A2(n_88),
.B(n_89),
.Y(n_4849)
);

CKINVDCx6p67_ASAP7_75t_R g4850 ( 
.A(n_4658),
.Y(n_4850)
);

AOI21xp5_ASAP7_75t_SL g4851 ( 
.A1(n_4598),
.A2(n_90),
.B(n_91),
.Y(n_4851)
);

O2A1O1Ixp33_ASAP7_75t_SL g4852 ( 
.A1(n_4521),
.A2(n_92),
.B(n_90),
.C(n_91),
.Y(n_4852)
);

OAI21x1_ASAP7_75t_L g4853 ( 
.A1(n_4503),
.A2(n_93),
.B(n_94),
.Y(n_4853)
);

OAI21x1_ASAP7_75t_L g4854 ( 
.A1(n_4687),
.A2(n_93),
.B(n_94),
.Y(n_4854)
);

AO21x2_ASAP7_75t_L g4855 ( 
.A1(n_4528),
.A2(n_96),
.B(n_97),
.Y(n_4855)
);

A2O1A1Ixp33_ASAP7_75t_L g4856 ( 
.A1(n_4531),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4657),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4542),
.Y(n_4858)
);

INVx1_ASAP7_75t_L g4859 ( 
.A(n_4542),
.Y(n_4859)
);

BUFx2_ASAP7_75t_L g4860 ( 
.A(n_4627),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4657),
.Y(n_4861)
);

OAI21x1_ASAP7_75t_L g4862 ( 
.A1(n_4690),
.A2(n_98),
.B(n_99),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4686),
.Y(n_4863)
);

OAI21x1_ASAP7_75t_L g4864 ( 
.A1(n_4693),
.A2(n_100),
.B(n_101),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4603),
.B(n_4629),
.Y(n_4865)
);

INVx2_ASAP7_75t_L g4866 ( 
.A(n_4616),
.Y(n_4866)
);

O2A1O1Ixp33_ASAP7_75t_L g4867 ( 
.A1(n_4581),
.A2(n_105),
.B(n_101),
.C(n_103),
.Y(n_4867)
);

AOI22x1_ASAP7_75t_L g4868 ( 
.A1(n_4532),
.A2(n_109),
.B1(n_105),
.B2(n_106),
.Y(n_4868)
);

INVx3_ASAP7_75t_L g4869 ( 
.A(n_4627),
.Y(n_4869)
);

OAI21x1_ASAP7_75t_L g4870 ( 
.A1(n_4520),
.A2(n_106),
.B(n_110),
.Y(n_4870)
);

BUFx10_ASAP7_75t_L g4871 ( 
.A(n_4594),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4686),
.Y(n_4872)
);

AOI21x1_ASAP7_75t_L g4873 ( 
.A1(n_4489),
.A2(n_111),
.B(n_112),
.Y(n_4873)
);

AOI21xp5_ASAP7_75t_L g4874 ( 
.A1(n_4536),
.A2(n_114),
.B(n_115),
.Y(n_4874)
);

OAI21x1_ASAP7_75t_L g4875 ( 
.A1(n_4695),
.A2(n_114),
.B(n_116),
.Y(n_4875)
);

AO31x2_ASAP7_75t_L g4876 ( 
.A1(n_4534),
.A2(n_4516),
.A3(n_4543),
.B(n_4485),
.Y(n_4876)
);

OAI21x1_ASAP7_75t_L g4877 ( 
.A1(n_4626),
.A2(n_116),
.B(n_118),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4678),
.B(n_119),
.Y(n_4878)
);

INVx1_ASAP7_75t_L g4879 ( 
.A(n_4686),
.Y(n_4879)
);

AOI21xp5_ASAP7_75t_L g4880 ( 
.A1(n_4675),
.A2(n_121),
.B(n_122),
.Y(n_4880)
);

OAI21x1_ASAP7_75t_L g4881 ( 
.A1(n_4577),
.A2(n_121),
.B(n_124),
.Y(n_4881)
);

AND2x2_ASAP7_75t_SL g4882 ( 
.A(n_4609),
.B(n_124),
.Y(n_4882)
);

INVx3_ASAP7_75t_L g4883 ( 
.A(n_4530),
.Y(n_4883)
);

INVx2_ASAP7_75t_SL g4884 ( 
.A(n_4530),
.Y(n_4884)
);

HB1xp67_ASAP7_75t_L g4885 ( 
.A(n_4510),
.Y(n_4885)
);

INVx3_ASAP7_75t_SL g4886 ( 
.A(n_4670),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4601),
.B(n_125),
.Y(n_4887)
);

INVx1_ASAP7_75t_L g4888 ( 
.A(n_4694),
.Y(n_4888)
);

OAI21x1_ASAP7_75t_L g4889 ( 
.A1(n_4493),
.A2(n_126),
.B(n_128),
.Y(n_4889)
);

INVx4_ASAP7_75t_L g4890 ( 
.A(n_4632),
.Y(n_4890)
);

OAI21x1_ASAP7_75t_L g4891 ( 
.A1(n_4558),
.A2(n_4642),
.B(n_4460),
.Y(n_4891)
);

HB1xp67_ASAP7_75t_L g4892 ( 
.A(n_4775),
.Y(n_4892)
);

INVx1_ASAP7_75t_L g4893 ( 
.A(n_4700),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4762),
.B(n_4586),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4700),
.Y(n_4895)
);

INVx4_ASAP7_75t_L g4896 ( 
.A(n_4713),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4707),
.Y(n_4897)
);

OAI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4776),
.A2(n_4488),
.B1(n_4480),
.B2(n_4622),
.Y(n_4898)
);

AOI21xp5_ASAP7_75t_L g4899 ( 
.A1(n_4823),
.A2(n_4672),
.B(n_4568),
.Y(n_4899)
);

INVx3_ASAP7_75t_L g4900 ( 
.A(n_4748),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4707),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_L g4902 ( 
.A(n_4733),
.B(n_4586),
.Y(n_4902)
);

OR2x2_ASAP7_75t_L g4903 ( 
.A(n_4739),
.B(n_4543),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4795),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4711),
.Y(n_4905)
);

BUFx2_ASAP7_75t_L g4906 ( 
.A(n_4790),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4711),
.Y(n_4907)
);

NOR2xp33_ASAP7_75t_L g4908 ( 
.A(n_4828),
.B(n_4479),
.Y(n_4908)
);

OR2x6_ASAP7_75t_L g4909 ( 
.A(n_4713),
.B(n_4632),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_SL g4910 ( 
.A1(n_4750),
.A2(n_4685),
.B1(n_4624),
.B2(n_4670),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_L g4911 ( 
.A(n_4765),
.B(n_4586),
.Y(n_4911)
);

BUFx3_ASAP7_75t_L g4912 ( 
.A(n_4726),
.Y(n_4912)
);

INVx2_ASAP7_75t_L g4913 ( 
.A(n_4795),
.Y(n_4913)
);

AOI22xp33_ASAP7_75t_L g4914 ( 
.A1(n_4803),
.A2(n_4607),
.B1(n_4529),
.B2(n_4561),
.Y(n_4914)
);

BUFx5_ASAP7_75t_L g4915 ( 
.A(n_4808),
.Y(n_4915)
);

CKINVDCx20_ASAP7_75t_R g4916 ( 
.A(n_4727),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4748),
.B(n_4602),
.Y(n_4917)
);

AOI21xp5_ASAP7_75t_L g4918 ( 
.A1(n_4827),
.A2(n_4547),
.B(n_4565),
.Y(n_4918)
);

AOI22xp33_ASAP7_75t_L g4919 ( 
.A1(n_4797),
.A2(n_4500),
.B1(n_4668),
.B2(n_4655),
.Y(n_4919)
);

NAND2xp5_ASAP7_75t_L g4920 ( 
.A(n_4782),
.B(n_4602),
.Y(n_4920)
);

AOI22xp33_ASAP7_75t_L g4921 ( 
.A1(n_4743),
.A2(n_4649),
.B1(n_4482),
.B2(n_4691),
.Y(n_4921)
);

CKINVDCx8_ASAP7_75t_R g4922 ( 
.A(n_4720),
.Y(n_4922)
);

OAI222xp33_ASAP7_75t_L g4923 ( 
.A1(n_4874),
.A2(n_4497),
.B1(n_4476),
.B2(n_4585),
.C1(n_4582),
.C2(n_4513),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4728),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4784),
.B(n_4602),
.Y(n_4925)
);

INVxp67_ASAP7_75t_SL g4926 ( 
.A(n_4742),
.Y(n_4926)
);

CKINVDCx5p33_ASAP7_75t_R g4927 ( 
.A(n_4777),
.Y(n_4927)
);

AOI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4743),
.A2(n_4517),
.B1(n_4526),
.B2(n_4487),
.Y(n_4928)
);

OAI22xp33_ASAP7_75t_L g4929 ( 
.A1(n_4776),
.A2(n_4497),
.B1(n_4459),
.B2(n_4563),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4728),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4746),
.Y(n_4931)
);

AOI22xp33_ASAP7_75t_SL g4932 ( 
.A1(n_4841),
.A2(n_4497),
.B1(n_4579),
.B2(n_4459),
.Y(n_4932)
);

OR2x2_ASAP7_75t_L g4933 ( 
.A(n_4746),
.B(n_4543),
.Y(n_4933)
);

NAND3xp33_ASAP7_75t_SL g4934 ( 
.A(n_4781),
.B(n_4662),
.C(n_4650),
.Y(n_4934)
);

AOI22xp33_ASAP7_75t_L g4935 ( 
.A1(n_4767),
.A2(n_4544),
.B1(n_4614),
.B2(n_4459),
.Y(n_4935)
);

AOI22xp33_ASAP7_75t_L g4936 ( 
.A1(n_4834),
.A2(n_4563),
.B1(n_4574),
.B2(n_4567),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_SL g4937 ( 
.A(n_4713),
.B(n_4832),
.Y(n_4937)
);

INVx1_ASAP7_75t_L g4938 ( 
.A(n_4699),
.Y(n_4938)
);

OR2x6_ASAP7_75t_L g4939 ( 
.A(n_4729),
.B(n_4563),
.Y(n_4939)
);

AO31x2_ASAP7_75t_L g4940 ( 
.A1(n_4789),
.A2(n_4684),
.A3(n_4551),
.B(n_4694),
.Y(n_4940)
);

HB1xp67_ASAP7_75t_L g4941 ( 
.A(n_4774),
.Y(n_4941)
);

AOI21xp33_ASAP7_75t_L g4942 ( 
.A1(n_4829),
.A2(n_129),
.B(n_130),
.Y(n_4942)
);

AOI21xp33_ASAP7_75t_L g4943 ( 
.A1(n_4801),
.A2(n_129),
.B(n_130),
.Y(n_4943)
);

AOI221xp5_ASAP7_75t_L g4944 ( 
.A1(n_4811),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.C(n_136),
.Y(n_4944)
);

AOI22xp33_ASAP7_75t_L g4945 ( 
.A1(n_4848),
.A2(n_4510),
.B1(n_4605),
.B2(n_4623),
.Y(n_4945)
);

OR2x2_ASAP7_75t_L g4946 ( 
.A(n_4709),
.B(n_4714),
.Y(n_4946)
);

CKINVDCx14_ASAP7_75t_R g4947 ( 
.A(n_4738),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_4804),
.B(n_4510),
.Y(n_4948)
);

OAI221xp5_ASAP7_75t_L g4949 ( 
.A1(n_4880),
.A2(n_139),
.B1(n_136),
.B2(n_137),
.C(n_140),
.Y(n_4949)
);

INVx2_ASAP7_75t_L g4950 ( 
.A(n_4774),
.Y(n_4950)
);

AND2x2_ASAP7_75t_L g4951 ( 
.A(n_4721),
.B(n_4461),
.Y(n_4951)
);

AND2x4_ASAP7_75t_L g4952 ( 
.A(n_4759),
.B(n_4605),
.Y(n_4952)
);

OR2x2_ASAP7_75t_L g4953 ( 
.A(n_4703),
.B(n_4549),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4716),
.Y(n_4954)
);

OAI22xp33_ASAP7_75t_L g4955 ( 
.A1(n_4832),
.A2(n_4694),
.B1(n_4605),
.B2(n_4549),
.Y(n_4955)
);

AO21x1_ASAP7_75t_L g4956 ( 
.A1(n_4836),
.A2(n_4623),
.B(n_140),
.Y(n_4956)
);

INVx2_ASAP7_75t_L g4957 ( 
.A(n_4800),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4725),
.B(n_4461),
.Y(n_4958)
);

AND2x2_ASAP7_75t_L g4959 ( 
.A(n_4725),
.B(n_4461),
.Y(n_4959)
);

AOI22xp5_ASAP7_75t_L g4960 ( 
.A1(n_4770),
.A2(n_4623),
.B1(n_4549),
.B2(n_144),
.Y(n_4960)
);

OAI22xp5_ASAP7_75t_L g4961 ( 
.A1(n_4831),
.A2(n_4470),
.B1(n_144),
.B2(n_141),
.Y(n_4961)
);

INVx3_ASAP7_75t_L g4962 ( 
.A(n_4740),
.Y(n_4962)
);

BUFx2_ASAP7_75t_L g4963 ( 
.A(n_4740),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4800),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4821),
.A2(n_4470),
.B1(n_145),
.B2(n_141),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4861),
.Y(n_4966)
);

INVx1_ASAP7_75t_L g4967 ( 
.A(n_4861),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4731),
.B(n_4470),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4710),
.B(n_143),
.Y(n_4969)
);

OAI22xp5_ASAP7_75t_L g4970 ( 
.A1(n_4832),
.A2(n_147),
.B1(n_143),
.B2(n_146),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4747),
.Y(n_4971)
);

O2A1O1Ixp33_ASAP7_75t_SL g4972 ( 
.A1(n_4856),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_4972)
);

AOI22xp5_ASAP7_75t_L g4973 ( 
.A1(n_4757),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_4973)
);

AOI22xp33_ASAP7_75t_SL g4974 ( 
.A1(n_4868),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_4974)
);

AOI22xp33_ASAP7_75t_L g4975 ( 
.A1(n_4798),
.A2(n_156),
.B1(n_152),
.B2(n_153),
.Y(n_4975)
);

AND2x4_ASAP7_75t_L g4976 ( 
.A(n_4866),
.B(n_153),
.Y(n_4976)
);

OAI22xp5_ASAP7_75t_L g4977 ( 
.A1(n_4778),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_4977)
);

INVx3_ASAP7_75t_L g4978 ( 
.A(n_4764),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4718),
.Y(n_4979)
);

BUFx3_ASAP7_75t_L g4980 ( 
.A(n_4805),
.Y(n_4980)
);

INVx2_ASAP7_75t_SL g4981 ( 
.A(n_4772),
.Y(n_4981)
);

NAND2xp33_ASAP7_75t_SL g4982 ( 
.A(n_4886),
.B(n_159),
.Y(n_4982)
);

OAI22xp33_ASAP7_75t_L g4983 ( 
.A1(n_4833),
.A2(n_162),
.B1(n_160),
.B2(n_161),
.Y(n_4983)
);

AOI22xp33_ASAP7_75t_L g4984 ( 
.A1(n_4826),
.A2(n_164),
.B1(n_160),
.B2(n_162),
.Y(n_4984)
);

INVx3_ASAP7_75t_L g4985 ( 
.A(n_4840),
.Y(n_4985)
);

AOI21xp5_ASAP7_75t_L g4986 ( 
.A1(n_4867),
.A2(n_611),
.B(n_165),
.Y(n_4986)
);

NOR2xp33_ASAP7_75t_L g4987 ( 
.A(n_4744),
.B(n_166),
.Y(n_4987)
);

OR2x2_ASAP7_75t_L g4988 ( 
.A(n_4863),
.B(n_610),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4865),
.B(n_166),
.Y(n_4989)
);

INVxp67_ASAP7_75t_L g4990 ( 
.A(n_4735),
.Y(n_4990)
);

INVx4_ASAP7_75t_SL g4991 ( 
.A(n_4833),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_4717),
.Y(n_4992)
);

AOI22xp33_ASAP7_75t_SL g4993 ( 
.A1(n_4868),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_4993)
);

AND2x4_ASAP7_75t_L g4994 ( 
.A(n_4860),
.B(n_168),
.Y(n_4994)
);

AND2x4_ASAP7_75t_L g4995 ( 
.A(n_4883),
.B(n_172),
.Y(n_4995)
);

OAI222xp33_ASAP7_75t_L g4996 ( 
.A1(n_4792),
.A2(n_175),
.B1(n_177),
.B2(n_173),
.C1(n_174),
.C2(n_176),
.Y(n_4996)
);

INVx1_ASAP7_75t_L g4997 ( 
.A(n_4863),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4879),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4879),
.Y(n_4999)
);

AOI22xp33_ASAP7_75t_SL g5000 ( 
.A1(n_4871),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4888),
.Y(n_5001)
);

AOI21xp5_ASAP7_75t_L g5002 ( 
.A1(n_4852),
.A2(n_608),
.B(n_176),
.Y(n_5002)
);

HB1xp67_ASAP7_75t_L g5003 ( 
.A(n_4755),
.Y(n_5003)
);

INVx2_ASAP7_75t_L g5004 ( 
.A(n_4717),
.Y(n_5004)
);

AO21x2_ASAP7_75t_L g5005 ( 
.A1(n_4888),
.A2(n_178),
.B(n_179),
.Y(n_5005)
);

HB1xp67_ASAP7_75t_L g5006 ( 
.A(n_4822),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4766),
.B(n_608),
.Y(n_5007)
);

OAI22xp5_ASAP7_75t_L g5008 ( 
.A1(n_4807),
.A2(n_4844),
.B1(n_4719),
.B2(n_4851),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4754),
.B(n_178),
.Y(n_5009)
);

AND2x2_ASAP7_75t_L g5010 ( 
.A(n_4850),
.B(n_180),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4857),
.Y(n_5011)
);

OR2x2_ASAP7_75t_L g5012 ( 
.A(n_4872),
.B(n_181),
.Y(n_5012)
);

HB1xp67_ASAP7_75t_L g5013 ( 
.A(n_4808),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_4812),
.Y(n_5014)
);

NAND3xp33_ASAP7_75t_L g5015 ( 
.A(n_4780),
.B(n_183),
.C(n_186),
.Y(n_5015)
);

NAND2x1_ASAP7_75t_L g5016 ( 
.A(n_4771),
.B(n_183),
.Y(n_5016)
);

AND2x2_ASAP7_75t_SL g5017 ( 
.A(n_4890),
.B(n_186),
.Y(n_5017)
);

NAND2x1p5_ASAP7_75t_L g5018 ( 
.A(n_4890),
.B(n_188),
.Y(n_5018)
);

CKINVDCx5p33_ASAP7_75t_R g5019 ( 
.A(n_4724),
.Y(n_5019)
);

AO21x1_ASAP7_75t_L g5020 ( 
.A1(n_4812),
.A2(n_190),
.B(n_191),
.Y(n_5020)
);

INVx2_ASAP7_75t_L g5021 ( 
.A(n_4702),
.Y(n_5021)
);

BUFx3_ASAP7_75t_L g5022 ( 
.A(n_4760),
.Y(n_5022)
);

NOR2xp33_ASAP7_75t_L g5023 ( 
.A(n_4871),
.B(n_193),
.Y(n_5023)
);

AO31x2_ASAP7_75t_L g5024 ( 
.A1(n_4837),
.A2(n_196),
.A3(n_193),
.B(n_195),
.Y(n_5024)
);

OAI21x1_ASAP7_75t_L g5025 ( 
.A1(n_4705),
.A2(n_195),
.B(n_197),
.Y(n_5025)
);

AOI22xp33_ASAP7_75t_L g5026 ( 
.A1(n_4882),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.Y(n_5026)
);

HB1xp67_ASAP7_75t_L g5027 ( 
.A(n_4819),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4885),
.Y(n_5028)
);

BUFx5_ASAP7_75t_L g5029 ( 
.A(n_4837),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4817),
.B(n_607),
.Y(n_5030)
);

OAI21x1_ASAP7_75t_L g5031 ( 
.A1(n_4708),
.A2(n_198),
.B(n_200),
.Y(n_5031)
);

INVx2_ASAP7_75t_L g5032 ( 
.A(n_4818),
.Y(n_5032)
);

OAI21x1_ASAP7_75t_L g5033 ( 
.A1(n_4706),
.A2(n_201),
.B(n_202),
.Y(n_5033)
);

OAI21xp5_ASAP7_75t_L g5034 ( 
.A1(n_4779),
.A2(n_201),
.B(n_205),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_4840),
.Y(n_5035)
);

HB1xp67_ASAP7_75t_L g5036 ( 
.A(n_4737),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4758),
.A2(n_208),
.B(n_210),
.Y(n_5037)
);

INVx4_ASAP7_75t_L g5038 ( 
.A(n_4704),
.Y(n_5038)
);

OAI221xp5_ASAP7_75t_L g5039 ( 
.A1(n_4761),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.C(n_212),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4842),
.B(n_607),
.Y(n_5040)
);

AND2x2_ASAP7_75t_L g5041 ( 
.A(n_4906),
.B(n_4704),
.Y(n_5041)
);

AND2x4_ASAP7_75t_L g5042 ( 
.A(n_4952),
.B(n_4937),
.Y(n_5042)
);

AND2x2_ASAP7_75t_L g5043 ( 
.A(n_4900),
.B(n_4869),
.Y(n_5043)
);

AOI221xp5_ASAP7_75t_L g5044 ( 
.A1(n_4923),
.A2(n_4825),
.B1(n_4745),
.B2(n_4887),
.C(n_4753),
.Y(n_5044)
);

BUFx3_ASAP7_75t_L g5045 ( 
.A(n_4912),
.Y(n_5045)
);

AOI21xp33_ASAP7_75t_L g5046 ( 
.A1(n_4932),
.A2(n_4824),
.B(n_4758),
.Y(n_5046)
);

BUFx6f_ASAP7_75t_L g5047 ( 
.A(n_4896),
.Y(n_5047)
);

AND2x2_ASAP7_75t_L g5048 ( 
.A(n_4900),
.B(n_4869),
.Y(n_5048)
);

OAI22xp5_ASAP7_75t_SL g5049 ( 
.A1(n_4922),
.A2(n_4947),
.B1(n_5038),
.B2(n_4896),
.Y(n_5049)
);

BUFx5_ASAP7_75t_L g5050 ( 
.A(n_5028),
.Y(n_5050)
);

OR2x2_ASAP7_75t_L g5051 ( 
.A(n_4892),
.B(n_4894),
.Y(n_5051)
);

AO21x2_ASAP7_75t_L g5052 ( 
.A1(n_4992),
.A2(n_4859),
.B(n_4858),
.Y(n_5052)
);

OAI22xp5_ASAP7_75t_L g5053 ( 
.A1(n_4975),
.A2(n_4883),
.B1(n_4884),
.B2(n_4712),
.Y(n_5053)
);

OAI22xp5_ASAP7_75t_L g5054 ( 
.A1(n_4936),
.A2(n_4771),
.B1(n_4839),
.B2(n_4843),
.Y(n_5054)
);

AOI21xp5_ASAP7_75t_L g5055 ( 
.A1(n_4918),
.A2(n_4756),
.B(n_4736),
.Y(n_5055)
);

AOI21xp33_ASAP7_75t_L g5056 ( 
.A1(n_5008),
.A2(n_4802),
.B(n_4806),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4893),
.Y(n_5057)
);

INVx1_ASAP7_75t_L g5058 ( 
.A(n_4895),
.Y(n_5058)
);

AOI21xp5_ASAP7_75t_L g5059 ( 
.A1(n_4899),
.A2(n_4796),
.B(n_4768),
.Y(n_5059)
);

AO31x2_ASAP7_75t_L g5060 ( 
.A1(n_5020),
.A2(n_4858),
.A3(n_4859),
.B(n_4741),
.Y(n_5060)
);

AOI22xp33_ASAP7_75t_L g5061 ( 
.A1(n_4934),
.A2(n_4891),
.B1(n_4855),
.B2(n_4701),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_4897),
.Y(n_5062)
);

INVx5_ASAP7_75t_L g5063 ( 
.A(n_5038),
.Y(n_5063)
);

NOR2x1_ASAP7_75t_L g5064 ( 
.A(n_4978),
.B(n_4839),
.Y(n_5064)
);

HB1xp67_ASAP7_75t_L g5065 ( 
.A(n_4941),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_4901),
.Y(n_5066)
);

OAI22xp5_ASAP7_75t_L g5067 ( 
.A1(n_4910),
.A2(n_4843),
.B1(n_4814),
.B2(n_4820),
.Y(n_5067)
);

AOI22xp33_ASAP7_75t_L g5068 ( 
.A1(n_4943),
.A2(n_4878),
.B1(n_4875),
.B2(n_4835),
.Y(n_5068)
);

AOI22xp33_ASAP7_75t_SL g5069 ( 
.A1(n_5017),
.A2(n_4877),
.B1(n_4820),
.B2(n_4847),
.Y(n_5069)
);

NOR2xp33_ASAP7_75t_SL g5070 ( 
.A(n_4927),
.B(n_4734),
.Y(n_5070)
);

AND2x2_ASAP7_75t_L g5071 ( 
.A(n_4963),
.B(n_4715),
.Y(n_5071)
);

AOI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4929),
.A2(n_4986),
.B(n_4898),
.Y(n_5072)
);

NOR2xp33_ASAP7_75t_L g5073 ( 
.A(n_4990),
.B(n_4813),
.Y(n_5073)
);

AOI221xp5_ASAP7_75t_L g5074 ( 
.A1(n_4942),
.A2(n_4813),
.B1(n_4846),
.B2(n_4830),
.C(n_4791),
.Y(n_5074)
);

AO22x2_ASAP7_75t_L g5075 ( 
.A1(n_5004),
.A2(n_4847),
.B1(n_4799),
.B2(n_4741),
.Y(n_5075)
);

INVx4_ASAP7_75t_SL g5076 ( 
.A(n_4980),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4911),
.B(n_4938),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4905),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4962),
.B(n_4715),
.Y(n_5079)
);

AOI22xp33_ASAP7_75t_L g5080 ( 
.A1(n_5015),
.A2(n_4751),
.B1(n_4799),
.B2(n_4854),
.Y(n_5080)
);

BUFx10_ASAP7_75t_L g5081 ( 
.A(n_5023),
.Y(n_5081)
);

NAND2xp5_ASAP7_75t_L g5082 ( 
.A(n_4954),
.B(n_4741),
.Y(n_5082)
);

OR2x6_ASAP7_75t_L g5083 ( 
.A(n_4909),
.B(n_4730),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_L g5084 ( 
.A(n_4902),
.B(n_4737),
.Y(n_5084)
);

OAI211xp5_ASAP7_75t_SL g5085 ( 
.A1(n_4914),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4907),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_5032),
.B(n_4737),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4964),
.B(n_4773),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4924),
.Y(n_5089)
);

OR2x6_ASAP7_75t_L g5090 ( 
.A(n_4909),
.B(n_4715),
.Y(n_5090)
);

OAI22xp5_ASAP7_75t_L g5091 ( 
.A1(n_4935),
.A2(n_4873),
.B1(n_4749),
.B2(n_4773),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4930),
.Y(n_5092)
);

AOI22xp33_ASAP7_75t_L g5093 ( 
.A1(n_4956),
.A2(n_4864),
.B1(n_4862),
.B2(n_4815),
.Y(n_5093)
);

AOI22xp33_ASAP7_75t_SL g5094 ( 
.A1(n_4949),
.A2(n_4845),
.B1(n_4853),
.B2(n_4870),
.Y(n_5094)
);

AO21x2_ASAP7_75t_L g5095 ( 
.A1(n_4926),
.A2(n_4838),
.B(n_4794),
.Y(n_5095)
);

AOI22xp33_ASAP7_75t_L g5096 ( 
.A1(n_5039),
.A2(n_4752),
.B1(n_4732),
.B2(n_4783),
.Y(n_5096)
);

NOR2xp33_ASAP7_75t_L g5097 ( 
.A(n_4916),
.B(n_5019),
.Y(n_5097)
);

AOI22xp33_ASAP7_75t_L g5098 ( 
.A1(n_4984),
.A2(n_4849),
.B1(n_4881),
.B2(n_4889),
.Y(n_5098)
);

AOI22xp33_ASAP7_75t_L g5099 ( 
.A1(n_4965),
.A2(n_4793),
.B1(n_4722),
.B2(n_4809),
.Y(n_5099)
);

AOI221xp5_ASAP7_75t_L g5100 ( 
.A1(n_4983),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.C(n_218),
.Y(n_5100)
);

AOI22xp33_ASAP7_75t_L g5101 ( 
.A1(n_4919),
.A2(n_4810),
.B1(n_4816),
.B2(n_4786),
.Y(n_5101)
);

OAI21x1_ASAP7_75t_L g5102 ( 
.A1(n_5021),
.A2(n_4723),
.B(n_4769),
.Y(n_5102)
);

AOI22xp5_ASAP7_75t_L g5103 ( 
.A1(n_4977),
.A2(n_4788),
.B1(n_4787),
.B2(n_4763),
.Y(n_5103)
);

INVx1_ASAP7_75t_L g5104 ( 
.A(n_5011),
.Y(n_5104)
);

OAI22xp5_ASAP7_75t_L g5105 ( 
.A1(n_4974),
.A2(n_4993),
.B1(n_4928),
.B2(n_4960),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_4917),
.B(n_4773),
.Y(n_5106)
);

OR2x2_ASAP7_75t_L g5107 ( 
.A(n_4946),
.B(n_4749),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_4966),
.Y(n_5108)
);

AOI22xp33_ASAP7_75t_L g5109 ( 
.A1(n_5037),
.A2(n_4749),
.B1(n_4876),
.B2(n_4785),
.Y(n_5109)
);

O2A1O1Ixp5_ASAP7_75t_L g5110 ( 
.A1(n_5016),
.A2(n_4785),
.B(n_4876),
.C(n_222),
.Y(n_5110)
);

AND2x4_ASAP7_75t_L g5111 ( 
.A(n_4952),
.B(n_4785),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4967),
.Y(n_5112)
);

CKINVDCx11_ASAP7_75t_R g5113 ( 
.A(n_4991),
.Y(n_5113)
);

INVxp67_ASAP7_75t_L g5114 ( 
.A(n_4908),
.Y(n_5114)
);

AOI221xp5_ASAP7_75t_L g5115 ( 
.A1(n_4972),
.A2(n_4996),
.B1(n_4944),
.B2(n_4970),
.C(n_5034),
.Y(n_5115)
);

INVx2_ASAP7_75t_L g5116 ( 
.A(n_4957),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_4904),
.Y(n_5117)
);

INVxp67_ASAP7_75t_SL g5118 ( 
.A(n_5036),
.Y(n_5118)
);

OAI221xp5_ASAP7_75t_L g5119 ( 
.A1(n_4973),
.A2(n_222),
.B1(n_219),
.B2(n_220),
.C(n_223),
.Y(n_5119)
);

OR2x2_ASAP7_75t_L g5120 ( 
.A(n_4920),
.B(n_4925),
.Y(n_5120)
);

BUFx4f_ASAP7_75t_L g5121 ( 
.A(n_5010),
.Y(n_5121)
);

AND2x2_ASAP7_75t_L g5122 ( 
.A(n_4962),
.B(n_4876),
.Y(n_5122)
);

OAI211xp5_ASAP7_75t_L g5123 ( 
.A1(n_5000),
.A2(n_226),
.B(n_220),
.C(n_225),
.Y(n_5123)
);

AND2x2_ASAP7_75t_L g5124 ( 
.A(n_4978),
.B(n_227),
.Y(n_5124)
);

NOR2xp33_ASAP7_75t_L g5125 ( 
.A(n_4989),
.B(n_5030),
.Y(n_5125)
);

INVx2_ASAP7_75t_L g5126 ( 
.A(n_4913),
.Y(n_5126)
);

BUFx3_ASAP7_75t_L g5127 ( 
.A(n_5022),
.Y(n_5127)
);

INVx2_ASAP7_75t_L g5128 ( 
.A(n_4931),
.Y(n_5128)
);

AOI221xp5_ASAP7_75t_L g5129 ( 
.A1(n_5002),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_5129)
);

BUFx2_ASAP7_75t_L g5130 ( 
.A(n_4985),
.Y(n_5130)
);

AOI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_4961),
.A2(n_228),
.B(n_230),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_4997),
.Y(n_5132)
);

AOI22xp33_ASAP7_75t_L g5133 ( 
.A1(n_4939),
.A2(n_235),
.B1(n_231),
.B2(n_232),
.Y(n_5133)
);

NAND3xp33_ASAP7_75t_L g5134 ( 
.A(n_5026),
.B(n_235),
.C(n_236),
.Y(n_5134)
);

OR2x2_ASAP7_75t_SL g5135 ( 
.A(n_4979),
.B(n_236),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_4998),
.Y(n_5136)
);

BUFx12f_ASAP7_75t_L g5137 ( 
.A(n_4994),
.Y(n_5137)
);

AOI22xp33_ASAP7_75t_L g5138 ( 
.A1(n_4939),
.A2(n_241),
.B1(n_238),
.B2(n_240),
.Y(n_5138)
);

INVx3_ASAP7_75t_L g5139 ( 
.A(n_4985),
.Y(n_5139)
);

AOI22xp33_ASAP7_75t_L g5140 ( 
.A1(n_4982),
.A2(n_244),
.B1(n_241),
.B2(n_242),
.Y(n_5140)
);

OR2x2_ASAP7_75t_L g5141 ( 
.A(n_4903),
.B(n_605),
.Y(n_5141)
);

AO21x2_ASAP7_75t_L g5142 ( 
.A1(n_5003),
.A2(n_242),
.B(n_244),
.Y(n_5142)
);

AND2x4_ASAP7_75t_L g5143 ( 
.A(n_4958),
.B(n_246),
.Y(n_5143)
);

OAI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_4921),
.A2(n_249),
.B1(n_246),
.B2(n_248),
.Y(n_5144)
);

OAI21xp33_ASAP7_75t_SL g5145 ( 
.A1(n_5025),
.A2(n_248),
.B(n_249),
.Y(n_5145)
);

AO21x2_ASAP7_75t_L g5146 ( 
.A1(n_4999),
.A2(n_250),
.B(n_252),
.Y(n_5146)
);

AOI221xp5_ASAP7_75t_L g5147 ( 
.A1(n_4969),
.A2(n_255),
.B1(n_252),
.B2(n_254),
.C(n_257),
.Y(n_5147)
);

OAI22xp33_ASAP7_75t_L g5148 ( 
.A1(n_4988),
.A2(n_261),
.B1(n_257),
.B2(n_259),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_4950),
.B(n_4951),
.Y(n_5149)
);

A2O1A1Ixp33_ASAP7_75t_L g5150 ( 
.A1(n_4987),
.A2(n_262),
.B(n_259),
.C(n_261),
.Y(n_5150)
);

CKINVDCx5p33_ASAP7_75t_R g5151 ( 
.A(n_4981),
.Y(n_5151)
);

AOI221x1_ASAP7_75t_SL g5152 ( 
.A1(n_5009),
.A2(n_265),
.B1(n_262),
.B2(n_264),
.C(n_266),
.Y(n_5152)
);

AO21x2_ASAP7_75t_L g5153 ( 
.A1(n_5001),
.A2(n_264),
.B(n_266),
.Y(n_5153)
);

AOI21xp5_ASAP7_75t_L g5154 ( 
.A1(n_4955),
.A2(n_267),
.B(n_268),
.Y(n_5154)
);

OAI22xp33_ASAP7_75t_L g5155 ( 
.A1(n_5012),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_5155)
);

OAI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_5031),
.A2(n_269),
.B(n_270),
.Y(n_5156)
);

OAI21x1_ASAP7_75t_L g5157 ( 
.A1(n_4933),
.A2(n_270),
.B(n_271),
.Y(n_5157)
);

AOI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4945),
.A2(n_271),
.B(n_272),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_5035),
.B(n_272),
.Y(n_5159)
);

AOI22xp33_ASAP7_75t_SL g5160 ( 
.A1(n_5005),
.A2(n_276),
.B1(n_273),
.B2(n_275),
.Y(n_5160)
);

AOI21xp5_ASAP7_75t_L g5161 ( 
.A1(n_4948),
.A2(n_604),
.B(n_273),
.Y(n_5161)
);

OAI221xp5_ASAP7_75t_L g5162 ( 
.A1(n_5018),
.A2(n_603),
.B1(n_278),
.B2(n_275),
.C(n_277),
.Y(n_5162)
);

OAI221xp5_ASAP7_75t_L g5163 ( 
.A1(n_5007),
.A2(n_5040),
.B1(n_4968),
.B2(n_4953),
.C(n_5006),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_5013),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5014),
.Y(n_5165)
);

OR2x6_ASAP7_75t_L g5166 ( 
.A(n_4995),
.B(n_279),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_5027),
.Y(n_5167)
);

INVxp67_ASAP7_75t_L g5168 ( 
.A(n_4976),
.Y(n_5168)
);

INVx2_ASAP7_75t_L g5169 ( 
.A(n_4915),
.Y(n_5169)
);

AOI21xp5_ASAP7_75t_L g5170 ( 
.A1(n_5033),
.A2(n_602),
.B(n_279),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_4971),
.Y(n_5171)
);

OAI22xp5_ASAP7_75t_L g5172 ( 
.A1(n_4995),
.A2(n_283),
.B1(n_280),
.B2(n_282),
.Y(n_5172)
);

AOI21xp5_ASAP7_75t_L g5173 ( 
.A1(n_4976),
.A2(n_280),
.B(n_283),
.Y(n_5173)
);

INVx2_ASAP7_75t_L g5174 ( 
.A(n_4915),
.Y(n_5174)
);

AOI22xp33_ASAP7_75t_L g5175 ( 
.A1(n_4991),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4959),
.B(n_4940),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4915),
.Y(n_5177)
);

OAI21x1_ASAP7_75t_L g5178 ( 
.A1(n_4915),
.A2(n_285),
.B(n_286),
.Y(n_5178)
);

AND2x4_ASAP7_75t_L g5179 ( 
.A(n_4994),
.B(n_287),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_4915),
.Y(n_5180)
);

OAI211xp5_ASAP7_75t_L g5181 ( 
.A1(n_4940),
.A2(n_291),
.B(n_287),
.C(n_290),
.Y(n_5181)
);

OAI221xp5_ASAP7_75t_L g5182 ( 
.A1(n_4940),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.C(n_293),
.Y(n_5182)
);

NAND2xp5_ASAP7_75t_L g5183 ( 
.A(n_5114),
.B(n_5024),
.Y(n_5183)
);

NAND2xp33_ASAP7_75t_R g5184 ( 
.A(n_5166),
.B(n_292),
.Y(n_5184)
);

INVx2_ASAP7_75t_L g5185 ( 
.A(n_5050),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_5050),
.Y(n_5186)
);

NOR2xp33_ASAP7_75t_R g5187 ( 
.A(n_5113),
.B(n_293),
.Y(n_5187)
);

INVx2_ASAP7_75t_L g5188 ( 
.A(n_5050),
.Y(n_5188)
);

BUFx3_ASAP7_75t_L g5189 ( 
.A(n_5137),
.Y(n_5189)
);

INVxp67_ASAP7_75t_L g5190 ( 
.A(n_5141),
.Y(n_5190)
);

OR2x6_ASAP7_75t_L g5191 ( 
.A(n_5049),
.B(n_5024),
.Y(n_5191)
);

NAND2xp33_ASAP7_75t_R g5192 ( 
.A(n_5166),
.B(n_294),
.Y(n_5192)
);

INVx1_ASAP7_75t_L g5193 ( 
.A(n_5057),
.Y(n_5193)
);

XOR2xp5_ASAP7_75t_L g5194 ( 
.A(n_5151),
.B(n_294),
.Y(n_5194)
);

INVxp67_ASAP7_75t_L g5195 ( 
.A(n_5142),
.Y(n_5195)
);

NAND2xp33_ASAP7_75t_R g5196 ( 
.A(n_5179),
.B(n_295),
.Y(n_5196)
);

XNOR2xp5_ASAP7_75t_L g5197 ( 
.A(n_5135),
.B(n_297),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_5072),
.B(n_5024),
.Y(n_5198)
);

BUFx2_ASAP7_75t_L g5199 ( 
.A(n_5090),
.Y(n_5199)
);

INVxp67_ASAP7_75t_L g5200 ( 
.A(n_5163),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_R g5201 ( 
.A(n_5070),
.B(n_297),
.Y(n_5201)
);

NAND2xp33_ASAP7_75t_SL g5202 ( 
.A(n_5041),
.B(n_298),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_5125),
.B(n_5029),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_5056),
.B(n_5029),
.Y(n_5204)
);

OR2x6_ASAP7_75t_L g5205 ( 
.A(n_5090),
.B(n_5029),
.Y(n_5205)
);

AND2x2_ASAP7_75t_L g5206 ( 
.A(n_5043),
.B(n_5029),
.Y(n_5206)
);

INVxp67_ASAP7_75t_L g5207 ( 
.A(n_5075),
.Y(n_5207)
);

NOR2xp33_ASAP7_75t_R g5208 ( 
.A(n_5081),
.B(n_298),
.Y(n_5208)
);

OR2x6_ASAP7_75t_L g5209 ( 
.A(n_5047),
.B(n_5029),
.Y(n_5209)
);

NOR2xp33_ASAP7_75t_L g5210 ( 
.A(n_5045),
.B(n_299),
.Y(n_5210)
);

NAND2xp33_ASAP7_75t_SL g5211 ( 
.A(n_5047),
.B(n_299),
.Y(n_5211)
);

AND2x2_ASAP7_75t_L g5212 ( 
.A(n_5048),
.B(n_300),
.Y(n_5212)
);

AND2x2_ASAP7_75t_SL g5213 ( 
.A(n_5121),
.B(n_5061),
.Y(n_5213)
);

AND2x2_ASAP7_75t_L g5214 ( 
.A(n_5042),
.B(n_301),
.Y(n_5214)
);

OR2x6_ASAP7_75t_L g5215 ( 
.A(n_5047),
.B(n_5055),
.Y(n_5215)
);

INVx2_ASAP7_75t_L g5216 ( 
.A(n_5050),
.Y(n_5216)
);

NAND2xp33_ASAP7_75t_R g5217 ( 
.A(n_5179),
.B(n_601),
.Y(n_5217)
);

AND2x4_ASAP7_75t_L g5218 ( 
.A(n_5042),
.B(n_303),
.Y(n_5218)
);

NAND2xp5_ASAP7_75t_L g5219 ( 
.A(n_5046),
.B(n_303),
.Y(n_5219)
);

OR2x6_ASAP7_75t_L g5220 ( 
.A(n_5083),
.B(n_304),
.Y(n_5220)
);

NAND2xp5_ASAP7_75t_SL g5221 ( 
.A(n_5067),
.B(n_305),
.Y(n_5221)
);

AND2x2_ASAP7_75t_L g5222 ( 
.A(n_5071),
.B(n_307),
.Y(n_5222)
);

CKINVDCx11_ASAP7_75t_R g5223 ( 
.A(n_5076),
.Y(n_5223)
);

AND2x2_ASAP7_75t_L g5224 ( 
.A(n_5079),
.B(n_309),
.Y(n_5224)
);

INVx1_ASAP7_75t_L g5225 ( 
.A(n_5058),
.Y(n_5225)
);

INVxp67_ASAP7_75t_L g5226 ( 
.A(n_5075),
.Y(n_5226)
);

NAND2xp5_ASAP7_75t_L g5227 ( 
.A(n_5168),
.B(n_311),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_5106),
.B(n_311),
.Y(n_5228)
);

NAND2xp33_ASAP7_75t_SL g5229 ( 
.A(n_5105),
.B(n_312),
.Y(n_5229)
);

BUFx6f_ASAP7_75t_L g5230 ( 
.A(n_5063),
.Y(n_5230)
);

CKINVDCx8_ASAP7_75t_R g5231 ( 
.A(n_5076),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_5159),
.B(n_313),
.Y(n_5232)
);

NAND2xp33_ASAP7_75t_R g5233 ( 
.A(n_5143),
.B(n_314),
.Y(n_5233)
);

XNOR2xp5_ASAP7_75t_L g5234 ( 
.A(n_5127),
.B(n_315),
.Y(n_5234)
);

NOR2xp33_ASAP7_75t_R g5235 ( 
.A(n_5081),
.B(n_315),
.Y(n_5235)
);

XNOR2xp5_ASAP7_75t_L g5236 ( 
.A(n_5152),
.B(n_317),
.Y(n_5236)
);

INVxp67_ASAP7_75t_L g5237 ( 
.A(n_5073),
.Y(n_5237)
);

CKINVDCx5p33_ASAP7_75t_R g5238 ( 
.A(n_5097),
.Y(n_5238)
);

NAND2x1p5_ASAP7_75t_L g5239 ( 
.A(n_5063),
.B(n_317),
.Y(n_5239)
);

INVx2_ASAP7_75t_L g5240 ( 
.A(n_5130),
.Y(n_5240)
);

NOR2xp33_ASAP7_75t_L g5241 ( 
.A(n_5063),
.B(n_318),
.Y(n_5241)
);

INVx2_ASAP7_75t_L g5242 ( 
.A(n_5139),
.Y(n_5242)
);

AND2x2_ASAP7_75t_L g5243 ( 
.A(n_5143),
.B(n_318),
.Y(n_5243)
);

NAND2xp33_ASAP7_75t_R g5244 ( 
.A(n_5083),
.B(n_319),
.Y(n_5244)
);

AND2x4_ASAP7_75t_L g5245 ( 
.A(n_5167),
.B(n_319),
.Y(n_5245)
);

OR2x6_ASAP7_75t_L g5246 ( 
.A(n_5154),
.B(n_320),
.Y(n_5246)
);

NAND2xp5_ASAP7_75t_L g5247 ( 
.A(n_5161),
.B(n_321),
.Y(n_5247)
);

NAND2xp33_ASAP7_75t_SL g5248 ( 
.A(n_5124),
.B(n_5146),
.Y(n_5248)
);

BUFx3_ASAP7_75t_L g5249 ( 
.A(n_5065),
.Y(n_5249)
);

AND2x2_ASAP7_75t_L g5250 ( 
.A(n_5149),
.B(n_324),
.Y(n_5250)
);

NAND2xp33_ASAP7_75t_R g5251 ( 
.A(n_5156),
.B(n_599),
.Y(n_5251)
);

NAND2xp33_ASAP7_75t_R g5252 ( 
.A(n_5173),
.B(n_599),
.Y(n_5252)
);

AND2x4_ASAP7_75t_L g5253 ( 
.A(n_5164),
.B(n_324),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_5062),
.Y(n_5254)
);

XNOR2xp5_ASAP7_75t_L g5255 ( 
.A(n_5069),
.B(n_325),
.Y(n_5255)
);

NAND2xp33_ASAP7_75t_R g5256 ( 
.A(n_5157),
.B(n_598),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_5172),
.Y(n_5257)
);

CKINVDCx11_ASAP7_75t_R g5258 ( 
.A(n_5053),
.Y(n_5258)
);

OR2x6_ASAP7_75t_L g5259 ( 
.A(n_5059),
.B(n_325),
.Y(n_5259)
);

CKINVDCx20_ASAP7_75t_R g5260 ( 
.A(n_5144),
.Y(n_5260)
);

AND2x4_ASAP7_75t_L g5261 ( 
.A(n_5111),
.B(n_326),
.Y(n_5261)
);

NAND2xp33_ASAP7_75t_SL g5262 ( 
.A(n_5153),
.B(n_327),
.Y(n_5262)
);

NOR2xp33_ASAP7_75t_R g5263 ( 
.A(n_5175),
.B(n_327),
.Y(n_5263)
);

NAND2xp33_ASAP7_75t_SL g5264 ( 
.A(n_5133),
.B(n_328),
.Y(n_5264)
);

NAND2xp33_ASAP7_75t_R g5265 ( 
.A(n_5178),
.B(n_597),
.Y(n_5265)
);

AND2x2_ASAP7_75t_L g5266 ( 
.A(n_5051),
.B(n_328),
.Y(n_5266)
);

NOR2xp33_ASAP7_75t_R g5267 ( 
.A(n_5140),
.B(n_329),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_5077),
.B(n_329),
.Y(n_5268)
);

NAND2xp33_ASAP7_75t_R g5269 ( 
.A(n_5158),
.B(n_5170),
.Y(n_5269)
);

NAND2xp33_ASAP7_75t_R g5270 ( 
.A(n_5131),
.B(n_597),
.Y(n_5270)
);

INVx1_ASAP7_75t_L g5271 ( 
.A(n_5066),
.Y(n_5271)
);

NOR2xp33_ASAP7_75t_R g5272 ( 
.A(n_5138),
.B(n_5080),
.Y(n_5272)
);

AND2x4_ASAP7_75t_L g5273 ( 
.A(n_5111),
.B(n_330),
.Y(n_5273)
);

NOR2xp33_ASAP7_75t_R g5274 ( 
.A(n_5068),
.B(n_330),
.Y(n_5274)
);

NAND2xp33_ASAP7_75t_R g5275 ( 
.A(n_5107),
.B(n_596),
.Y(n_5275)
);

NAND2xp33_ASAP7_75t_R g5276 ( 
.A(n_5082),
.B(n_331),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_5078),
.Y(n_5277)
);

NAND2xp33_ASAP7_75t_SL g5278 ( 
.A(n_5054),
.B(n_331),
.Y(n_5278)
);

NAND2xp5_ASAP7_75t_L g5279 ( 
.A(n_5084),
.B(n_332),
.Y(n_5279)
);

NAND2xp33_ASAP7_75t_R g5280 ( 
.A(n_5088),
.B(n_333),
.Y(n_5280)
);

INVx1_ASAP7_75t_L g5281 ( 
.A(n_5086),
.Y(n_5281)
);

CKINVDCx8_ASAP7_75t_R g5282 ( 
.A(n_5123),
.Y(n_5282)
);

NOR2xp33_ASAP7_75t_R g5283 ( 
.A(n_5098),
.B(n_333),
.Y(n_5283)
);

NAND2xp33_ASAP7_75t_SL g5284 ( 
.A(n_5091),
.B(n_334),
.Y(n_5284)
);

NAND2xp33_ASAP7_75t_R g5285 ( 
.A(n_5087),
.B(n_595),
.Y(n_5285)
);

INVx1_ASAP7_75t_L g5286 ( 
.A(n_5089),
.Y(n_5286)
);

NAND2xp33_ASAP7_75t_R g5287 ( 
.A(n_5176),
.B(n_595),
.Y(n_5287)
);

CKINVDCx12_ASAP7_75t_R g5288 ( 
.A(n_5120),
.Y(n_5288)
);

NAND2xp33_ASAP7_75t_R g5289 ( 
.A(n_5122),
.B(n_334),
.Y(n_5289)
);

NAND2xp33_ASAP7_75t_R g5290 ( 
.A(n_5115),
.B(n_594),
.Y(n_5290)
);

INVx1_ASAP7_75t_L g5291 ( 
.A(n_5092),
.Y(n_5291)
);

NAND2xp33_ASAP7_75t_SL g5292 ( 
.A(n_5085),
.B(n_335),
.Y(n_5292)
);

BUFx3_ASAP7_75t_L g5293 ( 
.A(n_5104),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5193),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5198),
.B(n_5074),
.Y(n_5295)
);

AND2x2_ASAP7_75t_L g5296 ( 
.A(n_5199),
.B(n_5118),
.Y(n_5296)
);

AND2x2_ASAP7_75t_L g5297 ( 
.A(n_5215),
.B(n_5064),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_5249),
.Y(n_5298)
);

AND2x2_ASAP7_75t_L g5299 ( 
.A(n_5215),
.B(n_5128),
.Y(n_5299)
);

AND2x4_ASAP7_75t_L g5300 ( 
.A(n_5230),
.B(n_5240),
.Y(n_5300)
);

INVx1_ASAP7_75t_L g5301 ( 
.A(n_5225),
.Y(n_5301)
);

BUFx3_ASAP7_75t_L g5302 ( 
.A(n_5223),
.Y(n_5302)
);

AND2x4_ASAP7_75t_SL g5303 ( 
.A(n_5218),
.B(n_5101),
.Y(n_5303)
);

INVx2_ASAP7_75t_R g5304 ( 
.A(n_5275),
.Y(n_5304)
);

INVx5_ASAP7_75t_L g5305 ( 
.A(n_5230),
.Y(n_5305)
);

AND2x2_ASAP7_75t_L g5306 ( 
.A(n_5205),
.B(n_5117),
.Y(n_5306)
);

INVx1_ASAP7_75t_L g5307 ( 
.A(n_5254),
.Y(n_5307)
);

OAI22xp33_ASAP7_75t_L g5308 ( 
.A1(n_5280),
.A2(n_5182),
.B1(n_5103),
.B2(n_5119),
.Y(n_5308)
);

NOR2xp33_ASAP7_75t_L g5309 ( 
.A(n_5231),
.B(n_5150),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5271),
.Y(n_5310)
);

OAI21xp5_ASAP7_75t_SL g5311 ( 
.A1(n_5221),
.A2(n_5044),
.B(n_5134),
.Y(n_5311)
);

AND2x4_ASAP7_75t_L g5312 ( 
.A(n_5230),
.B(n_5169),
.Y(n_5312)
);

HB1xp67_ASAP7_75t_L g5313 ( 
.A(n_5288),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5277),
.Y(n_5314)
);

INVx2_ASAP7_75t_L g5315 ( 
.A(n_5261),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_5281),
.Y(n_5316)
);

INVx3_ASAP7_75t_L g5317 ( 
.A(n_5205),
.Y(n_5317)
);

INVx2_ASAP7_75t_L g5318 ( 
.A(n_5261),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_5286),
.Y(n_5319)
);

OA21x2_ASAP7_75t_L g5320 ( 
.A1(n_5195),
.A2(n_5180),
.B(n_5177),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_5200),
.B(n_5190),
.Y(n_5321)
);

BUFx2_ASAP7_75t_L g5322 ( 
.A(n_5220),
.Y(n_5322)
);

NAND2xp5_ASAP7_75t_L g5323 ( 
.A(n_5237),
.B(n_5094),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_5191),
.B(n_5242),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5291),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5279),
.B(n_5148),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_5293),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5273),
.Y(n_5328)
);

AO31x2_ASAP7_75t_L g5329 ( 
.A1(n_5183),
.A2(n_5174),
.A3(n_5112),
.B(n_5132),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5273),
.Y(n_5330)
);

AND2x2_ASAP7_75t_L g5331 ( 
.A(n_5191),
.B(n_5126),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_5228),
.B(n_5155),
.Y(n_5332)
);

INVx2_ASAP7_75t_L g5333 ( 
.A(n_5218),
.Y(n_5333)
);

AND2x2_ASAP7_75t_L g5334 ( 
.A(n_5220),
.B(n_5116),
.Y(n_5334)
);

INVx3_ASAP7_75t_L g5335 ( 
.A(n_5209),
.Y(n_5335)
);

OAI221xp5_ASAP7_75t_L g5336 ( 
.A1(n_5290),
.A2(n_5129),
.B1(n_5147),
.B2(n_5160),
.C(n_5100),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_L g5337 ( 
.A(n_5253),
.B(n_5266),
.Y(n_5337)
);

HB1xp67_ASAP7_75t_L g5338 ( 
.A(n_5207),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_5253),
.Y(n_5339)
);

INVx1_ASAP7_75t_L g5340 ( 
.A(n_5227),
.Y(n_5340)
);

AND2x2_ASAP7_75t_L g5341 ( 
.A(n_5206),
.B(n_5108),
.Y(n_5341)
);

OR2x2_ASAP7_75t_L g5342 ( 
.A(n_5226),
.B(n_5248),
.Y(n_5342)
);

AO21x2_ASAP7_75t_L g5343 ( 
.A1(n_5208),
.A2(n_5181),
.B(n_5095),
.Y(n_5343)
);

AND2x2_ASAP7_75t_L g5344 ( 
.A(n_5209),
.B(n_5136),
.Y(n_5344)
);

INVx2_ASAP7_75t_L g5345 ( 
.A(n_5245),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_5245),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5268),
.Y(n_5347)
);

BUFx3_ASAP7_75t_L g5348 ( 
.A(n_5189),
.Y(n_5348)
);

INVx2_ASAP7_75t_L g5349 ( 
.A(n_5214),
.Y(n_5349)
);

INVxp67_ASAP7_75t_SL g5350 ( 
.A(n_5244),
.Y(n_5350)
);

INVx2_ASAP7_75t_L g5351 ( 
.A(n_5185),
.Y(n_5351)
);

INVx1_ASAP7_75t_L g5352 ( 
.A(n_5212),
.Y(n_5352)
);

INVx2_ASAP7_75t_L g5353 ( 
.A(n_5186),
.Y(n_5353)
);

AO21x2_ASAP7_75t_L g5354 ( 
.A1(n_5235),
.A2(n_5162),
.B(n_5165),
.Y(n_5354)
);

NAND2xp5_ASAP7_75t_L g5355 ( 
.A(n_5250),
.B(n_5099),
.Y(n_5355)
);

OR2x2_ASAP7_75t_L g5356 ( 
.A(n_5204),
.B(n_5060),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5224),
.Y(n_5357)
);

AND2x4_ASAP7_75t_L g5358 ( 
.A(n_5188),
.B(n_5052),
.Y(n_5358)
);

AND2x2_ASAP7_75t_L g5359 ( 
.A(n_5203),
.B(n_5171),
.Y(n_5359)
);

BUFx2_ASAP7_75t_L g5360 ( 
.A(n_5284),
.Y(n_5360)
);

AND2x2_ASAP7_75t_L g5361 ( 
.A(n_5258),
.B(n_5102),
.Y(n_5361)
);

AND2x2_ASAP7_75t_L g5362 ( 
.A(n_5213),
.B(n_5060),
.Y(n_5362)
);

INVx2_ASAP7_75t_SL g5363 ( 
.A(n_5216),
.Y(n_5363)
);

AND2x2_ASAP7_75t_L g5364 ( 
.A(n_5222),
.B(n_5060),
.Y(n_5364)
);

HB1xp67_ASAP7_75t_L g5365 ( 
.A(n_5289),
.Y(n_5365)
);

HB1xp67_ASAP7_75t_L g5366 ( 
.A(n_5285),
.Y(n_5366)
);

AND2x2_ASAP7_75t_L g5367 ( 
.A(n_5259),
.B(n_5109),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_5259),
.B(n_5110),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_5350),
.B(n_5257),
.Y(n_5369)
);

AOI21xp33_ASAP7_75t_L g5370 ( 
.A1(n_5313),
.A2(n_5269),
.B(n_5251),
.Y(n_5370)
);

AND2x4_ASAP7_75t_L g5371 ( 
.A(n_5305),
.B(n_5243),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5365),
.B(n_5272),
.Y(n_5372)
);

OAI221xp5_ASAP7_75t_SL g5373 ( 
.A1(n_5311),
.A2(n_5236),
.B1(n_5255),
.B2(n_5197),
.C(n_5246),
.Y(n_5373)
);

NAND2xp33_ASAP7_75t_SL g5374 ( 
.A(n_5366),
.B(n_5201),
.Y(n_5374)
);

AND2x2_ASAP7_75t_L g5375 ( 
.A(n_5322),
.B(n_5238),
.Y(n_5375)
);

AND2x2_ASAP7_75t_L g5376 ( 
.A(n_5322),
.B(n_5210),
.Y(n_5376)
);

NAND2xp5_ASAP7_75t_SL g5377 ( 
.A(n_5308),
.B(n_5278),
.Y(n_5377)
);

AND2x2_ASAP7_75t_L g5378 ( 
.A(n_5304),
.B(n_5239),
.Y(n_5378)
);

NAND2xp5_ASAP7_75t_L g5379 ( 
.A(n_5360),
.B(n_5260),
.Y(n_5379)
);

AOI22xp33_ASAP7_75t_L g5380 ( 
.A1(n_5304),
.A2(n_5229),
.B1(n_5283),
.B2(n_5274),
.Y(n_5380)
);

NAND2xp5_ASAP7_75t_L g5381 ( 
.A(n_5360),
.B(n_5219),
.Y(n_5381)
);

NAND3xp33_ASAP7_75t_L g5382 ( 
.A(n_5362),
.B(n_5276),
.C(n_5287),
.Y(n_5382)
);

AND2x2_ASAP7_75t_L g5383 ( 
.A(n_5333),
.B(n_5232),
.Y(n_5383)
);

AND2x2_ASAP7_75t_L g5384 ( 
.A(n_5333),
.B(n_5241),
.Y(n_5384)
);

OAI22xp5_ASAP7_75t_L g5385 ( 
.A1(n_5295),
.A2(n_5282),
.B1(n_5246),
.B2(n_5096),
.Y(n_5385)
);

AOI22xp33_ASAP7_75t_L g5386 ( 
.A1(n_5354),
.A2(n_5264),
.B1(n_5292),
.B2(n_5267),
.Y(n_5386)
);

NOR3xp33_ASAP7_75t_L g5387 ( 
.A(n_5336),
.B(n_5247),
.C(n_5321),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_5354),
.B(n_5234),
.Y(n_5388)
);

OAI21xp33_ASAP7_75t_L g5389 ( 
.A1(n_5362),
.A2(n_5263),
.B(n_5187),
.Y(n_5389)
);

OAI221xp5_ASAP7_75t_L g5390 ( 
.A1(n_5323),
.A2(n_5270),
.B1(n_5252),
.B2(n_5184),
.C(n_5192),
.Y(n_5390)
);

NAND2xp5_ASAP7_75t_L g5391 ( 
.A(n_5354),
.B(n_5202),
.Y(n_5391)
);

AOI22xp33_ASAP7_75t_SL g5392 ( 
.A1(n_5343),
.A2(n_5217),
.B1(n_5196),
.B2(n_5233),
.Y(n_5392)
);

OAI221xp5_ASAP7_75t_L g5393 ( 
.A1(n_5309),
.A2(n_5265),
.B1(n_5256),
.B2(n_5262),
.C(n_5211),
.Y(n_5393)
);

OAI221xp5_ASAP7_75t_L g5394 ( 
.A1(n_5368),
.A2(n_5194),
.B1(n_5093),
.B2(n_5145),
.C(n_339),
.Y(n_5394)
);

NAND2xp5_ASAP7_75t_L g5395 ( 
.A(n_5339),
.B(n_335),
.Y(n_5395)
);

AOI22xp33_ASAP7_75t_SL g5396 ( 
.A1(n_5343),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_5396)
);

AND2x2_ASAP7_75t_L g5397 ( 
.A(n_5302),
.B(n_340),
.Y(n_5397)
);

AND2x2_ASAP7_75t_L g5398 ( 
.A(n_5302),
.B(n_340),
.Y(n_5398)
);

NAND3xp33_ASAP7_75t_L g5399 ( 
.A(n_5368),
.B(n_341),
.C(n_344),
.Y(n_5399)
);

AND2x2_ASAP7_75t_L g5400 ( 
.A(n_5348),
.B(n_5298),
.Y(n_5400)
);

AND2x2_ASAP7_75t_L g5401 ( 
.A(n_5348),
.B(n_341),
.Y(n_5401)
);

OAI21xp33_ASAP7_75t_L g5402 ( 
.A1(n_5367),
.A2(n_344),
.B(n_345),
.Y(n_5402)
);

OAI22xp5_ASAP7_75t_L g5403 ( 
.A1(n_5361),
.A2(n_351),
.B1(n_347),
.B2(n_349),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5339),
.B(n_347),
.Y(n_5404)
);

NAND4xp25_ASAP7_75t_L g5405 ( 
.A(n_5298),
.B(n_593),
.C(n_352),
.D(n_349),
.Y(n_5405)
);

OAI21xp5_ASAP7_75t_SL g5406 ( 
.A1(n_5367),
.A2(n_351),
.B(n_353),
.Y(n_5406)
);

AND2x2_ASAP7_75t_L g5407 ( 
.A(n_5315),
.B(n_354),
.Y(n_5407)
);

OAI21xp5_ASAP7_75t_SL g5408 ( 
.A1(n_5361),
.A2(n_354),
.B(n_355),
.Y(n_5408)
);

NAND2xp5_ASAP7_75t_L g5409 ( 
.A(n_5349),
.B(n_355),
.Y(n_5409)
);

NAND2xp5_ASAP7_75t_SL g5410 ( 
.A(n_5297),
.B(n_356),
.Y(n_5410)
);

NAND4xp25_ASAP7_75t_L g5411 ( 
.A(n_5342),
.B(n_360),
.C(n_356),
.D(n_357),
.Y(n_5411)
);

OAI221xp5_ASAP7_75t_SL g5412 ( 
.A1(n_5342),
.A2(n_5332),
.B1(n_5326),
.B2(n_5355),
.C(n_5297),
.Y(n_5412)
);

OAI21xp33_ASAP7_75t_SL g5413 ( 
.A1(n_5324),
.A2(n_357),
.B(n_362),
.Y(n_5413)
);

OAI221xp5_ASAP7_75t_L g5414 ( 
.A1(n_5338),
.A2(n_362),
.B1(n_363),
.B2(n_364),
.C(n_365),
.Y(n_5414)
);

AND2x2_ASAP7_75t_L g5415 ( 
.A(n_5315),
.B(n_5318),
.Y(n_5415)
);

NAND3xp33_ASAP7_75t_L g5416 ( 
.A(n_5296),
.B(n_364),
.C(n_366),
.Y(n_5416)
);

INVx2_ASAP7_75t_L g5417 ( 
.A(n_5378),
.Y(n_5417)
);

AO221x2_ASAP7_75t_L g5418 ( 
.A1(n_5382),
.A2(n_5340),
.B1(n_5343),
.B2(n_5347),
.C(n_5327),
.Y(n_5418)
);

INVx2_ASAP7_75t_L g5419 ( 
.A(n_5375),
.Y(n_5419)
);

OAI31xp33_ASAP7_75t_L g5420 ( 
.A1(n_5390),
.A2(n_5388),
.A3(n_5374),
.B(n_5386),
.Y(n_5420)
);

INVx3_ASAP7_75t_L g5421 ( 
.A(n_5371),
.Y(n_5421)
);

BUFx6f_ASAP7_75t_L g5422 ( 
.A(n_5397),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5396),
.Y(n_5423)
);

OAI31xp33_ASAP7_75t_SL g5424 ( 
.A1(n_5392),
.A2(n_5324),
.A3(n_5364),
.B(n_5331),
.Y(n_5424)
);

AOI221xp5_ASAP7_75t_L g5425 ( 
.A1(n_5412),
.A2(n_5364),
.B1(n_5303),
.B2(n_5331),
.C(n_5300),
.Y(n_5425)
);

OAI221xp5_ASAP7_75t_L g5426 ( 
.A1(n_5392),
.A2(n_5317),
.B1(n_5305),
.B2(n_5346),
.C(n_5349),
.Y(n_5426)
);

OR2x2_ASAP7_75t_L g5427 ( 
.A(n_5372),
.B(n_5294),
.Y(n_5427)
);

INVx3_ASAP7_75t_L g5428 ( 
.A(n_5371),
.Y(n_5428)
);

AND2x4_ASAP7_75t_L g5429 ( 
.A(n_5400),
.B(n_5305),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_5415),
.Y(n_5430)
);

AND2x2_ASAP7_75t_L g5431 ( 
.A(n_5376),
.B(n_5296),
.Y(n_5431)
);

NAND2xp5_ASAP7_75t_L g5432 ( 
.A(n_5386),
.B(n_5318),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_5396),
.Y(n_5433)
);

HB1xp67_ASAP7_75t_L g5434 ( 
.A(n_5384),
.Y(n_5434)
);

INVx2_ASAP7_75t_L g5435 ( 
.A(n_5391),
.Y(n_5435)
);

NOR3xp33_ASAP7_75t_SL g5436 ( 
.A(n_5412),
.B(n_5330),
.C(n_5328),
.Y(n_5436)
);

BUFx2_ASAP7_75t_L g5437 ( 
.A(n_5413),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_5406),
.B(n_5345),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5407),
.Y(n_5439)
);

AOI22xp33_ASAP7_75t_SL g5440 ( 
.A1(n_5385),
.A2(n_5303),
.B1(n_5305),
.B2(n_5317),
.Y(n_5440)
);

HB1xp67_ASAP7_75t_L g5441 ( 
.A(n_5369),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_5409),
.Y(n_5442)
);

NOR2x1_ASAP7_75t_L g5443 ( 
.A(n_5399),
.B(n_5300),
.Y(n_5443)
);

AND2x2_ASAP7_75t_L g5444 ( 
.A(n_5383),
.B(n_5300),
.Y(n_5444)
);

INVx2_ASAP7_75t_L g5445 ( 
.A(n_5398),
.Y(n_5445)
);

HB1xp67_ASAP7_75t_L g5446 ( 
.A(n_5379),
.Y(n_5446)
);

INVx2_ASAP7_75t_L g5447 ( 
.A(n_5401),
.Y(n_5447)
);

INVx2_ASAP7_75t_L g5448 ( 
.A(n_5377),
.Y(n_5448)
);

HB1xp67_ASAP7_75t_L g5449 ( 
.A(n_5410),
.Y(n_5449)
);

NAND2xp5_ASAP7_75t_L g5450 ( 
.A(n_5408),
.B(n_5345),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5431),
.B(n_5357),
.Y(n_5451)
);

OR2x2_ASAP7_75t_L g5452 ( 
.A(n_5432),
.B(n_5381),
.Y(n_5452)
);

OR2x2_ASAP7_75t_L g5453 ( 
.A(n_5434),
.B(n_5411),
.Y(n_5453)
);

NAND2xp5_ASAP7_75t_L g5454 ( 
.A(n_5423),
.B(n_5387),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_5439),
.Y(n_5455)
);

AND2x2_ASAP7_75t_L g5456 ( 
.A(n_5431),
.B(n_5334),
.Y(n_5456)
);

INVx1_ASAP7_75t_L g5457 ( 
.A(n_5439),
.Y(n_5457)
);

NAND2xp5_ASAP7_75t_L g5458 ( 
.A(n_5423),
.B(n_5433),
.Y(n_5458)
);

AND2x4_ASAP7_75t_L g5459 ( 
.A(n_5421),
.B(n_5305),
.Y(n_5459)
);

OR2x2_ASAP7_75t_L g5460 ( 
.A(n_5445),
.B(n_5387),
.Y(n_5460)
);

AND2x2_ASAP7_75t_L g5461 ( 
.A(n_5444),
.B(n_5334),
.Y(n_5461)
);

NOR2x1_ASAP7_75t_L g5462 ( 
.A(n_5421),
.B(n_5416),
.Y(n_5462)
);

INVx1_ASAP7_75t_SL g5463 ( 
.A(n_5421),
.Y(n_5463)
);

AND2x2_ASAP7_75t_SL g5464 ( 
.A(n_5433),
.B(n_5380),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5430),
.Y(n_5465)
);

INVx1_ASAP7_75t_L g5466 ( 
.A(n_5430),
.Y(n_5466)
);

AND2x2_ASAP7_75t_L g5467 ( 
.A(n_5444),
.B(n_5352),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5445),
.Y(n_5468)
);

AND2x2_ASAP7_75t_L g5469 ( 
.A(n_5419),
.B(n_5370),
.Y(n_5469)
);

INVx1_ASAP7_75t_L g5470 ( 
.A(n_5447),
.Y(n_5470)
);

AND2x4_ASAP7_75t_L g5471 ( 
.A(n_5428),
.B(n_5312),
.Y(n_5471)
);

BUFx2_ASAP7_75t_SL g5472 ( 
.A(n_5428),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_5447),
.Y(n_5473)
);

AND2x2_ASAP7_75t_L g5474 ( 
.A(n_5456),
.B(n_5461),
.Y(n_5474)
);

INVx1_ASAP7_75t_L g5475 ( 
.A(n_5463),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5463),
.Y(n_5476)
);

INVx4_ASAP7_75t_L g5477 ( 
.A(n_5459),
.Y(n_5477)
);

NAND2xp5_ASAP7_75t_SL g5478 ( 
.A(n_5454),
.B(n_5420),
.Y(n_5478)
);

AND2x2_ASAP7_75t_L g5479 ( 
.A(n_5451),
.B(n_5419),
.Y(n_5479)
);

AOI22xp33_ASAP7_75t_L g5480 ( 
.A1(n_5464),
.A2(n_5418),
.B1(n_5420),
.B2(n_5437),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5472),
.Y(n_5481)
);

AND2x2_ASAP7_75t_L g5482 ( 
.A(n_5467),
.B(n_5422),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_L g5483 ( 
.A(n_5464),
.B(n_5436),
.Y(n_5483)
);

AND2x2_ASAP7_75t_L g5484 ( 
.A(n_5469),
.B(n_5422),
.Y(n_5484)
);

NOR2xp67_ASAP7_75t_L g5485 ( 
.A(n_5471),
.B(n_5428),
.Y(n_5485)
);

AND2x2_ASAP7_75t_L g5486 ( 
.A(n_5471),
.B(n_5422),
.Y(n_5486)
);

NAND4xp25_ASAP7_75t_L g5487 ( 
.A(n_5454),
.B(n_5440),
.C(n_5425),
.D(n_5424),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_5468),
.Y(n_5488)
);

AND2x4_ASAP7_75t_L g5489 ( 
.A(n_5459),
.B(n_5429),
.Y(n_5489)
);

INVx2_ASAP7_75t_SL g5490 ( 
.A(n_5459),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5470),
.Y(n_5491)
);

NAND2xp5_ASAP7_75t_L g5492 ( 
.A(n_5458),
.B(n_5437),
.Y(n_5492)
);

AND2x2_ASAP7_75t_L g5493 ( 
.A(n_5462),
.B(n_5422),
.Y(n_5493)
);

NOR3xp33_ASAP7_75t_L g5494 ( 
.A(n_5458),
.B(n_5426),
.C(n_5373),
.Y(n_5494)
);

INVx1_ASAP7_75t_L g5495 ( 
.A(n_5473),
.Y(n_5495)
);

NOR2xp33_ASAP7_75t_L g5496 ( 
.A(n_5481),
.B(n_5422),
.Y(n_5496)
);

CKINVDCx5p33_ASAP7_75t_R g5497 ( 
.A(n_5489),
.Y(n_5497)
);

CKINVDCx5p33_ASAP7_75t_R g5498 ( 
.A(n_5489),
.Y(n_5498)
);

NAND2x1_ASAP7_75t_L g5499 ( 
.A(n_5477),
.B(n_5429),
.Y(n_5499)
);

AND2x4_ASAP7_75t_L g5500 ( 
.A(n_5485),
.B(n_5429),
.Y(n_5500)
);

NOR2xp33_ASAP7_75t_L g5501 ( 
.A(n_5487),
.B(n_5450),
.Y(n_5501)
);

CKINVDCx5p33_ASAP7_75t_R g5502 ( 
.A(n_5486),
.Y(n_5502)
);

AO221x2_ASAP7_75t_L g5503 ( 
.A1(n_5483),
.A2(n_5448),
.B1(n_5455),
.B2(n_5457),
.C(n_5442),
.Y(n_5503)
);

OAI22xp33_ASAP7_75t_L g5504 ( 
.A1(n_5483),
.A2(n_5393),
.B1(n_5394),
.B2(n_5449),
.Y(n_5504)
);

OAI221xp5_ASAP7_75t_L g5505 ( 
.A1(n_5480),
.A2(n_5373),
.B1(n_5443),
.B2(n_5389),
.C(n_5448),
.Y(n_5505)
);

NAND2xp5_ASAP7_75t_L g5506 ( 
.A(n_5493),
.B(n_5417),
.Y(n_5506)
);

OR2x2_ASAP7_75t_L g5507 ( 
.A(n_5492),
.B(n_5453),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_5480),
.B(n_5417),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_5482),
.B(n_5446),
.Y(n_5509)
);

NAND2xp5_ASAP7_75t_L g5510 ( 
.A(n_5474),
.B(n_5443),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_5484),
.B(n_5438),
.Y(n_5511)
);

NAND2xp5_ASAP7_75t_L g5512 ( 
.A(n_5497),
.B(n_5490),
.Y(n_5512)
);

NOR2xp33_ASAP7_75t_L g5513 ( 
.A(n_5505),
.B(n_5478),
.Y(n_5513)
);

NOR2xp33_ASAP7_75t_L g5514 ( 
.A(n_5498),
.B(n_5478),
.Y(n_5514)
);

AND2x2_ASAP7_75t_L g5515 ( 
.A(n_5500),
.B(n_5479),
.Y(n_5515)
);

AND2x2_ASAP7_75t_L g5516 ( 
.A(n_5496),
.B(n_5441),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_5501),
.B(n_5475),
.Y(n_5517)
);

OAI21xp33_ASAP7_75t_L g5518 ( 
.A1(n_5511),
.A2(n_5494),
.B(n_5492),
.Y(n_5518)
);

OAI21xp33_ASAP7_75t_SL g5519 ( 
.A1(n_5508),
.A2(n_5477),
.B(n_5476),
.Y(n_5519)
);

NAND2xp5_ASAP7_75t_L g5520 ( 
.A(n_5502),
.B(n_5494),
.Y(n_5520)
);

AND2x2_ASAP7_75t_L g5521 ( 
.A(n_5510),
.B(n_5460),
.Y(n_5521)
);

INVx2_ASAP7_75t_L g5522 ( 
.A(n_5499),
.Y(n_5522)
);

NOR2xp33_ASAP7_75t_L g5523 ( 
.A(n_5506),
.B(n_5452),
.Y(n_5523)
);

INVx1_ASAP7_75t_L g5524 ( 
.A(n_5515),
.Y(n_5524)
);

AND2x2_ASAP7_75t_L g5525 ( 
.A(n_5516),
.B(n_5509),
.Y(n_5525)
);

AND2x2_ASAP7_75t_L g5526 ( 
.A(n_5521),
.B(n_5442),
.Y(n_5526)
);

AND2x2_ASAP7_75t_L g5527 ( 
.A(n_5514),
.B(n_5507),
.Y(n_5527)
);

INVxp67_ASAP7_75t_L g5528 ( 
.A(n_5522),
.Y(n_5528)
);

OR2x2_ASAP7_75t_L g5529 ( 
.A(n_5520),
.B(n_5503),
.Y(n_5529)
);

OR2x2_ASAP7_75t_L g5530 ( 
.A(n_5517),
.B(n_5503),
.Y(n_5530)
);

AOI21xp33_ASAP7_75t_SL g5531 ( 
.A1(n_5513),
.A2(n_5504),
.B(n_5491),
.Y(n_5531)
);

OAI21xp33_ASAP7_75t_SL g5532 ( 
.A1(n_5523),
.A2(n_5435),
.B(n_5465),
.Y(n_5532)
);

INVx1_ASAP7_75t_SL g5533 ( 
.A(n_5512),
.Y(n_5533)
);

AOI22xp5_ASAP7_75t_L g5534 ( 
.A1(n_5518),
.A2(n_5418),
.B1(n_5466),
.B2(n_5435),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5519),
.Y(n_5535)
);

OAI22xp33_ASAP7_75t_L g5536 ( 
.A1(n_5520),
.A2(n_5427),
.B1(n_5335),
.B2(n_5403),
.Y(n_5536)
);

INVxp67_ASAP7_75t_SL g5537 ( 
.A(n_5514),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_5515),
.Y(n_5538)
);

INVxp67_ASAP7_75t_SL g5539 ( 
.A(n_5530),
.Y(n_5539)
);

NOR3xp33_ASAP7_75t_L g5540 ( 
.A(n_5531),
.B(n_5495),
.C(n_5488),
.Y(n_5540)
);

AOI211xp5_ASAP7_75t_L g5541 ( 
.A1(n_5531),
.A2(n_5427),
.B(n_5414),
.C(n_5402),
.Y(n_5541)
);

INVx1_ASAP7_75t_L g5542 ( 
.A(n_5524),
.Y(n_5542)
);

OR2x2_ASAP7_75t_L g5543 ( 
.A(n_5538),
.B(n_5418),
.Y(n_5543)
);

AOI22xp5_ASAP7_75t_L g5544 ( 
.A1(n_5537),
.A2(n_5418),
.B1(n_5405),
.B2(n_5335),
.Y(n_5544)
);

OAI22xp33_ASAP7_75t_L g5545 ( 
.A1(n_5534),
.A2(n_5335),
.B1(n_5317),
.B2(n_5356),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5525),
.Y(n_5546)
);

INVx1_ASAP7_75t_L g5547 ( 
.A(n_5527),
.Y(n_5547)
);

AOI22xp33_ASAP7_75t_L g5548 ( 
.A1(n_5535),
.A2(n_5356),
.B1(n_5312),
.B2(n_5353),
.Y(n_5548)
);

INVx1_ASAP7_75t_L g5549 ( 
.A(n_5526),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_5528),
.Y(n_5550)
);

A2O1A1Ixp33_ASAP7_75t_L g5551 ( 
.A1(n_5544),
.A2(n_5541),
.B(n_5532),
.C(n_5540),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5547),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5543),
.Y(n_5553)
);

INVx1_ASAP7_75t_SL g5554 ( 
.A(n_5549),
.Y(n_5554)
);

NAND2xp5_ASAP7_75t_L g5555 ( 
.A(n_5546),
.B(n_5536),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5542),
.Y(n_5556)
);

INVx1_ASAP7_75t_L g5557 ( 
.A(n_5550),
.Y(n_5557)
);

OR2x2_ASAP7_75t_L g5558 ( 
.A(n_5539),
.B(n_5533),
.Y(n_5558)
);

AO22x2_ASAP7_75t_L g5559 ( 
.A1(n_5545),
.A2(n_5529),
.B1(n_5395),
.B2(n_5404),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_5548),
.Y(n_5560)
);

AND2x2_ASAP7_75t_L g5561 ( 
.A(n_5547),
.B(n_5337),
.Y(n_5561)
);

NAND2xp5_ASAP7_75t_L g5562 ( 
.A(n_5561),
.B(n_5314),
.Y(n_5562)
);

NAND2xp5_ASAP7_75t_L g5563 ( 
.A(n_5554),
.B(n_5316),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5558),
.Y(n_5564)
);

HB1xp67_ASAP7_75t_L g5565 ( 
.A(n_5559),
.Y(n_5565)
);

INVx1_ASAP7_75t_L g5566 ( 
.A(n_5559),
.Y(n_5566)
);

INVx1_ASAP7_75t_L g5567 ( 
.A(n_5552),
.Y(n_5567)
);

NAND3xp33_ASAP7_75t_SL g5568 ( 
.A(n_5551),
.B(n_5299),
.C(n_5301),
.Y(n_5568)
);

INVx1_ASAP7_75t_SL g5569 ( 
.A(n_5555),
.Y(n_5569)
);

OAI31xp33_ASAP7_75t_L g5570 ( 
.A1(n_5560),
.A2(n_5301),
.A3(n_5310),
.B(n_5307),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_L g5571 ( 
.A(n_5557),
.B(n_5325),
.Y(n_5571)
);

AOI221xp5_ASAP7_75t_L g5572 ( 
.A1(n_5556),
.A2(n_5307),
.B1(n_5310),
.B2(n_5319),
.C(n_5312),
.Y(n_5572)
);

NAND2xp5_ASAP7_75t_L g5573 ( 
.A(n_5553),
.B(n_5319),
.Y(n_5573)
);

INVx1_ASAP7_75t_L g5574 ( 
.A(n_5561),
.Y(n_5574)
);

OR2x2_ASAP7_75t_L g5575 ( 
.A(n_5558),
.B(n_5351),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_5561),
.B(n_5299),
.Y(n_5576)
);

AND2x2_ASAP7_75t_L g5577 ( 
.A(n_5561),
.B(n_5306),
.Y(n_5577)
);

XNOR2xp5_ASAP7_75t_L g5578 ( 
.A(n_5561),
.B(n_366),
.Y(n_5578)
);

AOI222xp33_ASAP7_75t_L g5579 ( 
.A1(n_5560),
.A2(n_5351),
.B1(n_5353),
.B2(n_5363),
.C1(n_5358),
.C2(n_5344),
.Y(n_5579)
);

OAI322xp33_ASAP7_75t_L g5580 ( 
.A1(n_5558),
.A2(n_5363),
.A3(n_5344),
.B1(n_5306),
.B2(n_5359),
.C1(n_5320),
.C2(n_5341),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_5577),
.Y(n_5581)
);

INVx1_ASAP7_75t_L g5582 ( 
.A(n_5576),
.Y(n_5582)
);

INVxp33_ASAP7_75t_SL g5583 ( 
.A(n_5565),
.Y(n_5583)
);

INVx1_ASAP7_75t_L g5584 ( 
.A(n_5578),
.Y(n_5584)
);

INVx1_ASAP7_75t_SL g5585 ( 
.A(n_5575),
.Y(n_5585)
);

INVx1_ASAP7_75t_SL g5586 ( 
.A(n_5569),
.Y(n_5586)
);

INVx1_ASAP7_75t_L g5587 ( 
.A(n_5566),
.Y(n_5587)
);

BUFx2_ASAP7_75t_L g5588 ( 
.A(n_5574),
.Y(n_5588)
);

INVx1_ASAP7_75t_L g5589 ( 
.A(n_5564),
.Y(n_5589)
);

INVx1_ASAP7_75t_L g5590 ( 
.A(n_5563),
.Y(n_5590)
);

INVx1_ASAP7_75t_L g5591 ( 
.A(n_5573),
.Y(n_5591)
);

HB1xp67_ASAP7_75t_L g5592 ( 
.A(n_5567),
.Y(n_5592)
);

NAND2x1_ASAP7_75t_SL g5593 ( 
.A(n_5568),
.B(n_5320),
.Y(n_5593)
);

HB1xp67_ASAP7_75t_L g5594 ( 
.A(n_5562),
.Y(n_5594)
);

CKINVDCx20_ASAP7_75t_R g5595 ( 
.A(n_5571),
.Y(n_5595)
);

INVx1_ASAP7_75t_L g5596 ( 
.A(n_5580),
.Y(n_5596)
);

INVx1_ASAP7_75t_SL g5597 ( 
.A(n_5570),
.Y(n_5597)
);

INVx1_ASAP7_75t_L g5598 ( 
.A(n_5572),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_5579),
.Y(n_5599)
);

INVx2_ASAP7_75t_SL g5600 ( 
.A(n_5577),
.Y(n_5600)
);

AND2x4_ASAP7_75t_L g5601 ( 
.A(n_5577),
.B(n_5358),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_5577),
.Y(n_5602)
);

INVx1_ASAP7_75t_L g5603 ( 
.A(n_5577),
.Y(n_5603)
);

XOR2x2_ASAP7_75t_L g5604 ( 
.A(n_5578),
.B(n_367),
.Y(n_5604)
);

INVx1_ASAP7_75t_L g5605 ( 
.A(n_5577),
.Y(n_5605)
);

INVx1_ASAP7_75t_L g5606 ( 
.A(n_5577),
.Y(n_5606)
);

INVx1_ASAP7_75t_L g5607 ( 
.A(n_5577),
.Y(n_5607)
);

OAI21xp33_ASAP7_75t_SL g5608 ( 
.A1(n_5593),
.A2(n_5359),
.B(n_5341),
.Y(n_5608)
);

A2O1A1Ixp33_ASAP7_75t_L g5609 ( 
.A1(n_5596),
.A2(n_5358),
.B(n_5320),
.C(n_5329),
.Y(n_5609)
);

AOI22xp33_ASAP7_75t_SL g5610 ( 
.A1(n_5583),
.A2(n_5329),
.B1(n_369),
.B2(n_370),
.Y(n_5610)
);

INVx1_ASAP7_75t_L g5611 ( 
.A(n_5604),
.Y(n_5611)
);

OR2x2_ASAP7_75t_L g5612 ( 
.A(n_5600),
.B(n_5329),
.Y(n_5612)
);

NAND3xp33_ASAP7_75t_SL g5613 ( 
.A(n_5586),
.B(n_367),
.C(n_371),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5592),
.Y(n_5614)
);

AOI22xp5_ASAP7_75t_SL g5615 ( 
.A1(n_5595),
.A2(n_5329),
.B1(n_372),
.B2(n_373),
.Y(n_5615)
);

INVx1_ASAP7_75t_L g5616 ( 
.A(n_5588),
.Y(n_5616)
);

AOI21xp5_ASAP7_75t_SL g5617 ( 
.A1(n_5589),
.A2(n_371),
.B(n_374),
.Y(n_5617)
);

CKINVDCx5p33_ASAP7_75t_R g5618 ( 
.A(n_5581),
.Y(n_5618)
);

AOI221xp5_ASAP7_75t_L g5619 ( 
.A1(n_5587),
.A2(n_5329),
.B1(n_377),
.B2(n_378),
.C(n_379),
.Y(n_5619)
);

OAI22xp5_ASAP7_75t_L g5620 ( 
.A1(n_5599),
.A2(n_374),
.B1(n_380),
.B2(n_381),
.Y(n_5620)
);

HB1xp67_ASAP7_75t_L g5621 ( 
.A(n_5601),
.Y(n_5621)
);

AOI221xp5_ASAP7_75t_L g5622 ( 
.A1(n_5597),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.C(n_386),
.Y(n_5622)
);

OAI22xp5_ASAP7_75t_L g5623 ( 
.A1(n_5602),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_5623)
);

AOI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_5603),
.A2(n_386),
.B1(n_388),
.B2(n_390),
.Y(n_5624)
);

INVx1_ASAP7_75t_L g5625 ( 
.A(n_5605),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5601),
.B(n_388),
.Y(n_5626)
);

OAI211xp5_ASAP7_75t_L g5627 ( 
.A1(n_5597),
.A2(n_391),
.B(n_393),
.C(n_394),
.Y(n_5627)
);

INVx2_ASAP7_75t_SL g5628 ( 
.A(n_5606),
.Y(n_5628)
);

OAI21x1_ASAP7_75t_L g5629 ( 
.A1(n_5607),
.A2(n_391),
.B(n_393),
.Y(n_5629)
);

OAI21xp5_ASAP7_75t_L g5630 ( 
.A1(n_5585),
.A2(n_394),
.B(n_395),
.Y(n_5630)
);

OAI21xp33_ASAP7_75t_L g5631 ( 
.A1(n_5582),
.A2(n_396),
.B(n_397),
.Y(n_5631)
);

O2A1O1Ixp33_ASAP7_75t_SL g5632 ( 
.A1(n_5598),
.A2(n_5590),
.B(n_5594),
.C(n_5584),
.Y(n_5632)
);

NAND2xp5_ASAP7_75t_L g5633 ( 
.A(n_5591),
.B(n_396),
.Y(n_5633)
);

NAND2xp5_ASAP7_75t_L g5634 ( 
.A(n_5601),
.B(n_398),
.Y(n_5634)
);

AOI321xp33_ASAP7_75t_L g5635 ( 
.A1(n_5596),
.A2(n_398),
.A3(n_399),
.B1(n_401),
.B2(n_403),
.C(n_407),
.Y(n_5635)
);

INVx2_ASAP7_75t_L g5636 ( 
.A(n_5601),
.Y(n_5636)
);

AOI311xp33_ASAP7_75t_L g5637 ( 
.A1(n_5616),
.A2(n_403),
.A3(n_408),
.B(n_409),
.C(n_410),
.Y(n_5637)
);

AOI21xp5_ASAP7_75t_L g5638 ( 
.A1(n_5632),
.A2(n_408),
.B(n_409),
.Y(n_5638)
);

AOI21xp33_ASAP7_75t_L g5639 ( 
.A1(n_5628),
.A2(n_411),
.B(n_412),
.Y(n_5639)
);

CKINVDCx16_ASAP7_75t_R g5640 ( 
.A(n_5621),
.Y(n_5640)
);

CKINVDCx20_ASAP7_75t_R g5641 ( 
.A(n_5618),
.Y(n_5641)
);

NAND2xp5_ASAP7_75t_L g5642 ( 
.A(n_5622),
.B(n_411),
.Y(n_5642)
);

OAI211xp5_ASAP7_75t_SL g5643 ( 
.A1(n_5614),
.A2(n_412),
.B(n_413),
.C(n_414),
.Y(n_5643)
);

OA22x2_ASAP7_75t_L g5644 ( 
.A1(n_5617),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_5644)
);

OAI211xp5_ASAP7_75t_L g5645 ( 
.A1(n_5635),
.A2(n_415),
.B(n_416),
.C(n_417),
.Y(n_5645)
);

NAND4xp75_ASAP7_75t_L g5646 ( 
.A(n_5625),
.B(n_417),
.C(n_418),
.D(n_419),
.Y(n_5646)
);

NAND3xp33_ASAP7_75t_L g5647 ( 
.A(n_5627),
.B(n_419),
.C(n_420),
.Y(n_5647)
);

NAND2xp5_ASAP7_75t_L g5648 ( 
.A(n_5636),
.B(n_420),
.Y(n_5648)
);

NOR4xp75_ASAP7_75t_L g5649 ( 
.A(n_5620),
.B(n_421),
.C(n_423),
.D(n_424),
.Y(n_5649)
);

NOR2xp33_ASAP7_75t_R g5650 ( 
.A(n_5613),
.B(n_5611),
.Y(n_5650)
);

NAND2xp5_ASAP7_75t_L g5651 ( 
.A(n_5608),
.B(n_421),
.Y(n_5651)
);

OAI21xp33_ASAP7_75t_SL g5652 ( 
.A1(n_5634),
.A2(n_423),
.B(n_424),
.Y(n_5652)
);

OAI21xp5_ASAP7_75t_L g5653 ( 
.A1(n_5609),
.A2(n_425),
.B(n_426),
.Y(n_5653)
);

OAI321xp33_ASAP7_75t_L g5654 ( 
.A1(n_5612),
.A2(n_425),
.A3(n_428),
.B1(n_430),
.B2(n_431),
.C(n_432),
.Y(n_5654)
);

INVx1_ASAP7_75t_SL g5655 ( 
.A(n_5626),
.Y(n_5655)
);

AOI22xp5_ASAP7_75t_L g5656 ( 
.A1(n_5631),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_5656)
);

OAI22xp33_ASAP7_75t_SL g5657 ( 
.A1(n_5633),
.A2(n_433),
.B1(n_434),
.B2(n_435),
.Y(n_5657)
);

OAI211xp5_ASAP7_75t_L g5658 ( 
.A1(n_5630),
.A2(n_436),
.B(n_437),
.C(n_438),
.Y(n_5658)
);

NAND2xp5_ASAP7_75t_SL g5659 ( 
.A(n_5610),
.B(n_436),
.Y(n_5659)
);

NAND2xp5_ASAP7_75t_L g5660 ( 
.A(n_5629),
.B(n_437),
.Y(n_5660)
);

AOI22xp5_ASAP7_75t_L g5661 ( 
.A1(n_5640),
.A2(n_5641),
.B1(n_5645),
.B2(n_5655),
.Y(n_5661)
);

AOI211xp5_ASAP7_75t_L g5662 ( 
.A1(n_5658),
.A2(n_5623),
.B(n_5619),
.C(n_5624),
.Y(n_5662)
);

AOI221x1_ASAP7_75t_L g5663 ( 
.A1(n_5638),
.A2(n_5615),
.B1(n_440),
.B2(n_441),
.C(n_442),
.Y(n_5663)
);

AND5x1_ASAP7_75t_L g5664 ( 
.A(n_5656),
.B(n_439),
.C(n_440),
.D(n_441),
.E(n_442),
.Y(n_5664)
);

AOI22xp5_ASAP7_75t_L g5665 ( 
.A1(n_5643),
.A2(n_5644),
.B1(n_5647),
.B2(n_5659),
.Y(n_5665)
);

OAI22xp5_ASAP7_75t_L g5666 ( 
.A1(n_5648),
.A2(n_443),
.B1(n_446),
.B2(n_448),
.Y(n_5666)
);

OAI221xp5_ASAP7_75t_L g5667 ( 
.A1(n_5652),
.A2(n_443),
.B1(n_446),
.B2(n_449),
.C(n_450),
.Y(n_5667)
);

OAI21xp33_ASAP7_75t_L g5668 ( 
.A1(n_5650),
.A2(n_449),
.B(n_450),
.Y(n_5668)
);

OAI22xp5_ASAP7_75t_L g5669 ( 
.A1(n_5642),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.Y(n_5669)
);

OAI21xp5_ASAP7_75t_L g5670 ( 
.A1(n_5651),
.A2(n_452),
.B(n_454),
.Y(n_5670)
);

NAND3xp33_ASAP7_75t_L g5671 ( 
.A(n_5637),
.B(n_456),
.C(n_458),
.Y(n_5671)
);

HB1xp67_ASAP7_75t_L g5672 ( 
.A(n_5649),
.Y(n_5672)
);

AOI21xp33_ASAP7_75t_L g5673 ( 
.A1(n_5660),
.A2(n_458),
.B(n_459),
.Y(n_5673)
);

OAI211xp5_ASAP7_75t_L g5674 ( 
.A1(n_5653),
.A2(n_459),
.B(n_460),
.C(n_462),
.Y(n_5674)
);

NAND3xp33_ASAP7_75t_L g5675 ( 
.A(n_5639),
.B(n_460),
.C(n_462),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5657),
.Y(n_5676)
);

OAI221xp5_ASAP7_75t_L g5677 ( 
.A1(n_5654),
.A2(n_5646),
.B1(n_465),
.B2(n_466),
.C(n_467),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_5644),
.Y(n_5678)
);

OAI22xp33_ASAP7_75t_L g5679 ( 
.A1(n_5661),
.A2(n_464),
.B1(n_469),
.B2(n_470),
.Y(n_5679)
);

BUFx2_ASAP7_75t_L g5680 ( 
.A(n_5672),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_L g5681 ( 
.A(n_5668),
.B(n_469),
.Y(n_5681)
);

XOR2x2_ASAP7_75t_L g5682 ( 
.A(n_5664),
.B(n_470),
.Y(n_5682)
);

AOI22xp5_ASAP7_75t_L g5683 ( 
.A1(n_5678),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5671),
.Y(n_5684)
);

INVx1_ASAP7_75t_L g5685 ( 
.A(n_5663),
.Y(n_5685)
);

HB1xp67_ASAP7_75t_L g5686 ( 
.A(n_5666),
.Y(n_5686)
);

AND2x2_ASAP7_75t_L g5687 ( 
.A(n_5676),
.B(n_472),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5667),
.Y(n_5688)
);

INVx1_ASAP7_75t_L g5689 ( 
.A(n_5675),
.Y(n_5689)
);

INVx1_ASAP7_75t_L g5690 ( 
.A(n_5674),
.Y(n_5690)
);

AOI22xp5_ASAP7_75t_L g5691 ( 
.A1(n_5665),
.A2(n_592),
.B1(n_475),
.B2(n_476),
.Y(n_5691)
);

NOR3xp33_ASAP7_75t_SL g5692 ( 
.A(n_5677),
.B(n_474),
.C(n_477),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5669),
.Y(n_5693)
);

NAND2xp5_ASAP7_75t_L g5694 ( 
.A(n_5670),
.B(n_478),
.Y(n_5694)
);

OR2x2_ASAP7_75t_L g5695 ( 
.A(n_5681),
.B(n_5673),
.Y(n_5695)
);

NOR2xp67_ASAP7_75t_SL g5696 ( 
.A(n_5685),
.B(n_5662),
.Y(n_5696)
);

INVx1_ASAP7_75t_L g5697 ( 
.A(n_5682),
.Y(n_5697)
);

NOR2xp33_ASAP7_75t_L g5698 ( 
.A(n_5687),
.B(n_478),
.Y(n_5698)
);

INVx5_ASAP7_75t_L g5699 ( 
.A(n_5680),
.Y(n_5699)
);

NAND3x1_ASAP7_75t_L g5700 ( 
.A(n_5694),
.B(n_479),
.C(n_481),
.Y(n_5700)
);

INVx5_ASAP7_75t_L g5701 ( 
.A(n_5679),
.Y(n_5701)
);

AND2x2_ASAP7_75t_L g5702 ( 
.A(n_5692),
.B(n_482),
.Y(n_5702)
);

INVx1_ASAP7_75t_SL g5703 ( 
.A(n_5691),
.Y(n_5703)
);

NAND5xp2_ASAP7_75t_L g5704 ( 
.A(n_5684),
.B(n_482),
.C(n_484),
.D(n_486),
.E(n_487),
.Y(n_5704)
);

NAND2x1p5_ASAP7_75t_L g5705 ( 
.A(n_5690),
.B(n_488),
.Y(n_5705)
);

NAND3xp33_ASAP7_75t_SL g5706 ( 
.A(n_5689),
.B(n_5688),
.C(n_5693),
.Y(n_5706)
);

NAND2xp5_ASAP7_75t_L g5707 ( 
.A(n_5683),
.B(n_5686),
.Y(n_5707)
);

INVx4_ASAP7_75t_SL g5708 ( 
.A(n_5687),
.Y(n_5708)
);

NOR2x1_ASAP7_75t_L g5709 ( 
.A(n_5685),
.B(n_488),
.Y(n_5709)
);

AOI211xp5_ASAP7_75t_L g5710 ( 
.A1(n_5679),
.A2(n_489),
.B(n_490),
.C(n_491),
.Y(n_5710)
);

NOR3xp33_ASAP7_75t_L g5711 ( 
.A(n_5680),
.B(n_592),
.C(n_490),
.Y(n_5711)
);

NAND2xp5_ASAP7_75t_SL g5712 ( 
.A(n_5699),
.B(n_489),
.Y(n_5712)
);

NAND3xp33_ASAP7_75t_L g5713 ( 
.A(n_5699),
.B(n_491),
.C(n_492),
.Y(n_5713)
);

NAND2xp5_ASAP7_75t_SL g5714 ( 
.A(n_5701),
.B(n_492),
.Y(n_5714)
);

NAND2xp5_ASAP7_75t_L g5715 ( 
.A(n_5698),
.B(n_493),
.Y(n_5715)
);

NOR2xp33_ASAP7_75t_R g5716 ( 
.A(n_5706),
.B(n_495),
.Y(n_5716)
);

NAND2xp5_ASAP7_75t_SL g5717 ( 
.A(n_5710),
.B(n_495),
.Y(n_5717)
);

XNOR2xp5_ASAP7_75t_L g5718 ( 
.A(n_5700),
.B(n_497),
.Y(n_5718)
);

NAND2xp5_ASAP7_75t_SL g5719 ( 
.A(n_5711),
.B(n_498),
.Y(n_5719)
);

NAND2xp5_ASAP7_75t_L g5720 ( 
.A(n_5705),
.B(n_498),
.Y(n_5720)
);

NOR2xp33_ASAP7_75t_R g5721 ( 
.A(n_5697),
.B(n_499),
.Y(n_5721)
);

NAND2xp33_ASAP7_75t_SL g5722 ( 
.A(n_5696),
.B(n_499),
.Y(n_5722)
);

NAND2xp5_ASAP7_75t_L g5723 ( 
.A(n_5709),
.B(n_500),
.Y(n_5723)
);

NAND2xp5_ASAP7_75t_L g5724 ( 
.A(n_5702),
.B(n_500),
.Y(n_5724)
);

HB1xp67_ASAP7_75t_L g5725 ( 
.A(n_5721),
.Y(n_5725)
);

NOR2xp33_ASAP7_75t_L g5726 ( 
.A(n_5720),
.B(n_5704),
.Y(n_5726)
);

OAI211xp5_ASAP7_75t_L g5727 ( 
.A1(n_5716),
.A2(n_5714),
.B(n_5722),
.C(n_5723),
.Y(n_5727)
);

NAND2xp5_ASAP7_75t_L g5728 ( 
.A(n_5712),
.B(n_5708),
.Y(n_5728)
);

NAND4xp25_ASAP7_75t_SL g5729 ( 
.A(n_5724),
.B(n_5703),
.C(n_5707),
.D(n_5695),
.Y(n_5729)
);

AO22x2_ASAP7_75t_L g5730 ( 
.A1(n_5715),
.A2(n_5713),
.B1(n_5719),
.B2(n_5717),
.Y(n_5730)
);

OAI221xp5_ASAP7_75t_L g5731 ( 
.A1(n_5718),
.A2(n_501),
.B1(n_503),
.B2(n_505),
.C(n_509),
.Y(n_5731)
);

INVx1_ASAP7_75t_L g5732 ( 
.A(n_5725),
.Y(n_5732)
);

AOI22xp5_ASAP7_75t_L g5733 ( 
.A1(n_5729),
.A2(n_505),
.B1(n_510),
.B2(n_511),
.Y(n_5733)
);

INVx1_ASAP7_75t_SL g5734 ( 
.A(n_5728),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5731),
.Y(n_5735)
);

INVx1_ASAP7_75t_L g5736 ( 
.A(n_5726),
.Y(n_5736)
);

OAI311xp33_ASAP7_75t_L g5737 ( 
.A1(n_5727),
.A2(n_510),
.A3(n_512),
.B1(n_513),
.C1(n_514),
.Y(n_5737)
);

INVx1_ASAP7_75t_L g5738 ( 
.A(n_5730),
.Y(n_5738)
);

NAND2x1_ASAP7_75t_L g5739 ( 
.A(n_5733),
.B(n_514),
.Y(n_5739)
);

NAND2xp5_ASAP7_75t_L g5740 ( 
.A(n_5738),
.B(n_515),
.Y(n_5740)
);

INVx2_ASAP7_75t_SL g5741 ( 
.A(n_5732),
.Y(n_5741)
);

INVx1_ASAP7_75t_L g5742 ( 
.A(n_5735),
.Y(n_5742)
);

XNOR2xp5_ASAP7_75t_L g5743 ( 
.A(n_5734),
.B(n_515),
.Y(n_5743)
);

HB1xp67_ASAP7_75t_L g5744 ( 
.A(n_5736),
.Y(n_5744)
);

BUFx2_ASAP7_75t_L g5745 ( 
.A(n_5744),
.Y(n_5745)
);

XNOR2x1_ASAP7_75t_L g5746 ( 
.A(n_5742),
.B(n_5737),
.Y(n_5746)
);

O2A1O1Ixp33_ASAP7_75t_L g5747 ( 
.A1(n_5741),
.A2(n_516),
.B(n_517),
.C(n_518),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_5743),
.Y(n_5748)
);

NAND2xp5_ASAP7_75t_SL g5749 ( 
.A(n_5740),
.B(n_519),
.Y(n_5749)
);

NAND4xp75_ASAP7_75t_L g5750 ( 
.A(n_5748),
.B(n_5739),
.C(n_521),
.D(n_522),
.Y(n_5750)
);

NAND4xp75_ASAP7_75t_L g5751 ( 
.A(n_5749),
.B(n_520),
.C(n_521),
.D(n_523),
.Y(n_5751)
);

NOR2x1_ASAP7_75t_L g5752 ( 
.A(n_5745),
.B(n_520),
.Y(n_5752)
);

INVx2_ASAP7_75t_L g5753 ( 
.A(n_5746),
.Y(n_5753)
);

AOI31xp33_ASAP7_75t_L g5754 ( 
.A1(n_5753),
.A2(n_5747),
.A3(n_525),
.B(n_526),
.Y(n_5754)
);

AOI22xp33_ASAP7_75t_L g5755 ( 
.A1(n_5752),
.A2(n_523),
.B1(n_525),
.B2(n_526),
.Y(n_5755)
);

AOI22xp33_ASAP7_75t_L g5756 ( 
.A1(n_5750),
.A2(n_5751),
.B1(n_528),
.B2(n_529),
.Y(n_5756)
);

OAI22xp5_ASAP7_75t_SL g5757 ( 
.A1(n_5753),
.A2(n_527),
.B1(n_529),
.B2(n_530),
.Y(n_5757)
);

AOI31xp33_ASAP7_75t_L g5758 ( 
.A1(n_5753),
.A2(n_530),
.A3(n_531),
.B(n_532),
.Y(n_5758)
);

AOI22xp5_ASAP7_75t_L g5759 ( 
.A1(n_5756),
.A2(n_534),
.B1(n_535),
.B2(n_536),
.Y(n_5759)
);

OAI311xp33_ASAP7_75t_L g5760 ( 
.A1(n_5754),
.A2(n_534),
.A3(n_537),
.B1(n_541),
.C1(n_542),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5757),
.Y(n_5761)
);

INVx1_ASAP7_75t_L g5762 ( 
.A(n_5758),
.Y(n_5762)
);

OAI22xp5_ASAP7_75t_L g5763 ( 
.A1(n_5755),
.A2(n_537),
.B1(n_542),
.B2(n_543),
.Y(n_5763)
);

INVx1_ASAP7_75t_L g5764 ( 
.A(n_5754),
.Y(n_5764)
);

INVx2_ASAP7_75t_L g5765 ( 
.A(n_5757),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5754),
.Y(n_5766)
);

INVx1_ASAP7_75t_L g5767 ( 
.A(n_5754),
.Y(n_5767)
);

XNOR2xp5_ASAP7_75t_L g5768 ( 
.A(n_5756),
.B(n_543),
.Y(n_5768)
);

OAI21xp33_ASAP7_75t_L g5769 ( 
.A1(n_5759),
.A2(n_544),
.B(n_545),
.Y(n_5769)
);

OR2x2_ASAP7_75t_L g5770 ( 
.A(n_5763),
.B(n_544),
.Y(n_5770)
);

INVx2_ASAP7_75t_L g5771 ( 
.A(n_5768),
.Y(n_5771)
);

AOI21xp5_ASAP7_75t_L g5772 ( 
.A1(n_5761),
.A2(n_545),
.B(n_546),
.Y(n_5772)
);

AOI21xp5_ASAP7_75t_L g5773 ( 
.A1(n_5762),
.A2(n_546),
.B(n_547),
.Y(n_5773)
);

OAI22x1_ASAP7_75t_L g5774 ( 
.A1(n_5765),
.A2(n_549),
.B1(n_552),
.B2(n_554),
.Y(n_5774)
);

HB1xp67_ASAP7_75t_L g5775 ( 
.A(n_5764),
.Y(n_5775)
);

NAND2xp5_ASAP7_75t_L g5776 ( 
.A(n_5766),
.B(n_549),
.Y(n_5776)
);

AOI21xp33_ASAP7_75t_SL g5777 ( 
.A1(n_5767),
.A2(n_552),
.B(n_554),
.Y(n_5777)
);

AOI22xp5_ASAP7_75t_L g5778 ( 
.A1(n_5760),
.A2(n_557),
.B1(n_558),
.B2(n_559),
.Y(n_5778)
);

OAI22xp33_ASAP7_75t_SL g5779 ( 
.A1(n_5770),
.A2(n_557),
.B1(n_558),
.B2(n_559),
.Y(n_5779)
);

AOI22xp33_ASAP7_75t_L g5780 ( 
.A1(n_5769),
.A2(n_5775),
.B1(n_5771),
.B2(n_5778),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5773),
.Y(n_5781)
);

AOI22xp33_ASAP7_75t_R g5782 ( 
.A1(n_5777),
.A2(n_560),
.B1(n_561),
.B2(n_563),
.Y(n_5782)
);

AOI222xp33_ASAP7_75t_L g5783 ( 
.A1(n_5774),
.A2(n_561),
.B1(n_563),
.B2(n_564),
.C1(n_565),
.C2(n_566),
.Y(n_5783)
);

OAI222xp33_ASAP7_75t_L g5784 ( 
.A1(n_5781),
.A2(n_5772),
.B1(n_5776),
.B2(n_567),
.C1(n_569),
.C2(n_572),
.Y(n_5784)
);

XNOR2xp5_ASAP7_75t_L g5785 ( 
.A(n_5780),
.B(n_590),
.Y(n_5785)
);

INVx3_ASAP7_75t_L g5786 ( 
.A(n_5782),
.Y(n_5786)
);

OR2x2_ASAP7_75t_L g5787 ( 
.A(n_5783),
.B(n_564),
.Y(n_5787)
);

AOI22xp5_ASAP7_75t_L g5788 ( 
.A1(n_5786),
.A2(n_5779),
.B1(n_567),
.B2(n_574),
.Y(n_5788)
);

AOI22x1_ASAP7_75t_L g5789 ( 
.A1(n_5787),
.A2(n_565),
.B1(n_574),
.B2(n_575),
.Y(n_5789)
);

AOI221xp5_ASAP7_75t_L g5790 ( 
.A1(n_5788),
.A2(n_5784),
.B1(n_5785),
.B2(n_577),
.C(n_578),
.Y(n_5790)
);

AOI22xp33_ASAP7_75t_L g5791 ( 
.A1(n_5790),
.A2(n_5789),
.B1(n_576),
.B2(n_577),
.Y(n_5791)
);

AOI211xp5_ASAP7_75t_L g5792 ( 
.A1(n_5791),
.A2(n_575),
.B(n_576),
.C(n_578),
.Y(n_5792)
);


endmodule