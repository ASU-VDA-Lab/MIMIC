module real_jpeg_31936_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_0),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_0),
.Y(n_314)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_0),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_60),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_1),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_1),
.B(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_1),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_1),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_1),
.B(n_433),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_1),
.Y(n_456)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_2),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_2),
.B(n_263),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_2),
.B(n_449),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g479 ( 
.A(n_2),
.B(n_480),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_19),
.B(n_538),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_3),
.B(n_539),
.Y(n_538)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_4),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_4),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_4),
.B(n_260),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_4),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_4),
.B(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_8),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_9),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_9),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_9),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_9),
.B(n_128),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_9),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_9),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_10),
.B(n_263),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_10),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_10),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g447 ( 
.A(n_10),
.B(n_200),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_10),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_10),
.B(n_491),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_11),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_11),
.Y(n_143)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_12),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_14),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_15),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_15),
.A2(n_124),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_15),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_15),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_15),
.B(n_359),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_15),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_15),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_15),
.B(n_496),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_16),
.Y(n_165)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_17),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_17),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_17),
.B(n_117),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_17),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_17),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_17),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_169),
.B1(n_536),
.B2(n_537),
.Y(n_19)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_20),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_168),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_105),
.Y(n_22)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_23),
.B(n_105),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_88),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_55),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.C(n_49),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.C(n_36),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_27),
.A2(n_28),
.B1(n_32),
.B2(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_27),
.B(n_115),
.C(n_119),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_28),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_27),
.A2(n_28),
.B1(n_273),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_28),
.B(n_273),
.C(n_276),
.Y(n_272)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_31),
.Y(n_159)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_31),
.Y(n_200)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_32),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_36),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_36),
.A2(n_63),
.B1(n_70),
.B2(n_71),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_36),
.A2(n_63),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_36),
.A2(n_63),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_38),
.Y(n_240)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_40),
.B(n_49),
.Y(n_91)
);

NOR2xp67_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_47),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_48),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_50),
.B(n_94),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_50),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_53),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_54),
.Y(n_242)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_54),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_75),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.C(n_70),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_63),
.B(n_259),
.C(n_262),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_119),
.C(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_66),
.B(n_140),
.Y(n_194)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_68),
.Y(n_327)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_71),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_70),
.A2(n_71),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_71),
.Y(n_231)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_74),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_123),
.C(n_127),
.Y(n_122)
);

XOR2x2_ASAP7_75t_L g144 ( 
.A(n_77),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_80),
.Y(n_295)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_83),
.B(n_198),
.C(n_201),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_84),
.B(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_103),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_103),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_100),
.Y(n_92)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_97),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_97),
.B(n_154),
.C(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_97),
.B(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_99),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_99),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_100),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.C(n_130),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_109),
.Y(n_206)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_122),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_114),
.B(n_122),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_116),
.B1(n_119),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_119),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_119),
.B(n_232),
.Y(n_317)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_121),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_121),
.Y(n_431)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_121),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_127),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_127),
.A2(n_146),
.B1(n_217),
.B2(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_131),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_148),
.C(n_152),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.C(n_144),
.Y(n_132)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_133),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OA21x2_ASAP7_75t_L g435 ( 
.A1(n_136),
.A2(n_232),
.B(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_136),
.B(n_232),
.Y(n_436)
);

OAI21xp33_ASAP7_75t_L g467 ( 
.A1(n_136),
.A2(n_232),
.B(n_436),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_137),
.A2(n_138),
.B1(n_144),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_143),
.Y(n_366)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_144),
.Y(n_250)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_152),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_161),
.C(n_166),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_156),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_154),
.B(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_154),
.B(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_154),
.B(n_429),
.Y(n_463)
);

INVx8_ASAP7_75t_L g505 ( 
.A(n_155),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_157),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_157),
.B(n_330),
.C(n_335),
.Y(n_344)
);

OR2x2_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_180),
.C(n_183),
.Y(n_179)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_166),
.A2(n_183),
.B1(n_184),
.B2(n_191),
.Y(n_244)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_169),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_251),
.B(n_533),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_207),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_171),
.A2(n_534),
.B(n_535),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_204),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_172),
.B(n_204),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_R g172 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_187),
.C(n_192),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_188),
.B1(n_189),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_181),
.B(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_181),
.B(n_266),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_182),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_182),
.Y(n_498)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_246),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_193),
.B(n_197),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_195),
.B(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_202),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_208),
.B(n_210),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_245),
.C(n_248),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g400 ( 
.A(n_211),
.B(n_401),
.Y(n_400)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_229),
.C(n_243),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_212),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_226),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g384 ( 
.A(n_213),
.B(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_215),
.A2(n_216),
.B1(n_226),
.B2(n_227),
.Y(n_385)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_222),
.Y(n_216)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_217),
.Y(n_343)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_222),
.Y(n_341)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_229),
.B(n_243),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.C(n_241),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_230),
.B(n_381),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.C(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_285)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_234),
.Y(n_493)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_237),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_241),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_245),
.B(n_248),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_413),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_387),
.B(n_409),
.Y(n_252)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_369),
.B(n_386),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_345),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_255),
.B(n_345),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_305),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_256),
.B(n_306),
.C(n_337),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_282),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_257),
.B(n_283),
.C(n_286),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.C(n_271),
.Y(n_257)
);

XOR2x2_ASAP7_75t_L g367 ( 
.A(n_258),
.B(n_368),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_265),
.B(n_272),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_270),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_270),
.B(n_431),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_270),
.B(n_508),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_273),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_275),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_276),
.B(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_279),
.Y(n_445)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_281),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_297),
.B2(n_304),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_294),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_289),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_291),
.Y(n_484)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g434 ( 
.A(n_292),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_293),
.Y(n_511)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_294),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_297),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g377 ( 
.A(n_297),
.B(n_378),
.C(n_379),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_299),
.Y(n_457)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

OA21x2_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_308),
.B(n_312),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_337),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_315),
.C(n_328),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_328),
.Y(n_347)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx4f_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_315),
.B(n_347),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.C(n_323),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_316),
.A2(n_317),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_318),
.A2(n_319),
.B1(n_323),
.B2(n_324),
.Y(n_425)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

XNOR2x2_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_335),
.Y(n_328)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XOR2x2_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_344),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_340),
.C(n_344),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJx2_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.C(n_367),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_346),
.B(n_417),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_349),
.B(n_367),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.C(n_355),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_354),
.A2(n_355),
.B1(n_356),
.B2(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_354),
.Y(n_422)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.C(n_364),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_357),
.A2(n_358),
.B1(n_362),
.B2(n_363),
.Y(n_471)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_364),
.B(n_471),
.Y(n_470)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_370),
.B(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_372),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_384),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_383),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_380),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_395),
.C(n_396),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_383),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_407),
.C(n_408),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_SL g413 ( 
.A(n_387),
.B(n_414),
.C(n_531),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_399),
.B1(n_402),
.B2(n_405),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_400),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_400),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.C(n_397),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_397),
.Y(n_404)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_406),
.Y(n_411)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_411),
.B(n_412),
.Y(n_409)
);

AO21x2_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_437),
.B(n_530),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_416),
.B(n_418),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.C(n_426),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_419),
.A2(n_420),
.B1(n_528),
.B2(n_529),
.Y(n_527)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_420),
.B(n_524),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_423),
.B(n_426),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_423),
.B(n_426),
.Y(n_529)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.C(n_435),
.Y(n_426)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_466),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_435),
.B1(n_467),
.B2(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_432),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_522),
.B(n_526),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_473),
.B(n_521),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_464),
.Y(n_439)
);

NOR2x1_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_464),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_453),
.C(n_463),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_442),
.B(n_518),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_447),
.C(n_452),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_503),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_447),
.A2(n_448),
.B1(n_451),
.B2(n_452),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_447),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_448),
.Y(n_452)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AO22x1_ASAP7_75t_L g518 ( 
.A1(n_453),
.A2(n_454),
.B1(n_463),
.B2(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_458),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_455),
.A2(n_458),
.B1(n_459),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_455),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx4_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_463),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_469),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_465),
.B(n_470),
.C(n_472),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_474),
.A2(n_515),
.B(n_520),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_499),
.B(n_514),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_488),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_476),
.B(n_488),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_478),
.B1(n_485),
.B2(n_486),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_479),
.B(n_482),
.C(n_485),
.Y(n_516)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_494),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_489),
.A2(n_490),
.B1(n_494),
.B2(n_495),
.Y(n_512)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx3_ASAP7_75t_SL g491 ( 
.A(n_492),
.Y(n_491)
);

INVx8_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_506),
.B(n_513),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx5_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_512),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_512),
.Y(n_513)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_517),
.Y(n_520)
);

NOR2x1p5_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule