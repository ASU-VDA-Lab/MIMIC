module fake_jpeg_2019_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_8),
.B(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_28),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_4),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_18),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_20),
.B1(n_14),
.B2(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_26),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_22),
.C(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_26),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_23),
.A2(n_15),
.B1(n_12),
.B2(n_9),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_30),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_9),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_11),
.Y(n_48)
);

A2O1A1O1Ixp25_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_49),
.B(n_50),
.C(n_16),
.D(n_12),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_16),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_37),
.B(n_32),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_51),
.B(n_28),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_58),
.C(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_57),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_30),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_56),
.C(n_38),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_45),
.B1(n_42),
.B2(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_1),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_53),
.B(n_54),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_60),
.B(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

BUFx12f_ASAP7_75t_SL g71 ( 
.A(n_68),
.Y(n_71)
);

AO221x1_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_38),
.B1(n_21),
.B2(n_3),
.C(n_2),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_71),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_73),
.B(n_70),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_72),
.C(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_7),
.B1(n_4),
.B2(n_3),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_3),
.Y(n_77)
);


endmodule