module fake_jpeg_11398_n_61 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_61);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_32),
.B1(n_17),
.B2(n_19),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_20),
.A2(n_24),
.B1(n_17),
.B2(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_30),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_22),
.B1(n_18),
.B2(n_7),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_41),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_37),
.B(n_33),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_42),
.B(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_5),
.Y(n_42)
);

OA21x2_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_5),
.B(n_6),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_22),
.B(n_18),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_10),
.C(n_11),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_48),
.B(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_46),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_55),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_47),
.B(n_51),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_57),
.B(n_52),
.Y(n_59)
);

XNOR2x1_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_46),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_58),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);


endmodule