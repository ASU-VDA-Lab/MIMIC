module fake_netlist_6_4168_n_845 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_845);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_845;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_41),
.Y(n_184)
);

INVxp33_ASAP7_75t_SL g185 ( 
.A(n_98),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_50),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_33),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_25),
.Y(n_191)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_128),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_3),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_149),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_139),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_12),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_133),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_116),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_110),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_71),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_24),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_46),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_106),
.Y(n_210)
);

BUFx2_ASAP7_75t_SL g211 ( 
.A(n_72),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_97),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_70),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_26),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_40),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_45),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_95),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_39),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_0),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_131),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_16),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_115),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_34),
.B(n_93),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_59),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_163),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_19),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_62),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_29),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_11),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_86),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_27),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_63),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_68),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_182),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_177),
.Y(n_253)
);

OA21x2_ASAP7_75t_L g254 ( 
.A1(n_227),
.A2(n_1),
.B(n_2),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_193),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_196),
.B(n_3),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_178),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

OA21x2_ASAP7_75t_L g264 ( 
.A1(n_184),
.A2(n_4),
.B(n_5),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_188),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_187),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

AOI22x1_ASAP7_75t_SL g272 ( 
.A1(n_224),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

AOI22x1_ASAP7_75t_SL g274 ( 
.A1(n_201),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_222),
.B(n_8),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_222),
.Y(n_277)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_205),
.B(n_20),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_179),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_214),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_204),
.B(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_211),
.Y(n_285)
);

OAI22x1_ASAP7_75t_R g286 ( 
.A1(n_214),
.A2(n_179),
.B1(n_186),
.B2(n_203),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_216),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_238),
.B(n_9),
.Y(n_289)
);

AOI22x1_ASAP7_75t_SL g290 ( 
.A1(n_186),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_280),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_L g295 ( 
.A1(n_258),
.A2(n_245),
.B1(n_276),
.B2(n_256),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_217),
.Y(n_297)
);

OR2x6_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_226),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_250),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_250),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_247),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_250),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_250),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_242),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_208),
.C(n_203),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_244),
.B(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_285),
.B(n_218),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_289),
.B(n_185),
.Y(n_314)
);

INVxp33_ASAP7_75t_SL g315 ( 
.A(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g319 ( 
.A1(n_256),
.A2(n_277),
.B1(n_271),
.B2(n_254),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_242),
.Y(n_320)
);

AND3x2_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_228),
.C(n_235),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

NOR2x1p5_ASAP7_75t_L g324 ( 
.A(n_246),
.B(n_208),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_248),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_252),
.B(n_185),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_248),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_244),
.B(n_225),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_261),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_275),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_261),
.Y(n_336)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_220),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_225),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_314),
.A2(n_278),
.B1(n_231),
.B2(n_219),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_278),
.B1(n_231),
.B2(n_241),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_293),
.B(n_285),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_301),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_333),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_295),
.B(n_190),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_324),
.Y(n_351)
);

INVxp33_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_342),
.B(n_269),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_296),
.B(n_300),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_243),
.C(n_192),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_293),
.B(n_253),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_323),
.Y(n_357)
);

BUFx6f_ASAP7_75t_SL g358 ( 
.A(n_298),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_331),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_309),
.B(n_191),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_SL g365 ( 
.A(n_306),
.B(n_269),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_309),
.B(n_195),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_323),
.B(n_269),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_319),
.B(n_197),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_263),
.Y(n_371)
);

OAI21xp33_ASAP7_75t_L g372 ( 
.A1(n_329),
.A2(n_268),
.B(n_265),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_310),
.B(n_273),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_306),
.Y(n_374)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_283),
.C(n_279),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_312),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_297),
.B(n_261),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_262),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_315),
.B(n_210),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_341),
.A2(n_288),
.B(n_287),
.C(n_266),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_305),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_311),
.A2(n_259),
.B(n_255),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_338),
.B(n_262),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_315),
.B(n_212),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_261),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_339),
.A2(n_264),
.B1(n_254),
.B2(n_278),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_305),
.B(n_317),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_302),
.B(n_215),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_SL g394 ( 
.A(n_340),
.B(n_281),
.Y(n_394)
);

NOR3xp33_ASAP7_75t_L g395 ( 
.A(n_340),
.B(n_270),
.C(n_262),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_334),
.B(n_221),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_298),
.B(n_279),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_305),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_291),
.B(n_267),
.Y(n_399)
);

NOR2xp67_ASAP7_75t_L g400 ( 
.A(n_294),
.B(n_270),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_317),
.B(n_270),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_318),
.B(n_267),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_298),
.B(n_287),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_298),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_291),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_320),
.Y(n_406)
);

INVx2_ASAP7_75t_SL g407 ( 
.A(n_292),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_334),
.B(n_223),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_320),
.B(n_267),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_292),
.B(n_288),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_334),
.B(n_255),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_354),
.A2(n_337),
.B(n_294),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_278),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_359),
.B(n_229),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_369),
.B(n_346),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_356),
.A2(n_230),
.B(n_232),
.C(n_260),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_390),
.A2(n_345),
.B(n_344),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_281),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_397),
.B(n_267),
.Y(n_420)
);

INVx11_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_278),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_322),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_410),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_390),
.B(n_322),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_357),
.A2(n_337),
.B(n_294),
.Y(n_429)
);

A2O1A1Ixp33_ASAP7_75t_L g430 ( 
.A1(n_372),
.A2(n_260),
.B(n_259),
.C(n_275),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_325),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_349),
.B(n_351),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_350),
.A2(n_264),
.B(n_254),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_362),
.B(n_284),
.Y(n_434)
);

AOI21xp33_ASAP7_75t_L g435 ( 
.A1(n_370),
.A2(n_264),
.B(n_286),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_325),
.B(n_327),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_379),
.B(n_327),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_366),
.B(n_290),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_21),
.Y(n_439)
);

AOI21xp33_ASAP7_75t_L g440 ( 
.A1(n_403),
.A2(n_10),
.B(n_13),
.Y(n_440)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_401),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_393),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_377),
.B(n_328),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_368),
.A2(n_337),
.B(n_335),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_347),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_348),
.B(n_328),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_360),
.B(n_330),
.Y(n_448)
);

O2A1O1Ixp33_ASAP7_75t_SL g449 ( 
.A1(n_396),
.A2(n_330),
.B(n_332),
.C(n_274),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_353),
.A2(n_337),
.B(n_335),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_361),
.B(n_332),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_364),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_367),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_391),
.A2(n_335),
.B(n_306),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_406),
.A2(n_335),
.B(n_306),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_376),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_363),
.B(n_275),
.Y(n_457)
);

O2A1O1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_384),
.A2(n_284),
.B(n_275),
.C(n_272),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_404),
.B(n_22),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_355),
.A2(n_284),
.B1(n_275),
.B2(n_335),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_284),
.C(n_306),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_378),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_374),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_23),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_408),
.A2(n_94),
.B(n_175),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_402),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_392),
.A2(n_92),
.B1(n_174),
.B2(n_173),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_358),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_28),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_411),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_374),
.B(n_30),
.Y(n_471)
);

OAI321xp33_ASAP7_75t_L g472 ( 
.A1(n_384),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_381),
.B(n_14),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_385),
.B(n_31),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_409),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_394),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_380),
.A2(n_373),
.B(n_371),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_400),
.A2(n_100),
.B(n_171),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_389),
.B(n_32),
.Y(n_481)
);

NAND2xp33_ASAP7_75t_L g482 ( 
.A(n_411),
.B(n_35),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g484 ( 
.A1(n_473),
.A2(n_355),
.B(n_388),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_416),
.B(n_442),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_427),
.A2(n_386),
.B(n_389),
.Y(n_486)
);

BUFx12f_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_443),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_418),
.A2(n_358),
.B1(n_386),
.B2(n_395),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_421),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_424),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_478),
.A2(n_399),
.B(n_365),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_431),
.A2(n_399),
.B(n_102),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_419),
.B(n_15),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_432),
.Y(n_495)
);

OAI21x1_ASAP7_75t_SL g496 ( 
.A1(n_413),
.A2(n_433),
.B(n_464),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_422),
.A2(n_101),
.B(n_170),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_437),
.A2(n_96),
.B(n_168),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_479),
.A2(n_176),
.B(n_91),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_470),
.A2(n_89),
.B(n_164),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_476),
.Y(n_501)
);

AO31x2_ASAP7_75t_L g502 ( 
.A1(n_430),
.A2(n_17),
.A3(n_18),
.B(n_19),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_470),
.A2(n_36),
.B(n_38),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_425),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_479),
.A2(n_42),
.B(n_43),
.Y(n_506)
);

OAI21xp33_ASAP7_75t_L g507 ( 
.A1(n_435),
.A2(n_44),
.B(n_47),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_466),
.B(n_434),
.Y(n_508)
);

AOI21x1_ASAP7_75t_L g509 ( 
.A1(n_451),
.A2(n_48),
.B(n_49),
.Y(n_509)
);

AO31x2_ASAP7_75t_L g510 ( 
.A1(n_417),
.A2(n_51),
.A3(n_52),
.B(n_53),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_475),
.B(n_54),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_438),
.B(n_56),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_475),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_436),
.A2(n_165),
.B(n_58),
.Y(n_514)
);

AOI211x1_ASAP7_75t_L g515 ( 
.A1(n_433),
.A2(n_57),
.B(n_60),
.C(n_61),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_436),
.A2(n_64),
.B(n_65),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_66),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_441),
.B(n_67),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_463),
.Y(n_519)
);

OAI21x1_ASAP7_75t_L g520 ( 
.A1(n_445),
.A2(n_69),
.B(n_73),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_450),
.A2(n_74),
.B(n_77),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_426),
.B(n_78),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_441),
.A2(n_79),
.B(n_80),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_457),
.A2(n_81),
.B(n_82),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_440),
.A2(n_83),
.B(n_84),
.C(n_85),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_428),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_461),
.A2(n_481),
.B(n_460),
.Y(n_527)
);

NOR4xp25_ASAP7_75t_L g528 ( 
.A(n_472),
.B(n_87),
.C(n_88),
.D(n_103),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_414),
.B(n_420),
.Y(n_529)
);

OA21x2_ASAP7_75t_L g530 ( 
.A1(n_454),
.A2(n_105),
.B(n_107),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_463),
.A2(n_471),
.B(n_455),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_460),
.B(n_108),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_459),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_441),
.A2(n_474),
.B(n_467),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_461),
.A2(n_472),
.B(n_412),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_448),
.A2(n_161),
.B(n_119),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_423),
.B(n_114),
.Y(n_537)
);

AO31x2_ASAP7_75t_L g538 ( 
.A1(n_480),
.A2(n_120),
.A3(n_121),
.B(n_123),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_458),
.B(n_124),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_456),
.B(n_127),
.Y(n_540)
);

OAI21x1_ASAP7_75t_SL g541 ( 
.A1(n_498),
.A2(n_465),
.B(n_444),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_485),
.A2(n_439),
.B1(n_446),
.B2(n_462),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_512),
.A2(n_453),
.B1(n_452),
.B2(n_477),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_484),
.A2(n_507),
.B1(n_532),
.B2(n_539),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_488),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_491),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_505),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_531),
.A2(n_456),
.B(n_429),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_486),
.A2(n_482),
.B(n_469),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_513),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_526),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

BUFx2_ASAP7_75t_SL g553 ( 
.A(n_490),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_492),
.A2(n_447),
.B(n_130),
.Y(n_554)
);

AO32x2_ASAP7_75t_L g555 ( 
.A1(n_489),
.A2(n_449),
.A3(n_447),
.B1(n_136),
.B2(n_138),
.Y(n_555)
);

A2O1A1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_484),
.A2(n_447),
.B(n_135),
.C(n_140),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_535),
.A2(n_447),
.B(n_142),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_508),
.B(n_129),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_513),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_519),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_496),
.A2(n_143),
.B(n_144),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_521),
.A2(n_145),
.B(n_146),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_519),
.Y(n_563)
);

AO31x2_ASAP7_75t_L g564 ( 
.A1(n_493),
.A2(n_147),
.A3(n_150),
.B(n_151),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_520),
.A2(n_506),
.B(n_499),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_501),
.B(n_152),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_501),
.B(n_154),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_511),
.A2(n_155),
.B(n_156),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_534),
.A2(n_158),
.B(n_159),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_513),
.B(n_160),
.Y(n_570)
);

NAND2x1p5_ASAP7_75t_L g571 ( 
.A(n_483),
.B(n_504),
.Y(n_571)
);

OA21x2_ASAP7_75t_L g572 ( 
.A1(n_527),
.A2(n_535),
.B(n_516),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_507),
.A2(n_494),
.B1(n_529),
.B2(n_483),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_517),
.A2(n_527),
.B(n_537),
.Y(n_574)
);

AO31x2_ASAP7_75t_L g575 ( 
.A1(n_525),
.A2(n_540),
.A3(n_522),
.B(n_533),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_514),
.A2(n_536),
.B(n_497),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_483),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_509),
.A2(n_500),
.B(n_503),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_510),
.B(n_538),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_515),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_528),
.B(n_515),
.Y(n_582)
);

INVx6_ASAP7_75t_L g583 ( 
.A(n_487),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_510),
.B(n_538),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_524),
.Y(n_585)
);

BUFx12f_ASAP7_75t_L g586 ( 
.A(n_502),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_518),
.A2(n_523),
.B(n_530),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_502),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_530),
.A2(n_524),
.B(n_510),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_538),
.B(n_490),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_513),
.B(n_483),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_580),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_551),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_588),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_544),
.B(n_573),
.Y(n_595)
);

CKINVDCx11_ASAP7_75t_R g596 ( 
.A(n_552),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_546),
.Y(n_597)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_565),
.A2(n_554),
.B(n_548),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_547),
.Y(n_599)
);

NAND2x1p5_ASAP7_75t_L g600 ( 
.A(n_561),
.B(n_568),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_560),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_563),
.Y(n_602)
);

OAI21x1_ASAP7_75t_SL g603 ( 
.A1(n_557),
.A2(n_549),
.B(n_569),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_550),
.B(n_559),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_555),
.B(n_557),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_566),
.A2(n_567),
.B1(n_583),
.B2(n_581),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_558),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_545),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_556),
.Y(n_611)
);

AOI21x1_ASAP7_75t_L g612 ( 
.A1(n_574),
.A2(n_587),
.B(n_589),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_555),
.B(n_572),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_562),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_581),
.A2(n_582),
.B1(n_586),
.B2(n_577),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_550),
.B(n_559),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_576),
.A2(n_549),
.B(n_587),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_571),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_591),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_579),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_579),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_555),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_582),
.B(n_590),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_590),
.B(n_584),
.Y(n_624)
);

OAI22xp5_ASAP7_75t_L g625 ( 
.A1(n_543),
.A2(n_542),
.B1(n_590),
.B2(n_585),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_570),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_584),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_542),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_543),
.A2(n_553),
.B1(n_578),
.B2(n_541),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_585),
.A2(n_578),
.B(n_575),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_564),
.B(n_575),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_564),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_564),
.B(n_575),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_583),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_545),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_623),
.B(n_594),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_607),
.B(n_605),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_592),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_592),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_610),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_623),
.B(n_602),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_605),
.B(n_609),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_627),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_599),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_620),
.B(n_621),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

AO31x2_ASAP7_75t_L g648 ( 
.A1(n_632),
.A2(n_625),
.A3(n_630),
.B(n_628),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_594),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_628),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_620),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_632),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_615),
.B(n_595),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_608),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_602),
.B(n_593),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_621),
.B(n_624),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_608),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_624),
.B(n_622),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_635),
.B(n_626),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_635),
.B(n_626),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_597),
.B(n_593),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_604),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_601),
.B(n_597),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_631),
.Y(n_664)
);

CKINVDCx11_ASAP7_75t_R g665 ( 
.A(n_604),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_631),
.Y(n_666)
);

OAI222xp33_ASAP7_75t_L g667 ( 
.A1(n_606),
.A2(n_611),
.B1(n_601),
.B2(n_622),
.C1(n_618),
.C2(n_629),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_604),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_627),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_627),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_604),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_619),
.B(n_634),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_616),
.B(n_611),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_633),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_606),
.B(n_613),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_613),
.B(n_627),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_612),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_616),
.B(n_617),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_612),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_614),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_616),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_617),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_616),
.B(n_600),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_600),
.B(n_598),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_600),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_603),
.Y(n_687)
);

INVxp67_ASAP7_75t_SL g688 ( 
.A(n_661),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_637),
.B(n_603),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_654),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_649),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_649),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_652),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_676),
.B(n_642),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_652),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_636),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_636),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_655),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_676),
.B(n_642),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_657),
.Y(n_700)
);

BUFx2_ASAP7_75t_L g701 ( 
.A(n_679),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_657),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_664),
.B(n_666),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_677),
.B(n_658),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_677),
.B(n_658),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_655),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_664),
.B(n_674),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_663),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_666),
.B(n_674),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_663),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_641),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_641),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_640),
.Y(n_713)
);

INVx4_ASAP7_75t_L g714 ( 
.A(n_665),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_643),
.B(n_660),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_659),
.B(n_668),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_653),
.A2(n_687),
.B1(n_656),
.B2(n_647),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_682),
.B(n_673),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_675),
.B(n_656),
.Y(n_719)
);

NAND2x1_ASAP7_75t_L g720 ( 
.A(n_644),
.B(n_685),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_675),
.B(n_648),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_645),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_648),
.B(n_687),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_648),
.B(n_687),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_645),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_638),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_646),
.Y(n_727)
);

INVx2_ASAP7_75t_SL g728 ( 
.A(n_656),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_650),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_715),
.B(n_653),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_701),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_701),
.B(n_679),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_704),
.B(n_705),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_693),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_704),
.B(n_648),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_695),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_713),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_691),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_705),
.B(n_648),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_694),
.B(n_656),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_700),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_L g742 ( 
.A(n_689),
.B(n_672),
.C(n_650),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_692),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_723),
.B(n_680),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_694),
.B(n_683),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_716),
.B(n_647),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_699),
.B(n_683),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_714),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_703),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_700),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_703),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_720),
.B(n_644),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_699),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_719),
.B(n_684),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_688),
.B(n_651),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_723),
.B(n_678),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_719),
.B(n_684),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_702),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_718),
.B(n_651),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_727),
.B(n_686),
.Y(n_760)
);

HB1xp67_ASAP7_75t_L g761 ( 
.A(n_698),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_724),
.B(n_680),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_735),
.B(n_724),
.Y(n_763)
);

INVxp33_ASAP7_75t_L g764 ( 
.A(n_746),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_735),
.B(n_721),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_737),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_734),
.Y(n_767)
);

OAI221xp5_ASAP7_75t_L g768 ( 
.A1(n_742),
.A2(n_717),
.B1(n_714),
.B2(n_647),
.C(n_697),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_748),
.B(n_714),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_739),
.B(n_721),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_739),
.B(n_709),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_731),
.B(n_696),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_730),
.B(n_706),
.Y(n_773)
);

AND2x6_ASAP7_75t_SL g774 ( 
.A(n_748),
.B(n_646),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_734),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_759),
.B(n_729),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_736),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_761),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_731),
.B(n_720),
.Y(n_779)
);

NAND2x1_ASAP7_75t_L g780 ( 
.A(n_760),
.B(n_727),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_763),
.B(n_753),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_767),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_773),
.B(n_733),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_775),
.Y(n_784)
);

AOI32xp33_ASAP7_75t_L g785 ( 
.A1(n_768),
.A2(n_732),
.A3(n_740),
.B1(n_733),
.B2(n_757),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_766),
.B(n_754),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_777),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_780),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_779),
.B(n_732),
.Y(n_789)
);

AOI21xp33_ASAP7_75t_L g790 ( 
.A1(n_764),
.A2(n_755),
.B(n_744),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_772),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_776),
.B(n_754),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_778),
.B(n_757),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_783),
.B(n_764),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_789),
.Y(n_795)
);

AOI211x1_ASAP7_75t_SL g796 ( 
.A1(n_790),
.A2(n_758),
.B(n_741),
.C(n_750),
.Y(n_796)
);

OAI21xp33_ASAP7_75t_L g797 ( 
.A1(n_785),
.A2(n_769),
.B(n_763),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_SL g798 ( 
.A1(n_788),
.A2(n_667),
.B(n_770),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_781),
.B(n_765),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_786),
.B(n_740),
.Y(n_800)
);

AOI21xp33_ASAP7_75t_L g801 ( 
.A1(n_787),
.A2(n_762),
.B(n_744),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_SL g802 ( 
.A(n_797),
.B(n_793),
.C(n_791),
.Y(n_802)
);

NAND2x1_ASAP7_75t_L g803 ( 
.A(n_795),
.B(n_788),
.Y(n_803)
);

AOI211xp5_ASAP7_75t_L g804 ( 
.A1(n_798),
.A2(n_782),
.B(n_784),
.C(n_792),
.Y(n_804)
);

NOR3x1_ASAP7_75t_L g805 ( 
.A(n_799),
.B(n_762),
.C(n_756),
.Y(n_805)
);

OAI211xp5_ASAP7_75t_SL g806 ( 
.A1(n_796),
.A2(n_743),
.B(n_738),
.C(n_749),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_794),
.B(n_789),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_807),
.B(n_800),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_804),
.B(n_801),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_805),
.B(n_802),
.Y(n_810)
);

NAND4xp25_ASAP7_75t_L g811 ( 
.A(n_806),
.B(n_662),
.C(n_756),
.D(n_765),
.Y(n_811)
);

NOR3x1_ASAP7_75t_L g812 ( 
.A(n_803),
.B(n_751),
.C(n_728),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_SL g813 ( 
.A(n_810),
.B(n_752),
.C(n_774),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_809),
.B(n_671),
.C(n_662),
.Y(n_814)
);

NAND4xp75_ASAP7_75t_L g815 ( 
.A(n_812),
.B(n_770),
.C(n_671),
.D(n_771),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_814),
.B(n_808),
.Y(n_816)
);

AND2x2_ASAP7_75t_SL g817 ( 
.A(n_813),
.B(n_811),
.Y(n_817)
);

NOR2x1_ASAP7_75t_L g818 ( 
.A(n_815),
.B(n_758),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_813),
.A2(n_752),
.B(n_711),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_817),
.A2(n_771),
.B1(n_747),
.B2(n_745),
.Y(n_820)
);

XOR2xp5_ASAP7_75t_L g821 ( 
.A(n_816),
.B(n_662),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_819),
.A2(n_760),
.B1(n_747),
.B2(n_745),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_818),
.Y(n_823)
);

NOR2x1_ASAP7_75t_L g824 ( 
.A(n_816),
.B(n_725),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_824),
.B(n_710),
.Y(n_825)
);

AOI211x1_ASAP7_75t_L g826 ( 
.A1(n_820),
.A2(n_708),
.B(n_707),
.C(n_709),
.Y(n_826)
);

NOR4xp25_ASAP7_75t_L g827 ( 
.A(n_823),
.B(n_722),
.C(n_712),
.D(n_741),
.Y(n_827)
);

NOR4xp25_ASAP7_75t_L g828 ( 
.A(n_821),
.B(n_822),
.C(n_750),
.D(n_702),
.Y(n_828)
);

AOI211xp5_ASAP7_75t_L g829 ( 
.A1(n_823),
.A2(n_760),
.B(n_707),
.C(n_646),
.Y(n_829)
);

CKINVDCx16_ASAP7_75t_R g830 ( 
.A(n_821),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_SL g831 ( 
.A1(n_825),
.A2(n_698),
.B(n_728),
.Y(n_831)
);

NAND4xp25_ASAP7_75t_L g832 ( 
.A(n_829),
.B(n_646),
.C(n_727),
.D(n_685),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_830),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_L g834 ( 
.A(n_826),
.B(n_670),
.C(n_669),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_833),
.B(n_828),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_831),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_832),
.B(n_827),
.C(n_670),
.Y(n_837)
);

AOI31xp33_ASAP7_75t_L g838 ( 
.A1(n_834),
.A2(n_669),
.A3(n_638),
.B(n_639),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_835),
.A2(n_726),
.B(n_639),
.Y(n_839)
);

XOR2x1_ASAP7_75t_L g840 ( 
.A(n_836),
.B(n_726),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_SL g841 ( 
.A1(n_837),
.A2(n_838),
.B1(n_644),
.B2(n_678),
.Y(n_841)
);

XNOR2xp5_ASAP7_75t_L g842 ( 
.A(n_840),
.B(n_841),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_842),
.B(n_839),
.Y(n_843)
);

NAND2x2_ASAP7_75t_L g844 ( 
.A(n_843),
.B(n_644),
.Y(n_844)
);

AOI21xp33_ASAP7_75t_SL g845 ( 
.A1(n_844),
.A2(n_681),
.B(n_690),
.Y(n_845)
);


endmodule