module real_aes_18267_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_844, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_844;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_635;
wire n_287;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g840 ( .A(n_0), .B(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_1), .A2(n_34), .B1(n_147), .B2(n_162), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_2), .A2(n_9), .B1(n_552), .B2(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g841 ( .A(n_3), .Y(n_841) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_4), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_5), .A2(n_10), .B1(n_563), .B2(n_564), .Y(n_562) );
OR2x2_ASAP7_75t_L g110 ( .A(n_6), .B(n_30), .Y(n_110) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_7), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g580 ( .A(n_8), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_11), .B(n_141), .Y(n_241) );
AOI22xp33_ASAP7_75t_SL g102 ( .A1(n_12), .A2(n_103), .B1(n_835), .B2(n_842), .Y(n_102) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_13), .A2(n_98), .B1(n_301), .B2(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_14), .A2(n_31), .B1(n_531), .B2(n_575), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g111 ( .A1(n_15), .A2(n_18), .B1(n_112), .B2(n_113), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_15), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_16), .B(n_141), .Y(n_528) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_17), .A2(n_46), .B(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g113 ( .A(n_18), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_19), .B(n_168), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_20), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_21), .A2(n_38), .B1(n_149), .B2(n_306), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_22), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_23), .A2(n_44), .B1(n_149), .B2(n_552), .Y(n_633) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_24), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_25), .B(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_26), .B(n_165), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g589 ( .A(n_27), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_28), .B(n_155), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_29), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_32), .A2(n_82), .B1(n_147), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_33), .A2(n_37), .B1(n_147), .B2(n_527), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_35), .A2(n_49), .B1(n_552), .B2(n_554), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_36), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_39), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g117 ( .A(n_40), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_41), .A2(n_52), .B1(n_493), .B2(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g494 ( .A(n_41), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_42), .B(n_150), .Y(n_160) );
BUFx3_ASAP7_75t_L g109 ( .A(n_43), .Y(n_109) );
INVx1_ASAP7_75t_L g502 ( .A(n_43), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_45), .B(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g226 ( .A(n_47), .B(n_172), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_48), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_50), .B(n_165), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_51), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g493 ( .A(n_52), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_53), .A2(n_69), .B1(n_306), .B2(n_554), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_54), .A2(n_72), .B1(n_147), .B2(n_527), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_55), .B(n_207), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_56), .A2(n_142), .B(n_218), .C(n_219), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_57), .A2(n_94), .B1(n_552), .B2(n_564), .Y(n_586) );
INVx1_ASAP7_75t_L g134 ( .A(n_58), .Y(n_134) );
AND2x4_ASAP7_75t_L g152 ( .A(n_59), .B(n_153), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_60), .A2(n_61), .B1(n_149), .B2(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_62), .B(n_155), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_63), .B(n_172), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_64), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_65), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g153 ( .A(n_66), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_67), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_68), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_70), .B(n_147), .Y(n_202) );
NAND3xp33_ASAP7_75t_L g161 ( .A(n_71), .B(n_150), .C(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_73), .B(n_147), .Y(n_233) );
INVx2_ASAP7_75t_L g144 ( .A(n_74), .Y(n_144) );
CKINVDCx14_ASAP7_75t_R g122 ( .A(n_75), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_75), .A2(n_122), .B1(n_492), .B2(n_495), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_76), .B(n_170), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_77), .B(n_141), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_78), .B(n_238), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_79), .A2(n_95), .B1(n_149), .B2(n_218), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_80), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_81), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_83), .A2(n_89), .B1(n_165), .B2(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g506 ( .A(n_84), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_85), .B(n_141), .Y(n_302) );
NAND2xp33_ASAP7_75t_SL g253 ( .A(n_86), .B(n_235), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_87), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_88), .B(n_155), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_90), .Y(n_569) );
INVx1_ASAP7_75t_L g485 ( .A(n_91), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_91), .B(n_501), .Y(n_500) );
NAND2xp33_ASAP7_75t_L g532 ( .A(n_92), .B(n_141), .Y(n_532) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_93), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_96), .B(n_172), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g249 ( .A(n_97), .B(n_170), .C(n_235), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_99), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_100), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_101), .B(n_165), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g103 ( .A(n_104), .B(n_508), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_118), .B(n_486), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AOI22x1_ASAP7_75t_L g508 ( .A1(n_106), .A2(n_509), .B1(n_831), .B2(n_833), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .C(n_114), .Y(n_106) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_107), .B(n_512), .Y(n_511) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g830 ( .A(n_108), .B(n_828), .Y(n_830) );
INVxp67_ASAP7_75t_L g838 ( .A(n_108), .Y(n_838) );
NOR2x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
INVx1_ASAP7_75t_L g503 ( .A(n_110), .Y(n_503) );
INVx1_ASAP7_75t_L g512 ( .A(n_111), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_114), .A2(n_487), .B(n_506), .Y(n_486) );
BUFx6f_ASAP7_75t_L g832 ( .A(n_114), .Y(n_832) );
CKINVDCx11_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_119), .A2(n_510), .B(n_829), .Y(n_509) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_481), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
BUFx2_ASAP7_75t_L g489 ( .A(n_123), .Y(n_489) );
NAND2x1p5_ASAP7_75t_SL g123 ( .A(n_124), .B(n_415), .Y(n_123) );
NOR2x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_351), .Y(n_124) );
NAND4xp25_ASAP7_75t_L g125 ( .A(n_126), .B(n_271), .C(n_312), .D(n_341), .Y(n_125) );
O2A1O1Ixp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_190), .B(n_197), .C(n_255), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_156), .Y(n_127) );
INVx2_ASAP7_75t_L g193 ( .A(n_128), .Y(n_193) );
AND2x2_ASAP7_75t_L g339 ( .A(n_128), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_128), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_128), .B(n_257), .Y(n_434) );
OR2x2_ASAP7_75t_L g470 ( .A(n_128), .B(n_386), .Y(n_470) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g367 ( .A(n_129), .B(n_157), .Y(n_367) );
NOR2xp67_ASAP7_75t_L g393 ( .A(n_129), .B(n_195), .Y(n_393) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g328 ( .A(n_130), .Y(n_328) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_135), .B(n_154), .Y(n_130) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_131), .A2(n_158), .B(n_171), .Y(n_157) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_131), .A2(n_135), .B(n_154), .Y(n_259) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_131), .A2(n_158), .B(n_171), .Y(n_294) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g155 ( .A(n_132), .Y(n_155) );
AND2x4_ASAP7_75t_SL g242 ( .A(n_132), .B(n_151), .Y(n_242) );
INVx1_ASAP7_75t_SL g245 ( .A(n_132), .Y(n_245) );
INVx2_ASAP7_75t_SL g523 ( .A(n_132), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_132), .B(n_543), .Y(n_542) );
BUFx3_ASAP7_75t_L g578 ( .A(n_132), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_132), .B(n_580), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_132), .B(n_589), .Y(n_588) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_145), .B(n_151), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_140), .B(n_142), .Y(n_136) );
INVx2_ASAP7_75t_L g301 ( .A(n_138), .Y(n_301) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_139), .Y(n_141) );
INVx3_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_139), .Y(n_162) );
INVx1_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
INVx2_ASAP7_75t_L g221 ( .A(n_139), .Y(n_221) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_139), .Y(n_235) );
INVx1_ASAP7_75t_L g252 ( .A(n_139), .Y(n_252) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g247 ( .A1(n_141), .A2(n_248), .B(n_249), .Y(n_247) );
INVx3_ASAP7_75t_L g552 ( .A(n_141), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_142), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_142), .A2(n_233), .B(n_234), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_142), .A2(n_251), .B(n_253), .Y(n_250) );
BUFx4f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx8_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx1_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
INVx2_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_150), .Y(n_145) );
OAI22xp33_ASAP7_75t_L g223 ( .A1(n_147), .A2(n_149), .B1(n_224), .B2(n_225), .Y(n_223) );
INVx4_ASAP7_75t_L g527 ( .A(n_147), .Y(n_527) );
INVx1_ASAP7_75t_L g554 ( .A(n_147), .Y(n_554) );
INVx1_ASAP7_75t_L g564 ( .A(n_147), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_149), .A2(n_160), .B(n_161), .Y(n_159) );
INVx2_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx6_ASAP7_75t_L g179 ( .A(n_150), .Y(n_179) );
O2A1O1Ixp5_ASAP7_75t_L g299 ( .A1(n_150), .A2(n_300), .B(n_301), .C(n_302), .Y(n_299) );
O2A1O1Ixp5_ASAP7_75t_L g525 ( .A1(n_150), .A2(n_526), .B(n_527), .C(n_528), .Y(n_525) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_151), .A2(n_159), .B(n_163), .Y(n_158) );
OAI21x1_ASAP7_75t_L g200 ( .A1(n_151), .A2(n_201), .B(n_204), .Y(n_200) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_151), .A2(n_247), .B(n_250), .Y(n_246) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_151), .A2(n_299), .B(n_303), .Y(n_298) );
BUFx10_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx10_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
INVx1_ASAP7_75t_L g534 ( .A(n_152), .Y(n_534) );
INVx2_ASAP7_75t_L g541 ( .A(n_155), .Y(n_541) );
AND2x2_ASAP7_75t_L g265 ( .A(n_156), .B(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_156), .B(n_295), .Y(n_311) );
AND2x2_ASAP7_75t_L g319 ( .A(n_156), .B(n_320), .Y(n_319) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_156), .Y(n_342) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_175), .Y(n_156) );
INVx1_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
INVx1_ASAP7_75t_L g257 ( .A(n_157), .Y(n_257) );
AND2x2_ASAP7_75t_L g329 ( .A(n_157), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g390 ( .A(n_157), .B(n_296), .Y(n_390) );
INVx2_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
AOI21x1_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_167), .B(n_169), .Y(n_163) );
INVx1_ASAP7_75t_L g563 ( .A(n_165), .Y(n_563) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_SL g566 ( .A(n_170), .Y(n_566) );
INVx1_ASAP7_75t_L g598 ( .A(n_170), .Y(n_598) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g209 ( .A(n_173), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_173), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_173), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g185 ( .A(n_174), .Y(n_185) );
INVx2_ASAP7_75t_L g189 ( .A(n_174), .Y(n_189) );
INVx1_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
AND2x2_ASAP7_75t_L g258 ( .A(n_175), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_175), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_175), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g373 ( .A(n_175), .B(n_328), .Y(n_373) );
OR2x2_ASAP7_75t_L g386 ( .A(n_175), .B(n_294), .Y(n_386) );
OR2x2_ASAP7_75t_L g396 ( .A(n_175), .B(n_259), .Y(n_396) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_185), .A3(n_186), .B(n_187), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_179), .B1(n_180), .B2(n_182), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_179), .A2(n_530), .B(n_532), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_179), .A2(n_182), .B1(n_539), .B2(n_540), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_179), .A2(n_182), .B1(n_551), .B2(n_553), .Y(n_550) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_179), .A2(n_562), .B1(n_565), .B2(n_566), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_179), .A2(n_182), .B1(n_574), .B2(n_576), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_179), .A2(n_566), .B1(n_586), .B2(n_587), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_179), .A2(n_595), .B1(n_597), .B2(n_598), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_179), .A2(n_182), .B1(n_632), .B2(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g577 ( .A(n_181), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_182), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g208 ( .A(n_183), .Y(n_208) );
BUFx3_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g239 ( .A(n_184), .Y(n_239) );
INVx2_ASAP7_75t_L g214 ( .A(n_185), .Y(n_214) );
NOR2xp33_ASAP7_75t_SL g568 ( .A(n_185), .B(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_185), .B(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g215 ( .A(n_186), .Y(n_215) );
AO31x2_ASAP7_75t_L g537 ( .A1(n_186), .A2(n_538), .A3(n_541), .B(n_542), .Y(n_537) );
AO31x2_ASAP7_75t_L g560 ( .A1(n_186), .A2(n_561), .A3(n_567), .B(n_568), .Y(n_560) );
AO31x2_ASAP7_75t_L g572 ( .A1(n_186), .A2(n_573), .A3(n_578), .B(n_579), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_189), .Y(n_187) );
BUFx2_ASAP7_75t_L g567 ( .A(n_189), .Y(n_567) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x4_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_193), .B(n_412), .Y(n_458) );
INVx1_ASAP7_75t_L g314 ( .A(n_194), .Y(n_314) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
AND2x2_ASAP7_75t_L g398 ( .A(n_196), .B(n_259), .Y(n_398) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_227), .Y(n_197) );
AND2x2_ASAP7_75t_L g269 ( .A(n_198), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g333 ( .A(n_198), .Y(n_333) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_211), .Y(n_198) );
BUFx2_ASAP7_75t_L g440 ( .A(n_199), .Y(n_440) );
OAI21xp33_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_209), .B(n_210), .Y(n_199) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_200), .A2(n_209), .B(n_210), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_208), .Y(n_204) );
OAI21x1_ASAP7_75t_L g297 ( .A1(n_209), .A2(n_298), .B(n_307), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_209), .A2(n_298), .B(n_307), .Y(n_330) );
AND2x2_ASAP7_75t_L g277 ( .A(n_211), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g263 ( .A(n_212), .B(n_244), .Y(n_263) );
INVx2_ASAP7_75t_L g289 ( .A(n_212), .Y(n_289) );
AOI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_226), .Y(n_212) );
NOR2xp67_ASAP7_75t_SL g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g555 ( .A(n_214), .Y(n_555) );
INVx1_ASAP7_75t_L g549 ( .A(n_215), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_217), .B(n_222), .Y(n_216) );
INVx1_ASAP7_75t_L g240 ( .A(n_218), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
INVx2_ASAP7_75t_SL g596 ( .A(n_221), .Y(n_596) );
AND2x2_ASAP7_75t_L g437 ( .A(n_227), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_243), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx4_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
BUFx2_ASAP7_75t_L g270 ( .A(n_229), .Y(n_270) );
OR2x2_ASAP7_75t_L g274 ( .A(n_229), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g336 ( .A(n_229), .B(n_278), .Y(n_336) );
AND2x4_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_236), .B(n_242), .Y(n_231) );
INVx2_ASAP7_75t_L g306 ( .A(n_235), .Y(n_306) );
INVx1_ASAP7_75t_L g531 ( .A(n_235), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B1(n_240), .B2(n_241), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_238), .A2(n_304), .B(n_305), .Y(n_303) );
INVx2_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g323 ( .A(n_243), .Y(n_323) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_243), .Y(n_337) );
INVx2_ASAP7_75t_L g362 ( .A(n_243), .Y(n_362) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g275 ( .A(n_244), .Y(n_275) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_254), .Y(n_244) );
INVx1_ASAP7_75t_L g575 ( .A(n_252), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_260), .B1(n_264), .B2(n_268), .Y(n_255) );
INVx1_ASAP7_75t_L g347 ( .A(n_256), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g358 ( .A(n_257), .Y(n_358) );
AND2x2_ASAP7_75t_L g375 ( .A(n_258), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_258), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g267 ( .A(n_259), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_260), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_263), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_261), .B(n_277), .Y(n_370) );
AND2x2_ASAP7_75t_L g378 ( .A(n_261), .B(n_344), .Y(n_378) );
AND2x2_ASAP7_75t_L g454 ( .A(n_261), .B(n_401), .Y(n_454) );
BUFx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g287 ( .A(n_262), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g310 ( .A(n_262), .B(n_278), .Y(n_310) );
OR2x2_ASAP7_75t_L g322 ( .A(n_262), .B(n_323), .Y(n_322) );
NAND2x1_ASAP7_75t_L g356 ( .A(n_262), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g361 ( .A(n_262), .Y(n_361) );
INVx2_ASAP7_75t_L g355 ( .A(n_263), .Y(n_355) );
AND2x2_ASAP7_75t_L g381 ( .A(n_263), .B(n_345), .Y(n_381) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
INVx1_ASAP7_75t_L g384 ( .A(n_266), .Y(n_384) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g368 ( .A(n_267), .B(n_296), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g379 ( .A1(n_268), .A2(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g441 ( .A(n_270), .B(n_381), .Y(n_441) );
INVx1_ASAP7_75t_L g477 ( .A(n_270), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_280), .B(n_284), .Y(n_271) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_272), .A2(n_321), .A3(n_426), .B1(n_427), .B2(n_428), .C1(n_429), .C2(n_432), .Y(n_425) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NOR3xp33_ASAP7_75t_L g413 ( .A(n_274), .B(n_276), .C(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g290 ( .A(n_275), .B(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g421 ( .A(n_275), .B(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_275), .Y(n_473) );
OR2x2_ASAP7_75t_L g369 ( .A(n_276), .B(n_322), .Y(n_369) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g357 ( .A(n_278), .Y(n_357) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_281), .Y(n_418) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g389 ( .A(n_282), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_283), .B(n_412), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_292), .B(n_308), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_286), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
AND2x2_ASAP7_75t_L g344 ( .A(n_288), .B(n_345), .Y(n_344) );
AND3x2_ASAP7_75t_L g388 ( .A(n_288), .B(n_290), .C(n_361), .Y(n_388) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g350 ( .A(n_289), .Y(n_350) );
AND2x2_ASAP7_75t_L g401 ( .A(n_289), .B(n_362), .Y(n_401) );
INVx2_ASAP7_75t_L g424 ( .A(n_289), .Y(n_424) );
AND2x2_ASAP7_75t_L g428 ( .A(n_290), .B(n_424), .Y(n_428) );
INVx2_ASAP7_75t_L g345 ( .A(n_291), .Y(n_345) );
OR2x2_ASAP7_75t_L g479 ( .A(n_291), .B(n_362), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_292), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g431 ( .A(n_293), .Y(n_431) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_330), .Y(n_340) );
AND2x2_ASAP7_75t_L g376 ( .A(n_294), .B(n_296), .Y(n_376) );
AND2x2_ASAP7_75t_L g372 ( .A(n_295), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_295), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g444 ( .A(n_295), .Y(n_444) );
BUFx3_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g315 ( .A(n_296), .Y(n_315) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_296), .Y(n_320) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_296), .Y(n_366) );
INVx1_ASAP7_75t_L g412 ( .A(n_296), .Y(n_412) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_321), .B(n_324), .Y(n_312) );
OAI31xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .A3(n_316), .B(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g395 ( .A(n_315), .Y(n_395) );
OAI32xp33_ASAP7_75t_L g353 ( .A1(n_316), .A2(n_325), .A3(n_354), .B1(n_358), .B2(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g346 ( .A(n_322), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_331), .B1(n_334), .B2(n_338), .Y(n_324) );
OAI22xp33_ASAP7_75t_SL g409 ( .A1(n_325), .A2(n_370), .B1(n_410), .B2(n_411), .Y(n_409) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
INVx2_ASAP7_75t_L g467 ( .A(n_327), .Y(n_467) );
BUFx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g422 ( .A(n_330), .Y(n_422) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g348 ( .A(n_336), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g423 ( .A(n_336), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g474 ( .A(n_336), .Y(n_474) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g414 ( .A(n_340), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_347), .B2(n_348), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_343), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AND2x2_ASAP7_75t_L g400 ( .A(n_345), .B(n_361), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_348), .A2(n_406), .B(n_409), .C(n_413), .Y(n_405) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_350), .Y(n_463) );
INVx1_ASAP7_75t_L g480 ( .A(n_350), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g351 ( .A(n_352), .B(n_374), .C(n_387), .D(n_405), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_353), .B(n_363), .Y(n_352) );
OR2x6_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_357), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g462 ( .A(n_360), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_369), .B1(n_370), .B2(n_371), .Y(n_363) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_365), .B(n_368), .Y(n_364) );
BUFx2_ASAP7_75t_L g377 ( .A(n_365), .Y(n_377) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_371), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g426 ( .A(n_373), .B(n_412), .Y(n_426) );
O2A1O1Ixp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_377), .B(n_378), .C(n_379), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_376), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g436 ( .A(n_383), .B(n_437), .Y(n_436) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_391), .B2(n_399), .C(n_402), .Y(n_387) );
AND2x2_ASAP7_75t_L g466 ( .A(n_390), .B(n_467), .Y(n_466) );
NAND3xp33_ASAP7_75t_SL g391 ( .A(n_392), .B(n_394), .C(n_397), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_395), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_395), .B(n_431), .Y(n_461) );
INVx1_ASAP7_75t_L g404 ( .A(n_396), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_396), .Y(n_408) );
AND2x2_ASAP7_75t_L g449 ( .A(n_398), .B(n_438), .Y(n_449) );
NAND2xp33_ASAP7_75t_SL g450 ( .A(n_398), .B(n_420), .Y(n_450) );
AND2x4_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_L g410 ( .A(n_401), .Y(n_410) );
NOR3x1_ASAP7_75t_L g415 ( .A(n_416), .B(n_445), .C(n_464), .Y(n_415) );
NAND3xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_425), .C(n_435), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g438 ( .A(n_422), .Y(n_438) );
INVx2_ASAP7_75t_L g427 ( .A(n_424), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_426), .A2(n_469), .B1(n_476), .B2(n_844), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g447 ( .A1(n_427), .A2(n_439), .B(n_448), .C(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AO21x1_ASAP7_75t_L g451 ( .A1(n_430), .A2(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g443 ( .A(n_434), .B(n_444), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B1(n_441), .B2(n_442), .Y(n_435) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND4xp75_ASAP7_75t_L g445 ( .A(n_446), .B(n_451), .C(n_455), .D(n_459), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_468), .C(n_475), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_471), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVxp67_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
AND2x4_ASAP7_75t_L g476 ( .A(n_477), .B(n_478), .Y(n_476) );
NOR2x1p5_ASAP7_75t_SL g478 ( .A(n_479), .B(n_480), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_482), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_484), .B(n_840), .Y(n_839) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g828 ( .A(n_485), .Y(n_828) );
OAI22xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B1(n_490), .B2(n_504), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g505 ( .A(n_491), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_492), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_496), .B(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g507 ( .A(n_499), .Y(n_507) );
AND2x6_ASAP7_75t_SL g499 ( .A(n_500), .B(n_503), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp33_ASAP7_75t_SL g510 ( .A(n_511), .B(n_513), .Y(n_510) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_513), .Y(n_834) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_514), .B(n_825), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_515), .B(n_769), .Y(n_514) );
NOR3x1_ASAP7_75t_L g515 ( .A(n_516), .B(n_687), .C(n_724), .Y(n_515) );
NAND4xp75_ASAP7_75t_L g516 ( .A(n_517), .B(n_607), .C(n_641), .D(n_671), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OAI32xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_544), .A3(n_581), .B1(n_590), .B2(n_602), .Y(n_518) );
OR2x2_ASAP7_75t_L g590 ( .A(n_519), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_520), .A2(n_799), .B(n_801), .Y(n_798) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_536), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_521), .B(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g670 ( .A(n_521), .B(n_616), .Y(n_670) );
AND2x2_ASAP7_75t_L g765 ( .A(n_521), .B(n_583), .Y(n_765) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx2_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
OAI21x1_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_535), .Y(n_522) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_523), .A2(n_524), .B(n_535), .Y(n_647) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_529), .B(n_533), .Y(n_524) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g599 ( .A(n_534), .Y(n_599) );
INVx2_ASAP7_75t_L g638 ( .A(n_536), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_536), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_537), .Y(n_625) );
INVx1_ASAP7_75t_L g669 ( .A(n_537), .Y(n_669) );
AND2x2_ASAP7_75t_L g713 ( .A(n_537), .B(n_647), .Y(n_713) );
OR2x2_ASAP7_75t_L g767 ( .A(n_537), .B(n_593), .Y(n_767) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_545), .A2(n_693), .B1(n_785), .B2(n_787), .Y(n_784) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
INVx4_ASAP7_75t_L g610 ( .A(n_546), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_546), .A2(n_592), .B1(n_622), .B2(n_624), .Y(n_621) );
OR2x2_ASAP7_75t_L g627 ( .A(n_546), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g746 ( .A(n_546), .B(n_645), .Y(n_746) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g666 ( .A(n_547), .B(n_559), .Y(n_666) );
AND2x2_ASAP7_75t_L g757 ( .A(n_547), .B(n_629), .Y(n_757) );
AND2x2_ASAP7_75t_L g812 ( .A(n_547), .B(n_572), .Y(n_812) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g606 ( .A(n_548), .Y(n_606) );
AND2x4_ASAP7_75t_L g733 ( .A(n_548), .B(n_629), .Y(n_733) );
AO31x2_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .A3(n_555), .B(n_556), .Y(n_548) );
AO31x2_ASAP7_75t_L g584 ( .A1(n_549), .A2(n_567), .A3(n_585), .B(n_588), .Y(n_584) );
AO31x2_ASAP7_75t_L g630 ( .A1(n_555), .A2(n_599), .A3(n_631), .B(n_634), .Y(n_630) );
NAND2x1_ASAP7_75t_L g609 ( .A(n_558), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_558), .B(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g558 ( .A(n_559), .B(n_570), .Y(n_558) );
INVx2_ASAP7_75t_L g604 ( .A(n_559), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_559), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g652 ( .A(n_559), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_559), .B(n_654), .Y(n_679) );
AND2x2_ASAP7_75t_L g682 ( .A(n_559), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g742 ( .A(n_559), .Y(n_742) );
INVx4_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_560), .B(n_571), .Y(n_620) );
BUFx2_ASAP7_75t_L g658 ( .A(n_560), .Y(n_658) );
AND2x2_ASAP7_75t_L g707 ( .A(n_560), .B(n_572), .Y(n_707) );
AND2x2_ASAP7_75t_L g749 ( .A(n_560), .B(n_630), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_560), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_572), .B(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g660 ( .A(n_572), .B(n_630), .Y(n_660) );
INVx1_ASAP7_75t_L g683 ( .A(n_572), .Y(n_683) );
INVx2_ASAP7_75t_L g703 ( .A(n_572), .Y(n_703) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_572), .Y(n_748) );
AO31x2_ASAP7_75t_L g593 ( .A1(n_578), .A2(n_594), .A3(n_599), .B(n_600), .Y(n_593) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g667 ( .A(n_582), .B(n_668), .Y(n_667) );
NOR2x1p5_ASAP7_75t_L g773 ( .A(n_582), .B(n_767), .Y(n_773) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g592 ( .A(n_583), .B(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g623 ( .A(n_583), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_583), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_583), .B(n_699), .Y(n_698) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g615 ( .A(n_584), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g673 ( .A(n_584), .B(n_593), .Y(n_673) );
BUFx2_ASAP7_75t_L g786 ( .A(n_584), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_590), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g824 ( .A(n_590), .Y(n_824) );
INVx2_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g760 ( .A(n_592), .Y(n_760) );
AND2x4_ASAP7_75t_L g783 ( .A(n_592), .B(n_713), .Y(n_783) );
AND2x2_ASAP7_75t_L g807 ( .A(n_592), .B(n_808), .Y(n_807) );
INVx2_ASAP7_75t_L g616 ( .A(n_593), .Y(n_616) );
BUFx2_ASAP7_75t_L g640 ( .A(n_593), .Y(n_640) );
INVx1_ASAP7_75t_L g696 ( .A(n_593), .Y(n_696) );
OR2x2_ASAP7_75t_L g818 ( .A(n_593), .B(n_675), .Y(n_818) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g664 ( .A(n_604), .Y(n_664) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_605), .Y(n_681) );
INVx1_ASAP7_75t_L g685 ( .A(n_605), .Y(n_685) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g626 ( .A(n_606), .Y(n_626) );
OR2x2_ASAP7_75t_L g663 ( .A(n_606), .B(n_655), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B(n_617), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_612), .A2(n_706), .B1(n_708), .B2(n_711), .Y(n_705) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
OR2x2_ASAP7_75t_L g751 ( .A(n_614), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g759 ( .A(n_614), .Y(n_759) );
AND2x2_ASAP7_75t_L g772 ( .A(n_614), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g734 ( .A(n_615), .B(n_713), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B1(n_627), .B2(n_636), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g686 ( .A(n_620), .Y(n_686) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g644 ( .A(n_623), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g712 ( .A(n_623), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g721 ( .A(n_623), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_623), .B(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_624), .B(n_793), .Y(n_792) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g709 ( .A(n_626), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g723 ( .A(n_626), .Y(n_723) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g655 ( .A(n_630), .Y(n_655) );
AND2x4_ASAP7_75t_L g702 ( .A(n_630), .B(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_630), .Y(n_718) );
INVx1_ASAP7_75t_L g782 ( .A(n_630), .Y(n_782) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AND2x4_ASAP7_75t_L g674 ( .A(n_638), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g691 ( .A(n_638), .Y(n_691) );
INVx1_ASAP7_75t_L g649 ( .A(n_640), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_650), .B1(n_661), .B2(n_667), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_644), .B(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_646), .Y(n_699) );
INVx1_ASAP7_75t_L g675 ( .A(n_647), .Y(n_675) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_651), .B(n_656), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_652), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g804 ( .A(n_653), .Y(n_804) );
INVx1_ASAP7_75t_L g823 ( .A(n_653), .Y(n_823) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NAND2x1_ASAP7_75t_L g800 ( .A(n_657), .B(n_723), .Y(n_800) );
AND2x4_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g816 ( .A(n_658), .Y(n_816) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
INVx2_ASAP7_75t_L g754 ( .A(n_662), .Y(n_754) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx2_ASAP7_75t_L g743 ( .A(n_663), .Y(n_743) );
AND2x4_ASAP7_75t_L g745 ( .A(n_664), .B(n_702), .Y(n_745) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_668), .A2(n_814), .B1(n_817), .B2(n_819), .Y(n_813) );
AND2x4_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g738 ( .A(n_669), .Y(n_738) );
INVx1_ASAP7_75t_L g692 ( .A(n_670), .Y(n_692) );
AND2x4_ASAP7_75t_L g785 ( .A(n_670), .B(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g793 ( .A(n_670), .B(n_794), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_676), .Y(n_671) );
AND2x4_ASAP7_75t_SL g672 ( .A(n_673), .B(n_674), .Y(n_672) );
INVx1_ASAP7_75t_SL g736 ( .A(n_673), .Y(n_736) );
INVx2_ASAP7_75t_L g752 ( .A(n_673), .Y(n_752) );
INVx1_ASAP7_75t_L g779 ( .A(n_674), .Y(n_779) );
AND2x2_ASAP7_75t_L g810 ( .A(n_674), .B(n_721), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .C(n_684), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_681), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g722 ( .A(n_682), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_682), .B(n_757), .Y(n_790) );
INVx1_ASAP7_75t_L g710 ( .A(n_683), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_685), .B(n_749), .Y(n_775) );
INVx1_ASAP7_75t_L g730 ( .A(n_686), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_704), .C(n_714), .Y(n_687) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_693), .B(n_700), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
INVx1_ASAP7_75t_L g808 ( .A(n_691), .Y(n_808) );
AND2x4_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI32xp33_ASAP7_75t_L g744 ( .A1(n_695), .A2(n_745), .A3(n_746), .B1(n_747), .B2(n_750), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_695), .B(n_779), .Y(n_778) );
BUFx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g728 ( .A(n_702), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g763 ( .A(n_702), .B(n_723), .Y(n_763) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_707), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g768 ( .A(n_707), .B(n_717), .Y(n_768) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g796 ( .A(n_710), .Y(n_796) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g714 ( .A1(n_712), .A2(n_715), .B1(n_719), .B2(n_722), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_713), .B(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_715), .A2(n_773), .B1(n_810), .B2(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g811 ( .A(n_717), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_719), .A2(n_762), .B1(n_764), .B2(n_768), .Y(n_761) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g803 ( .A(n_723), .Y(n_803) );
NAND4xp25_ASAP7_75t_L g724 ( .A(n_725), .B(n_744), .C(n_753), .D(n_761), .Y(n_724) );
O2A1O1Ixp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_731), .B(n_734), .C(n_735), .Y(n_725) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AND2x4_ASAP7_75t_L g789 ( .A(n_733), .B(n_748), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_733), .B(n_816), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_740), .A2(n_778), .B1(n_780), .B2(n_783), .Y(n_777) );
AND2x4_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OAI21xp5_ASAP7_75t_L g806 ( .A1(n_745), .A2(n_750), .B(n_807), .Y(n_806) );
AND2x4_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI21xp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_758), .Y(n_753) );
INVx2_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NOR2xp33_ASAP7_75t_R g758 ( .A(n_759), .B(n_760), .Y(n_758) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_768), .A2(n_785), .B1(n_822), .B2(n_824), .Y(n_821) );
NOR3x1_ASAP7_75t_L g769 ( .A(n_770), .B(n_791), .C(n_805), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_784), .Y(n_770) );
AOI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B(n_776), .Y(n_771) );
INVx1_ASAP7_75t_L g797 ( .A(n_772), .Y(n_797) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
INVxp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g820 ( .A(n_782), .Y(n_820) );
INVx1_ASAP7_75t_L g794 ( .A(n_786), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_790), .Y(n_787) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_788), .A2(n_792), .B1(n_795), .B2(n_797), .C(n_798), .Y(n_791) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
NAND4xp25_ASAP7_75t_SL g805 ( .A(n_806), .B(n_809), .C(n_813), .D(n_821), .Y(n_805) );
AND2x2_ASAP7_75t_L g819 ( .A(n_812), .B(n_820), .Y(n_819) );
INVxp67_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx4_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
BUFx12f_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_SL g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_836), .Y(n_835) );
BUFx12f_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
BUFx6f_ASAP7_75t_SL g842 ( .A(n_837), .Y(n_842) );
OR2x6_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
endmodule