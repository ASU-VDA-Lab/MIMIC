module fake_netlist_6_2567_n_3029 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_3029);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_3029;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_2647;
wire n_2997;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_883;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_461;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_873;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_405;
wire n_2660;
wire n_538;
wire n_3028;
wire n_2981;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_494;
wire n_539;
wire n_493;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_1815;
wire n_659;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1605;
wire n_1330;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_2693;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_2537;
wire n_2897;
wire n_851;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_417;
wire n_2857;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_1284;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_884;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_2442;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_600;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_2990;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_497;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_401;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3004;
wire n_2830;
wire n_2781;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_664;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_419;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_392;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_621;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_466;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_609;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_579;
wire n_2789;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_411;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_1548;
wire n_799;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_2759;
wire n_1229;
wire n_2945;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_400;
wire n_739;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_506;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1737;
wire n_2430;
wire n_653;
wire n_1464;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_414;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_1537;
wire n_779;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_390;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_924;
wire n_475;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_2600;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_2899;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_120),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_222),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_61),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_315),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_100),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_35),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_215),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_121),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_107),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_299),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_72),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_324),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_68),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_34),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_332),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_61),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_345),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_347),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_128),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_319),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_375),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_137),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_342),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_71),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_360),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_56),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_195),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_77),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_32),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_0),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_120),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_317),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_289),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_201),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_288),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_228),
.Y(n_430)
);

BUFx10_ASAP7_75t_L g431 ( 
.A(n_104),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_349),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_335),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_263),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_339),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_297),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_353),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_48),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_265),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_165),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_309),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_38),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_205),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_179),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_232),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_307),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_305),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_138),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_116),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_102),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_44),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_65),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_241),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_202),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_350),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_139),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_70),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_387),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_362),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_112),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_191),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_50),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_53),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_135),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_101),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_200),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_139),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_55),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_36),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_85),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_100),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_152),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_8),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_209),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_72),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_184),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_198),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_370),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_226),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_84),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_159),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_238),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_128),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_74),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_314),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_91),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_363),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_384),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_300),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_110),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_293),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_115),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_116),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_93),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_327),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_271),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_369),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_348),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_267),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_56),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_249),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_127),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_380),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_230),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_320),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_284),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_174),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_325),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_142),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_340),
.Y(n_512)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_163),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_5),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_216),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_259),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_5),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_211),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_283),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_366),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_6),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_34),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_206),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_88),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_346),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_109),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_93),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_243),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_86),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_213),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_180),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_62),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_164),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_6),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_258),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_180),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_141),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_90),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_9),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_379),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_367),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_329),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_341),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_28),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_376),
.Y(n_545)
);

BUFx2_ASAP7_75t_SL g546 ( 
.A(n_136),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_47),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_229),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_286),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_304),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_356),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_202),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_214),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_132),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_64),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_246),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_364),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_373),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_385),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_279),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_331),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_134),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_208),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_377),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_328),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_344),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_45),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_105),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_89),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_156),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_32),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_176),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_4),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_186),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_42),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_74),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_388),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_378),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_69),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_135),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_127),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_183),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_79),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_386),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_355),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_21),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_12),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_27),
.Y(n_588)
);

BUFx10_ASAP7_75t_L g589 ( 
.A(n_219),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_176),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_131),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_365),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_270),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_193),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_383),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_381),
.Y(n_596)
);

INVxp33_ASAP7_75t_SL g597 ( 
.A(n_336),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_330),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_204),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_89),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_123),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_119),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_117),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_185),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_150),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_240),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_25),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_218),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_382),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_334),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_261),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_9),
.Y(n_612)
);

BUFx5_ASAP7_75t_L g613 ( 
.A(n_110),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_322),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_266),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_70),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_290),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_169),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_358),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_83),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_295),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_53),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_62),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_133),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_52),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_255),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_77),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_95),
.Y(n_628)
);

BUFx10_ASAP7_75t_L g629 ( 
.A(n_10),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_310),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_298),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_185),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_144),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_169),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_69),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_357),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_67),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_11),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_80),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_273),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_59),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_81),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_134),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_11),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_187),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_114),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_179),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_389),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_372),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_158),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_65),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_244),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_275),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_234),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_312),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_143),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_66),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_49),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_190),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_13),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_130),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_4),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_13),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_236),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_326),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_359),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_323),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_76),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_374),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_98),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_115),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_78),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_197),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_31),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_153),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_125),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_368),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_67),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_64),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_343),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_8),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_291),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_23),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_186),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_248),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_167),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_143),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_36),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_212),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_83),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_101),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_20),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_84),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_141),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_285),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_276),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_613),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_613),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_613),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_403),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_613),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_613),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_613),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_513),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_403),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_613),
.Y(n_707)
);

BUFx2_ASAP7_75t_L g708 ( 
.A(n_474),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_613),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_525),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_390),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_390),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_392),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_626),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_392),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_394),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_394),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_569),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_395),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_611),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_396),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_474),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_402),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_602),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_396),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_525),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_602),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_391),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_391),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_605),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_391),
.Y(n_731)
);

INVxp33_ASAP7_75t_L g732 ( 
.A(n_463),
.Y(n_732)
);

INVxp33_ASAP7_75t_SL g733 ( 
.A(n_547),
.Y(n_733)
);

CKINVDCx16_ASAP7_75t_R g734 ( 
.A(n_429),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_391),
.Y(n_735)
);

INVxp67_ASAP7_75t_SL g736 ( 
.A(n_611),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_543),
.Y(n_737)
);

CKINVDCx20_ASAP7_75t_R g738 ( 
.A(n_449),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_405),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_391),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_605),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_651),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_472),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_398),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_398),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_406),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_406),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_407),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_543),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_411),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_411),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_426),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_426),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_432),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_432),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_436),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_436),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_437),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_437),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_651),
.Y(n_760)
);

CKINVDCx16_ASAP7_75t_R g761 ( 
.A(n_431),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_472),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_444),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_444),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_457),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_431),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_457),
.Y(n_767)
);

INVxp33_ASAP7_75t_SL g768 ( 
.A(n_546),
.Y(n_768)
);

INVxp67_ASAP7_75t_SL g769 ( 
.A(n_563),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_476),
.Y(n_770)
);

INVxp33_ASAP7_75t_SL g771 ( 
.A(n_546),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_476),
.Y(n_772)
);

BUFx5_ASAP7_75t_L g773 ( 
.A(n_501),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_465),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_501),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_563),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_598),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_508),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_508),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_510),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_510),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_472),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_399),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_399),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_518),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_518),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_520),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_520),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_523),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_408),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_523),
.Y(n_791)
);

HB1xp67_ASAP7_75t_L g792 ( 
.A(n_418),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_541),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_541),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_549),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_420),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_549),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_598),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_550),
.Y(n_799)
);

CKINVDCx16_ASAP7_75t_R g800 ( 
.A(n_431),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_471),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_550),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_553),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_472),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_483),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_421),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_553),
.Y(n_807)
);

INVxp33_ASAP7_75t_SL g808 ( 
.A(n_422),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_559),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_559),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_565),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_565),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_626),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_596),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_578),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_578),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_472),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_595),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_424),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_626),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_522),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_486),
.Y(n_822)
);

INVxp33_ASAP7_75t_SL g823 ( 
.A(n_425),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_509),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_595),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_527),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_606),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_522),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_428),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_537),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_522),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_601),
.Y(n_832)
);

HB1xp67_ASAP7_75t_L g833 ( 
.A(n_441),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_596),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_632),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_400),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_522),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_522),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_769),
.B(n_427),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_734),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_728),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

OAI22x1_ASAP7_75t_SL g843 ( 
.A1(n_738),
.A2(n_650),
.B1(n_676),
.B2(n_635),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_738),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_762),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_777),
.B(n_427),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_782),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_705),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_733),
.A2(n_597),
.B1(n_456),
.B2(n_481),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_782),
.Y(n_850)
);

INVx6_ASAP7_75t_L g851 ( 
.A(n_714),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_804),
.Y(n_852)
);

BUFx8_ASAP7_75t_L g853 ( 
.A(n_708),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_728),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_733),
.A2(n_718),
.B1(n_736),
.B2(n_720),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_804),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_714),
.Y(n_857)
);

OA21x2_ASAP7_75t_L g858 ( 
.A1(n_702),
.A2(n_704),
.B(n_703),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_714),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_817),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_SL g861 ( 
.A1(n_774),
.A2(n_683),
.B1(n_416),
.B2(n_455),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_814),
.B(n_596),
.Y(n_862)
);

AND2x6_ASAP7_75t_L g863 ( 
.A(n_714),
.B(n_626),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_817),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_729),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_821),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_729),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_798),
.B(n_503),
.Y(n_868)
);

BUFx8_ASAP7_75t_L g869 ( 
.A(n_708),
.Y(n_869)
);

BUFx8_ASAP7_75t_SL g870 ( 
.A(n_774),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_SL g871 ( 
.A1(n_801),
.A2(n_423),
.B1(n_625),
.B2(n_581),
.Y(n_871)
);

OAI22x1_ASAP7_75t_R g872 ( 
.A1(n_801),
.A2(n_452),
.B1(n_453),
.B2(n_450),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_714),
.Y(n_873)
);

AND2x6_ASAP7_75t_L g874 ( 
.A(n_813),
.B(n_626),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_834),
.B(n_503),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_706),
.A2(n_730),
.B1(n_742),
.B2(n_722),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_821),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_731),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_731),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_813),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_813),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_805),
.A2(n_548),
.B1(n_558),
.B2(n_414),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_813),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_813),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_735),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_761),
.A2(n_592),
.B1(n_682),
.B2(n_560),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_760),
.A2(n_594),
.B1(n_459),
.B2(n_467),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_820),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_735),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_820),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_740),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_740),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_820),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_710),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_743),
.Y(n_895)
);

OA21x2_ASAP7_75t_L g896 ( 
.A1(n_707),
.A2(n_653),
.B(n_606),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_743),
.Y(n_897)
);

INVx5_ASAP7_75t_L g898 ( 
.A(n_820),
.Y(n_898)
);

INVx5_ASAP7_75t_L g899 ( 
.A(n_710),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_732),
.A2(n_462),
.B1(n_473),
.B2(n_470),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_792),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_828),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_726),
.Y(n_903)
);

AND2x6_ASAP7_75t_L g904 ( 
.A(n_697),
.B(n_440),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_828),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_831),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_831),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_837),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_705),
.Y(n_909)
);

NOR2x1_ASAP7_75t_L g910 ( 
.A(n_837),
.B(n_653),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_726),
.B(n_464),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_737),
.B(n_440),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_737),
.B(n_491),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_719),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_724),
.A2(n_482),
.B1(n_485),
.B2(n_477),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_749),
.B(n_491),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_838),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_749),
.B(n_519),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_838),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_776),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_711),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_709),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_800),
.A2(n_808),
.B1(n_823),
.B2(n_771),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_776),
.Y(n_924)
);

BUFx8_ASAP7_75t_SL g925 ( 
.A(n_805),
.Y(n_925)
);

INVx5_ASAP7_75t_L g926 ( 
.A(n_766),
.Y(n_926)
);

OA21x2_ASAP7_75t_L g927 ( 
.A1(n_697),
.A2(n_689),
.B(n_599),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_712),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_808),
.A2(n_494),
.B1(n_496),
.B2(n_495),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_698),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_713),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_698),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_715),
.B(n_519),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_716),
.B(n_599),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_717),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_724),
.A2(n_504),
.B1(n_517),
.B2(n_511),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_699),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_773),
.B(n_608),
.Y(n_938)
);

OAI22x1_ASAP7_75t_SL g939 ( 
.A1(n_822),
.A2(n_524),
.B1(n_526),
.B2(n_521),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_721),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_725),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_766),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_699),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_823),
.B(n_768),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_744),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_719),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_745),
.Y(n_947)
);

OA21x2_ASAP7_75t_L g948 ( 
.A1(n_700),
.A2(n_689),
.B(n_640),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_700),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_783),
.B(n_464),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_773),
.B(n_608),
.Y(n_951)
);

CKINVDCx11_ASAP7_75t_R g952 ( 
.A(n_822),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_784),
.B(n_573),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_773),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_768),
.B(n_415),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_746),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_824),
.Y(n_957)
);

BUFx3_ASAP7_75t_L g958 ( 
.A(n_747),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_750),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_773),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_751),
.B(n_640),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_752),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_870),
.Y(n_963)
);

CKINVDCx20_ASAP7_75t_R g964 ( 
.A(n_870),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_842),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_921),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_962),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_842),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_925),
.Y(n_969)
);

INVxp33_ASAP7_75t_L g970 ( 
.A(n_872),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_857),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_928),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_925),
.Y(n_973)
);

OR2x2_ASAP7_75t_L g974 ( 
.A(n_876),
.B(n_833),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_952),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_894),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_952),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_840),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_R g979 ( 
.A(n_914),
.B(n_723),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_848),
.B(n_771),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_857),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_840),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_848),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_914),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_909),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_909),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_853),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_853),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_911),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_853),
.Y(n_990)
);

CKINVDCx20_ASAP7_75t_R g991 ( 
.A(n_844),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_869),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_859),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_955),
.B(n_723),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_931),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_845),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_844),
.B(n_739),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_894),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_935),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_859),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_940),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_926),
.B(n_739),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_941),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_957),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_901),
.B(n_748),
.Y(n_1005)
);

BUFx10_ASAP7_75t_L g1006 ( 
.A(n_944),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_945),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_957),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_946),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_946),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_903),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_903),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_869),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_R g1014 ( 
.A(n_926),
.B(n_748),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_845),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_869),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_886),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_947),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_923),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_847),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_882),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_849),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_847),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_855),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_959),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_920),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_920),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_929),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_859),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_958),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_859),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_843),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_861),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_939),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_900),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_958),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_915),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_930),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_930),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_936),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_R g1041 ( 
.A(n_926),
.B(n_790),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_887),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_871),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_859),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_911),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_862),
.B(n_753),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_839),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_926),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_862),
.B(n_754),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_926),
.B(n_773),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_937),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_937),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_899),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_932),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_943),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_850),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_943),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_949),
.Y(n_1058)
);

CKINVDCx16_ASAP7_75t_R g1059 ( 
.A(n_950),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_846),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_850),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_868),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_950),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_953),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_953),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_875),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_949),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_899),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_852),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_932),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_918),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_918),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_932),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_932),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_918),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_862),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_852),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_942),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_942),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_956),
.Y(n_1080)
);

CKINVDCx20_ASAP7_75t_R g1081 ( 
.A(n_942),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_942),
.B(n_755),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_857),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_942),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_912),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_856),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_913),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_899),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_899),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_916),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_956),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_890),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_899),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_924),
.B(n_773),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_924),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_924),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_924),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_956),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_933),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_922),
.B(n_773),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_933),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_933),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_934),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_934),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_934),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_956),
.Y(n_1106)
);

AND2x6_ASAP7_75t_L g1107 ( 
.A(n_910),
.B(n_685),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_856),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_961),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_858),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_961),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_860),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_961),
.Y(n_1113)
);

CKINVDCx20_ASAP7_75t_R g1114 ( 
.A(n_896),
.Y(n_1114)
);

CKINVDCx16_ASAP7_75t_R g1115 ( 
.A(n_904),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_841),
.B(n_790),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_956),
.B(n_796),
.Y(n_1117)
);

XNOR2xp5_ASAP7_75t_L g1118 ( 
.A(n_896),
.B(n_824),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_904),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_896),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_904),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_904),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_854),
.Y(n_1123)
);

XNOR2xp5_ASAP7_75t_L g1124 ( 
.A(n_927),
.B(n_826),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_R g1125 ( 
.A(n_865),
.B(n_796),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_922),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_922),
.B(n_773),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_860),
.Y(n_1128)
);

CKINVDCx20_ASAP7_75t_R g1129 ( 
.A(n_938),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_922),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_904),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_904),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_1110),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1110),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_971),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1011),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1123),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1063),
.B(n_741),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_966),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_967),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_SL g1141 ( 
.A(n_1006),
.Y(n_1141)
);

AND3x4_ASAP7_75t_L g1142 ( 
.A(n_1011),
.B(n_830),
.C(n_826),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_971),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_1045),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_965),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1047),
.B(n_1062),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1090),
.B(n_806),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_994),
.B(n_806),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1085),
.B(n_858),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1087),
.B(n_819),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_965),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_968),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_968),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_989),
.B(n_685),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_972),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_996),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_996),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_995),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_999),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_989),
.B(n_756),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1030),
.B(n_757),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1129),
.A2(n_829),
.B1(n_819),
.B2(n_499),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1001),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_1046),
.B(n_400),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1003),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1015),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_991),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1007),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1059),
.B(n_829),
.Y(n_1169)
);

AND2x2_ASAP7_75t_SL g1170 ( 
.A(n_1115),
.B(n_927),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1018),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1076),
.B(n_1065),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1025),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1015),
.Y(n_1174)
);

AND2x6_ASAP7_75t_L g1175 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_984),
.B(n_830),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1049),
.B(n_858),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1020),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1020),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1064),
.B(n_741),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1036),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1026),
.B(n_701),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1027),
.B(n_727),
.Y(n_1183)
);

BUFx8_ASAP7_75t_SL g1184 ( 
.A(n_969),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1005),
.B(n_836),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_971),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1023),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_976),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_998),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1114),
.A2(n_948),
.B1(n_927),
.B2(n_413),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_1089),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1071),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1082),
.B(n_922),
.Y(n_1193)
);

AND2x2_ASAP7_75t_SL g1194 ( 
.A(n_974),
.B(n_948),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_1023),
.Y(n_1195)
);

INVx5_ASAP7_75t_L g1196 ( 
.A(n_1107),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1120),
.B(n_954),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1124),
.B(n_532),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1056),
.Y(n_1199)
);

AND2x2_ASAP7_75t_SL g1200 ( 
.A(n_980),
.B(n_948),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1056),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1117),
.B(n_532),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1061),
.Y(n_1203)
);

AND2x6_ASAP7_75t_L g1204 ( 
.A(n_1126),
.B(n_410),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_971),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_1072),
.B(n_758),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1061),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_1075),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1118),
.B(n_534),
.C(n_529),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1069),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1102),
.B(n_1103),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1069),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1082),
.B(n_954),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1054),
.B(n_1070),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1038),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1102),
.B(n_954),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1004),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_971),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1066),
.B(n_497),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1012),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1073),
.B(n_960),
.Y(n_1221)
);

AND2x6_ASAP7_75t_L g1222 ( 
.A(n_1130),
.B(n_410),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1039),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1103),
.B(n_759),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1074),
.B(n_960),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1035),
.B(n_507),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_981),
.Y(n_1227)
);

BUFx2_ASAP7_75t_L g1228 ( 
.A(n_1008),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1077),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1051),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1052),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1081),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1104),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1055),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1057),
.B(n_960),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1035),
.B(n_512),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1077),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1058),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1067),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1006),
.B(n_832),
.Y(n_1240)
);

INVx5_ASAP7_75t_L g1241 ( 
.A(n_1107),
.Y(n_1241)
);

BUFx2_ASAP7_75t_L g1242 ( 
.A(n_997),
.Y(n_1242)
);

AO22x2_ASAP7_75t_L g1243 ( 
.A1(n_1037),
.A2(n_679),
.B1(n_627),
.B2(n_439),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_969),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1084),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1060),
.B(n_649),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1104),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1086),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1105),
.B(n_654),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1086),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1105),
.B(n_763),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1108),
.Y(n_1252)
);

NOR3xp33_ASAP7_75t_L g1253 ( 
.A(n_1022),
.B(n_679),
.C(n_627),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1006),
.B(n_1109),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1009),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1108),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1112),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1112),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1128),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1109),
.B(n_536),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1128),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_993),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1111),
.B(n_1113),
.Y(n_1263)
);

NAND2xp33_ASAP7_75t_L g1264 ( 
.A(n_1119),
.B(n_863),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1099),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1111),
.B(n_867),
.Y(n_1266)
);

AND2x2_ASAP7_75t_SL g1267 ( 
.A(n_1080),
.B(n_690),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1101),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1113),
.B(n_764),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1091),
.Y(n_1270)
);

INVxp33_ASAP7_75t_SL g1271 ( 
.A(n_979),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1098),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_981),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1033),
.A2(n_835),
.B1(n_832),
.B2(n_544),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1119),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1107),
.A2(n_514),
.B1(n_607),
.B2(n_413),
.Y(n_1276)
);

INVx3_ASAP7_75t_L g1277 ( 
.A(n_993),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1106),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1010),
.B(n_835),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_985),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1042),
.B(n_538),
.Y(n_1281)
);

AO22x2_ASAP7_75t_L g1282 ( 
.A1(n_1037),
.A2(n_439),
.B1(n_445),
.B2(n_443),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_993),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1000),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_981),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1000),
.Y(n_1286)
);

AND2x6_ASAP7_75t_L g1287 ( 
.A(n_1100),
.B(n_443),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1000),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1029),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_981),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_985),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_986),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1029),
.Y(n_1293)
);

BUFx10_ASAP7_75t_L g1294 ( 
.A(n_978),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1029),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1116),
.B(n_431),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1031),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1031),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1031),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1121),
.B(n_765),
.Y(n_1300)
);

OR2x6_ASAP7_75t_L g1301 ( 
.A(n_1002),
.B(n_514),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1044),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1121),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1044),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1044),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1092),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_981),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1125),
.B(n_629),
.Y(n_1308)
);

AND2x2_ASAP7_75t_SL g1309 ( 
.A(n_1127),
.B(n_690),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1092),
.B(n_878),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1028),
.B(n_552),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1092),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1122),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1122),
.B(n_951),
.Y(n_1314)
);

AND2x6_ASAP7_75t_L g1315 ( 
.A(n_1050),
.B(n_445),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1083),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1107),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_986),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1107),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1107),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1048),
.B(n_889),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1083),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1048),
.B(n_891),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1083),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_1132),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1131),
.B(n_393),
.Y(n_1326)
);

INVx5_ASAP7_75t_L g1327 ( 
.A(n_1134),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1248),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1190),
.A2(n_1040),
.B1(n_1019),
.B2(n_1017),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1252),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1148),
.B(n_1014),
.Y(n_1331)
);

INVx5_ASAP7_75t_L g1332 ( 
.A(n_1134),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1148),
.B(n_1185),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1194),
.B(n_1041),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1194),
.B(n_1078),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1226),
.B(n_984),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1145),
.Y(n_1337)
);

OAI221xp5_ASAP7_75t_L g1338 ( 
.A1(n_1226),
.A2(n_1021),
.B1(n_478),
.B2(n_770),
.C(n_772),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1236),
.B(n_983),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1134),
.B(n_1131),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1136),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1145),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_SL g1343 ( 
.A(n_1271),
.B(n_978),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1190),
.B(n_1079),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1256),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1236),
.B(n_1132),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1134),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1141),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1151),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1133),
.A2(n_983),
.B1(n_1024),
.B2(n_1043),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1160),
.B(n_1088),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1146),
.B(n_982),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1146),
.B(n_982),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1175),
.A2(n_589),
.B1(n_619),
.B2(n_907),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1257),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1160),
.B(n_1093),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1258),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1160),
.B(n_1095),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1175),
.B(n_1096),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1147),
.B(n_1281),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1175),
.B(n_1097),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_SL g1362 ( 
.A(n_1133),
.B(n_987),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1175),
.B(n_906),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1151),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1133),
.B(n_987),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1259),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1175),
.A2(n_589),
.B1(n_619),
.B2(n_690),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1152),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1182),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1154),
.B(n_906),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1154),
.B(n_906),
.Y(n_1371)
);

INVx3_ASAP7_75t_L g1372 ( 
.A(n_1262),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1154),
.B(n_906),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1149),
.B(n_919),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1147),
.B(n_1300),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1300),
.B(n_919),
.Y(n_1376)
);

INVxp33_ASAP7_75t_L g1377 ( 
.A(n_1183),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_SL g1378 ( 
.A(n_1200),
.B(n_988),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1262),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1186),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1200),
.B(n_988),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1170),
.B(n_990),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1300),
.B(n_919),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1261),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1180),
.B(n_767),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1152),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1136),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1170),
.B(n_990),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1262),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1153),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1249),
.B(n_919),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1153),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1281),
.B(n_970),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1156),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1156),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1177),
.A2(n_1213),
.B(n_1309),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1249),
.B(n_397),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1197),
.B(n_992),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1157),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1139),
.B(n_401),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1138),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1164),
.A2(n_1197),
.B1(n_1287),
.B2(n_1309),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1140),
.B(n_404),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1260),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_SL g1405 ( 
.A(n_1271),
.B(n_992),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1157),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1150),
.B(n_963),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1325),
.B(n_1013),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_SL g1409 ( 
.A(n_1325),
.B(n_1016),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1166),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1174),
.Y(n_1411)
);

NOR2xp67_ASAP7_75t_L g1412 ( 
.A(n_1233),
.B(n_975),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1174),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1178),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1178),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1150),
.B(n_975),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1277),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1179),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1155),
.B(n_409),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1325),
.B(n_1094),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1158),
.B(n_412),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1314),
.A2(n_1193),
.B(n_1317),
.Y(n_1422)
);

AND2x6_ASAP7_75t_SL g1423 ( 
.A(n_1311),
.B(n_451),
.Y(n_1423)
);

INVx8_ASAP7_75t_L g1424 ( 
.A(n_1164),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1159),
.B(n_417),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1277),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1179),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1187),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1163),
.B(n_419),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1187),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1233),
.B(n_690),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1313),
.A2(n_433),
.B1(n_434),
.B2(n_430),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1165),
.B(n_435),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1199),
.Y(n_1434)
);

INVx3_ASAP7_75t_L g1435 ( 
.A(n_1277),
.Y(n_1435)
);

NOR3xp33_ASAP7_75t_L g1436 ( 
.A(n_1311),
.B(n_973),
.C(n_977),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1219),
.B(n_977),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1221),
.A2(n_898),
.B(n_1053),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1168),
.B(n_438),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1202),
.A2(n_1301),
.B1(n_1198),
.B2(n_1266),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1171),
.B(n_442),
.Y(n_1441)
);

INVx3_ASAP7_75t_L g1442 ( 
.A(n_1283),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_R g1443 ( 
.A(n_1244),
.B(n_973),
.Y(n_1443)
);

AND2x6_ASAP7_75t_SL g1444 ( 
.A(n_1279),
.B(n_451),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1186),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1201),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1173),
.B(n_446),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1219),
.B(n_964),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1215),
.B(n_447),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1203),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1246),
.B(n_1034),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1223),
.B(n_448),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1230),
.B(n_1231),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1203),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1325),
.B(n_1053),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1234),
.B(n_454),
.Y(n_1456)
);

AND2x6_ASAP7_75t_SL g1457 ( 
.A(n_1246),
.B(n_458),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1238),
.B(n_460),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1162),
.B(n_1034),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1239),
.B(n_461),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1313),
.B(n_480),
.Y(n_1461)
);

INVx2_ASAP7_75t_SL g1462 ( 
.A(n_1206),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1224),
.B(n_775),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1283),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1164),
.B(n_484),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1210),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1164),
.B(n_1224),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1164),
.B(n_487),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1210),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1212),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1206),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1196),
.B(n_1068),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1212),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1237),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1327),
.A2(n_1307),
.B(n_1314),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1360),
.B(n_1209),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1375),
.B(n_1254),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1368),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1333),
.B(n_1346),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1336),
.B(n_1291),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1338),
.A2(n_1211),
.B(n_1172),
.C(n_1253),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1404),
.B(n_1331),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1385),
.B(n_1224),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1385),
.B(n_1169),
.Y(n_1484)
);

BUFx2_ASAP7_75t_SL g1485 ( 
.A(n_1412),
.Y(n_1485)
);

O2A1O1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1339),
.A2(n_1211),
.B(n_1172),
.C(n_1260),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1337),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1327),
.B(n_1263),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1397),
.B(n_1251),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1251),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_1377),
.B(n_1255),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1380),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1377),
.B(n_1144),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1327),
.A2(n_1307),
.B(n_1216),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1401),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1380),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1368),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1420),
.A2(n_1216),
.B(n_1270),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1396),
.A2(n_1320),
.B(n_1319),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1344),
.A2(n_1275),
.B1(n_1303),
.B2(n_1263),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_SL g1501 ( 
.A1(n_1440),
.A2(n_1278),
.B(n_1272),
.C(n_1286),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1348),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1463),
.B(n_1251),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1327),
.A2(n_1307),
.B(n_1205),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1369),
.B(n_1296),
.Y(n_1505)
);

O2A1O1Ixp33_ASAP7_75t_L g1506 ( 
.A1(n_1329),
.A2(n_1137),
.B(n_1268),
.C(n_1265),
.Y(n_1506)
);

NOR2xp67_ASAP7_75t_L g1507 ( 
.A(n_1352),
.B(n_1247),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1327),
.A2(n_1205),
.B(n_1186),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1422),
.A2(n_1235),
.B(n_1225),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_SL g1510 ( 
.A(n_1332),
.B(n_1402),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1353),
.B(n_1308),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1391),
.B(n_1269),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1337),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1367),
.A2(n_1276),
.B1(n_1282),
.B2(n_1287),
.Y(n_1514)
);

A2O1A1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1393),
.A2(n_1276),
.B(n_1269),
.C(n_1275),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1407),
.B(n_1416),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1469),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1437),
.B(n_1280),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1469),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_R g1520 ( 
.A(n_1343),
.B(n_1244),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1332),
.A2(n_1205),
.B(n_1186),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1341),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1453),
.B(n_1269),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1462),
.B(n_1263),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1332),
.A2(n_1218),
.B(n_1205),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1332),
.A2(n_1227),
.B(n_1218),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1342),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1392),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1332),
.Y(n_1529)
);

INVx4_ASAP7_75t_L g1530 ( 
.A(n_1380),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1342),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1334),
.A2(n_1335),
.B1(n_1467),
.B2(n_1303),
.Y(n_1532)
);

AO21x1_ASAP7_75t_L g1533 ( 
.A1(n_1378),
.A2(n_1310),
.B(n_1214),
.Y(n_1533)
);

OAI321xp33_ASAP7_75t_L g1534 ( 
.A1(n_1451),
.A2(n_1202),
.A3(n_1138),
.B1(n_1301),
.B2(n_469),
.C(n_466),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1341),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1374),
.A2(n_1250),
.B(n_1326),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1462),
.B(n_1206),
.Y(n_1537)
);

AOI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1420),
.A2(n_1227),
.B(n_1218),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1340),
.A2(n_1227),
.B(n_1218),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1349),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1471),
.B(n_1161),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1340),
.A2(n_1321),
.B1(n_1323),
.B2(n_1192),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1376),
.A2(n_1290),
.B(n_1227),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1471),
.B(n_1161),
.Y(n_1544)
);

OAI21xp5_ASAP7_75t_L g1545 ( 
.A1(n_1370),
.A2(n_1250),
.B(n_1326),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1350),
.B(n_1292),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_L g1547 ( 
.A1(n_1383),
.A2(n_1316),
.B(n_1290),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1398),
.A2(n_1181),
.B(n_1161),
.C(n_1220),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1363),
.A2(n_1316),
.B(n_1290),
.Y(n_1549)
);

NOR2xp67_ASAP7_75t_L g1550 ( 
.A(n_1408),
.B(n_1188),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1371),
.A2(n_1316),
.B(n_1290),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1410),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1347),
.Y(n_1553)
);

AO21x1_ASAP7_75t_L g1554 ( 
.A1(n_1378),
.A2(n_1295),
.B(n_1289),
.Y(n_1554)
);

NOR2xp33_ASAP7_75t_L g1555 ( 
.A(n_1382),
.B(n_1318),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1373),
.A2(n_1316),
.B(n_1143),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1351),
.B(n_1301),
.Y(n_1557)
);

CKINVDCx10_ASAP7_75t_R g1558 ( 
.A(n_1443),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1411),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1414),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1455),
.A2(n_1273),
.B(n_1135),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1455),
.A2(n_1285),
.B(n_1264),
.Y(n_1562)
);

A2O1A1Ixp33_ASAP7_75t_SL g1563 ( 
.A1(n_1476),
.A2(n_1354),
.B(n_1347),
.C(n_1465),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1479),
.B(n_1398),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1487),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1516),
.B(n_1167),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1509),
.A2(n_1424),
.B(n_1264),
.Y(n_1567)
);

O2A1O1Ixp5_ASAP7_75t_L g1568 ( 
.A1(n_1516),
.A2(n_1476),
.B(n_1510),
.C(n_1554),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1528),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_R g1570 ( 
.A(n_1502),
.B(n_1405),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_L g1571 ( 
.A1(n_1480),
.A2(n_1176),
.B(n_1459),
.Y(n_1571)
);

INVx4_ASAP7_75t_L g1572 ( 
.A(n_1492),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1552),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1511),
.B(n_1356),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1486),
.B(n_1381),
.Y(n_1575)
);

INVx11_ASAP7_75t_L g1576 ( 
.A(n_1558),
.Y(n_1576)
);

A2O1A1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1515),
.A2(n_1424),
.B(n_1328),
.C(n_1345),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1492),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1482),
.B(n_1358),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1523),
.B(n_1483),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1484),
.B(n_1382),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1559),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1535),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1487),
.Y(n_1584)
);

OAI21xp33_ASAP7_75t_L g1585 ( 
.A1(n_1480),
.A2(n_1176),
.B(n_1240),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1489),
.A2(n_1424),
.B(n_1361),
.Y(n_1586)
);

BUFx8_ASAP7_75t_L g1587 ( 
.A(n_1505),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1518),
.B(n_1217),
.Y(n_1588)
);

NOR2xp67_ASAP7_75t_L g1589 ( 
.A(n_1491),
.B(n_1220),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1492),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1513),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1560),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1490),
.B(n_1388),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1478),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_SL g1595 ( 
.A(n_1481),
.B(n_1142),
.C(n_1242),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1555),
.A2(n_1388),
.B1(n_1381),
.B2(n_1142),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1510),
.A2(n_1424),
.B(n_1359),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1491),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1492),
.Y(n_1599)
);

O2A1O1Ixp5_ASAP7_75t_L g1600 ( 
.A1(n_1533),
.A2(n_1365),
.B(n_1362),
.C(n_1408),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1503),
.B(n_1387),
.Y(n_1601)
);

AOI33xp33_ASAP7_75t_L g1602 ( 
.A1(n_1506),
.A2(n_469),
.A3(n_466),
.B1(n_475),
.B2(n_468),
.B3(n_458),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1512),
.B(n_1387),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1513),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1495),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1497),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1536),
.A2(n_1241),
.B(n_1196),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1524),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1529),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1517),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1531),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1496),
.Y(n_1612)
);

AOI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1498),
.A2(n_1428),
.B(n_1418),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1477),
.B(n_1400),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1546),
.A2(n_1274),
.B1(n_1448),
.B2(n_1141),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1613),
.A2(n_1538),
.B(n_1499),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1567),
.A2(n_1515),
.B(n_1494),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1568),
.A2(n_1542),
.B(n_1477),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1594),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_SL g1621 ( 
.A(n_1575),
.B(n_1485),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1576),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1571),
.A2(n_1514),
.B(n_1534),
.C(n_1548),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1613),
.A2(n_1539),
.B(n_1562),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1586),
.A2(n_1545),
.B(n_1549),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1606),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1600),
.A2(n_1575),
.B(n_1614),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1583),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1610),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1608),
.B(n_1488),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1607),
.A2(n_1475),
.B(n_1532),
.Y(n_1631)
);

AOI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1597),
.A2(n_1500),
.B(n_1543),
.Y(n_1632)
);

INVx4_ASAP7_75t_L g1633 ( 
.A(n_1590),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1565),
.A2(n_1547),
.B(n_1551),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1564),
.A2(n_1548),
.B(n_1507),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1565),
.A2(n_1556),
.B(n_1561),
.Y(n_1636)
);

AO32x2_ASAP7_75t_L g1637 ( 
.A1(n_1602),
.A2(n_1282),
.A3(n_1432),
.B1(n_1243),
.B2(n_1530),
.Y(n_1637)
);

AO21x2_ASAP7_75t_L g1638 ( 
.A1(n_1577),
.A2(n_1501),
.B(n_1508),
.Y(n_1638)
);

O2A1O1Ixp5_ASAP7_75t_L g1639 ( 
.A1(n_1577),
.A2(n_1563),
.B(n_1518),
.C(n_1362),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1584),
.A2(n_1504),
.B(n_1521),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1580),
.B(n_1555),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1563),
.A2(n_1501),
.B(n_1529),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1584),
.A2(n_1526),
.B(n_1525),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1591),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1598),
.B(n_1493),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1602),
.A2(n_1514),
.B(n_1557),
.C(n_1493),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1593),
.A2(n_1488),
.B(n_1468),
.Y(n_1647)
);

AOI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1603),
.A2(n_1574),
.B(n_1595),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1605),
.Y(n_1649)
);

OAI21xp5_ASAP7_75t_L g1650 ( 
.A1(n_1589),
.A2(n_1461),
.B(n_1419),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1588),
.B(n_1537),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1572),
.Y(n_1652)
);

BUFx8_ASAP7_75t_L g1653 ( 
.A(n_1608),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1576),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1569),
.Y(n_1655)
);

CKINVDCx14_ASAP7_75t_R g1656 ( 
.A(n_1570),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_L g1657 ( 
.A1(n_1591),
.A2(n_1438),
.B(n_1531),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1585),
.A2(n_1436),
.B1(n_1228),
.B2(n_1141),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_SL g1659 ( 
.A(n_1590),
.B(n_1496),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1601),
.B(n_1208),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_SL g1661 ( 
.A1(n_1581),
.A2(n_1365),
.B(n_1409),
.C(n_1519),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1604),
.A2(n_1379),
.B(n_1372),
.Y(n_1662)
);

NAND2x1_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1530),
.Y(n_1663)
);

AOI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1596),
.A2(n_1550),
.B1(n_1208),
.B2(n_1032),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1590),
.Y(n_1665)
);

OAI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1624),
.A2(n_1625),
.B(n_1632),
.Y(n_1666)
);

OAI211xp5_ASAP7_75t_L g1667 ( 
.A1(n_1664),
.A2(n_1615),
.B(n_1520),
.C(n_1032),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1620),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1622),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1622),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1626),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1619),
.B(n_1583),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1618),
.A2(n_1658),
.B1(n_1651),
.B2(n_1660),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_SL g1674 ( 
.A1(n_1621),
.A2(n_1582),
.B(n_1573),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1653),
.A2(n_1282),
.B1(n_1243),
.B2(n_1520),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1624),
.A2(n_1631),
.B(n_1617),
.Y(n_1676)
);

CKINVDCx11_ASAP7_75t_R g1677 ( 
.A(n_1649),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1627),
.A2(n_779),
.B(n_778),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1629),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1655),
.Y(n_1680)
);

AO21x2_ASAP7_75t_L g1681 ( 
.A1(n_1642),
.A2(n_1409),
.B(n_1592),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1644),
.Y(n_1682)
);

NAND2x1p5_ASAP7_75t_L g1683 ( 
.A(n_1641),
.B(n_1630),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1645),
.A2(n_1202),
.B1(n_1423),
.B2(n_1245),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1644),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1630),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1662),
.Y(n_1687)
);

OA21x2_ASAP7_75t_L g1688 ( 
.A1(n_1616),
.A2(n_781),
.B(n_780),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1630),
.B(n_1572),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1641),
.B(n_1457),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1648),
.A2(n_1243),
.B1(n_661),
.B2(n_675),
.Y(n_1691)
);

AOI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1647),
.A2(n_1452),
.B(n_1449),
.Y(n_1692)
);

BUFx2_ASAP7_75t_L g1693 ( 
.A(n_1653),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1639),
.A2(n_1458),
.B(n_1456),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1635),
.A2(n_1611),
.B(n_1472),
.Y(n_1695)
);

INVx4_ASAP7_75t_L g1696 ( 
.A(n_1665),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_L g1697 ( 
.A(n_1628),
.B(n_1587),
.Y(n_1697)
);

INVxp33_ASAP7_75t_L g1698 ( 
.A(n_1665),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1662),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1633),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1633),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1616),
.A2(n_786),
.B(n_785),
.Y(n_1702)
);

INVx6_ASAP7_75t_L g1703 ( 
.A(n_1653),
.Y(n_1703)
);

OAI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1636),
.A2(n_1604),
.B(n_1611),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1634),
.A2(n_1657),
.B(n_1640),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1661),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1665),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1657),
.A2(n_1609),
.B(n_1364),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1638),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1650),
.A2(n_1202),
.B1(n_1245),
.B2(n_1232),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1623),
.B(n_1646),
.C(n_1587),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1638),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1665),
.Y(n_1714)
);

AO31x2_ASAP7_75t_L g1715 ( 
.A1(n_1623),
.A2(n_1612),
.A3(n_1578),
.B(n_1572),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1646),
.B(n_1587),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1643),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1663),
.B(n_1633),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_L g1719 ( 
.A1(n_1656),
.A2(n_575),
.B1(n_576),
.B2(n_570),
.C(n_554),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1654),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1652),
.B(n_1138),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1652),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1659),
.A2(n_1609),
.B(n_1364),
.Y(n_1723)
);

BUFx2_ASAP7_75t_SL g1724 ( 
.A(n_1656),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1637),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1637),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1637),
.A2(n_788),
.B(n_787),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1637),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1654),
.A2(n_1191),
.B1(n_1294),
.B2(n_1232),
.Y(n_1729)
);

BUFx3_ASAP7_75t_L g1730 ( 
.A(n_1628),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1620),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1620),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_L g1733 ( 
.A1(n_1648),
.A2(n_1460),
.B(n_1421),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1619),
.A2(n_1348),
.B1(n_1294),
.B2(n_1191),
.Y(n_1734)
);

AOI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1617),
.A2(n_1241),
.B(n_1196),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1624),
.A2(n_1386),
.B(n_1349),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1618),
.B(n_1612),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1664),
.A2(n_1522),
.B1(n_1544),
.B2(n_1541),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1641),
.A2(n_661),
.B1(n_675),
.B2(n_573),
.Y(n_1739)
);

OAI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1624),
.A2(n_1390),
.B(n_1386),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1617),
.A2(n_1241),
.B(n_1196),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1623),
.A2(n_1267),
.B(n_638),
.C(n_681),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1664),
.A2(n_1301),
.B1(n_1431),
.B2(n_1425),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1651),
.B(n_1431),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1624),
.A2(n_1394),
.B(n_1390),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1665),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1664),
.A2(n_1294),
.B1(n_1429),
.B2(n_1403),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1620),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1617),
.A2(n_1241),
.B(n_1267),
.Y(n_1749)
);

INVx4_ASAP7_75t_L g1750 ( 
.A(n_1665),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1644),
.Y(n_1751)
);

INVxp67_ASAP7_75t_L g1752 ( 
.A(n_1681),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1733),
.A2(n_1347),
.B(n_1472),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1696),
.Y(n_1754)
);

BUFx2_ASAP7_75t_R g1755 ( 
.A(n_1724),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1696),
.Y(n_1756)
);

AO31x2_ASAP7_75t_L g1757 ( 
.A1(n_1710),
.A2(n_1578),
.A3(n_791),
.B(n_793),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1668),
.B(n_789),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1673),
.B(n_1590),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1671),
.Y(n_1760)
);

INVx3_ASAP7_75t_L g1761 ( 
.A(n_1696),
.Y(n_1761)
);

AO21x2_ASAP7_75t_L g1762 ( 
.A1(n_1666),
.A2(n_1439),
.B(n_1433),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1679),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1730),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1680),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1731),
.B(n_794),
.Y(n_1766)
);

BUFx6f_ASAP7_75t_L g1767 ( 
.A(n_1677),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1732),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1748),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1666),
.A2(n_1553),
.B(n_1355),
.Y(n_1770)
);

AO31x2_ASAP7_75t_L g1771 ( 
.A1(n_1710),
.A2(n_1578),
.A3(n_797),
.B(n_799),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1726),
.B(n_795),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1749),
.A2(n_1445),
.B(n_1380),
.Y(n_1773)
);

A2O1A1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1712),
.A2(n_638),
.B(n_681),
.C(n_607),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1751),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1682),
.Y(n_1776)
);

OAI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1706),
.A2(n_1553),
.B(n_1357),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1690),
.A2(n_629),
.B1(n_475),
.B2(n_479),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1730),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1683),
.B(n_468),
.Y(n_1780)
);

BUFx12f_ASAP7_75t_L g1781 ( 
.A(n_1669),
.Y(n_1781)
);

OA21x2_ASAP7_75t_L g1782 ( 
.A1(n_1706),
.A2(n_803),
.B(n_802),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1713),
.Y(n_1783)
);

AO21x2_ASAP7_75t_L g1784 ( 
.A1(n_1705),
.A2(n_1447),
.B(n_1441),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1685),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1751),
.Y(n_1786)
);

NAND2x1p5_ASAP7_75t_L g1787 ( 
.A(n_1678),
.B(n_1590),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1683),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1735),
.A2(n_1445),
.B(n_1380),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1741),
.A2(n_1678),
.B(n_1742),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1708),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_1670),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1714),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1692),
.A2(n_809),
.B(n_807),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1686),
.B(n_1599),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1737),
.B(n_1189),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1725),
.B(n_810),
.Y(n_1797)
);

OA21x2_ASAP7_75t_L g1798 ( 
.A1(n_1676),
.A2(n_812),
.B(n_811),
.Y(n_1798)
);

INVx8_ASAP7_75t_L g1799 ( 
.A(n_1670),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1728),
.B(n_815),
.Y(n_1800)
);

NAND2x1p5_ASAP7_75t_L g1801 ( 
.A(n_1700),
.B(n_1599),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1676),
.A2(n_818),
.B(n_816),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1672),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1715),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1742),
.A2(n_1445),
.B(n_1496),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1694),
.A2(n_1695),
.B(n_1688),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1675),
.A2(n_1431),
.B1(n_488),
.B2(n_492),
.Y(n_1807)
);

OR2x6_ASAP7_75t_L g1808 ( 
.A(n_1672),
.B(n_1707),
.Y(n_1808)
);

OA21x2_ASAP7_75t_L g1809 ( 
.A1(n_1713),
.A2(n_827),
.B(n_825),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1715),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1689),
.B(n_1599),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1672),
.B(n_479),
.Y(n_1812)
);

AO21x2_ASAP7_75t_L g1813 ( 
.A1(n_1717),
.A2(n_1366),
.B(n_1330),
.Y(n_1813)
);

OA21x2_ASAP7_75t_L g1814 ( 
.A1(n_1709),
.A2(n_492),
.B(n_488),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1693),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1728),
.B(n_502),
.Y(n_1816)
);

AOI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1718),
.A2(n_1431),
.B(n_1384),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1689),
.B(n_502),
.Y(n_1818)
);

AOI222xp33_ASAP7_75t_L g1819 ( 
.A1(n_1690),
.A2(n_555),
.B1(n_533),
.B2(n_562),
.C1(n_539),
.C2(n_531),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1689),
.B(n_1599),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1715),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1715),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1681),
.B(n_1695),
.Y(n_1823)
);

BUFx10_ASAP7_75t_L g1824 ( 
.A(n_1669),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1746),
.Y(n_1825)
);

BUFx12f_ASAP7_75t_L g1826 ( 
.A(n_1677),
.Y(n_1826)
);

AO21x2_ASAP7_75t_L g1827 ( 
.A1(n_1717),
.A2(n_533),
.B(n_531),
.Y(n_1827)
);

OAI21x1_ASAP7_75t_L g1828 ( 
.A1(n_1709),
.A2(n_1540),
.B(n_1527),
.Y(n_1828)
);

OA21x2_ASAP7_75t_L g1829 ( 
.A1(n_1704),
.A2(n_1740),
.B(n_1736),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1727),
.B(n_539),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1703),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1704),
.Y(n_1832)
);

AOI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1684),
.A2(n_562),
.B(n_567),
.C(n_555),
.Y(n_1833)
);

AOI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1718),
.A2(n_568),
.B(n_567),
.Y(n_1834)
);

CKINVDCx20_ASAP7_75t_R g1835 ( 
.A(n_1720),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1691),
.A2(n_1287),
.B(n_1315),
.Y(n_1836)
);

BUFx2_ASAP7_75t_L g1837 ( 
.A(n_1746),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1700),
.B(n_1599),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1736),
.A2(n_1450),
.B(n_1430),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1734),
.B(n_1348),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1674),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1746),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1744),
.B(n_568),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1722),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1698),
.B(n_571),
.Y(n_1845)
);

A2O1A1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1716),
.A2(n_572),
.B(n_574),
.C(n_571),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1687),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1722),
.Y(n_1848)
);

INVx4_ASAP7_75t_SL g1849 ( 
.A(n_1703),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1698),
.B(n_572),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1716),
.B(n_574),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1701),
.B(n_1470),
.Y(n_1852)
);

BUFx3_ASAP7_75t_L g1853 ( 
.A(n_1703),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1687),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1699),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1697),
.B(n_579),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1711),
.B(n_1444),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1740),
.A2(n_1474),
.B(n_1395),
.Y(n_1858)
);

AO31x2_ASAP7_75t_L g1859 ( 
.A1(n_1699),
.A2(n_582),
.A3(n_583),
.B(n_579),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1727),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1688),
.Y(n_1861)
);

AOI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1718),
.A2(n_1727),
.B(n_1743),
.Y(n_1862)
);

AOI21x1_ASAP7_75t_L g1863 ( 
.A1(n_1738),
.A2(n_583),
.B(n_582),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1750),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1701),
.B(n_1394),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1745),
.Y(n_1866)
);

AOI21xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1729),
.A2(n_590),
.B(n_588),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1745),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1702),
.Y(n_1869)
);

AOI21x1_ASAP7_75t_L g1870 ( 
.A1(n_1702),
.A2(n_590),
.B(n_588),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1721),
.Y(n_1871)
);

INVx3_ASAP7_75t_L g1872 ( 
.A(n_1750),
.Y(n_1872)
);

OAI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1723),
.A2(n_1399),
.B(n_1395),
.Y(n_1873)
);

OAI21x1_ASAP7_75t_L g1874 ( 
.A1(n_1723),
.A2(n_1406),
.B(n_1399),
.Y(n_1874)
);

AO31x2_ASAP7_75t_L g1875 ( 
.A1(n_1750),
.A2(n_624),
.A3(n_628),
.B(n_623),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1697),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1691),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1739),
.Y(n_1878)
);

BUFx8_ASAP7_75t_L g1879 ( 
.A(n_1667),
.Y(n_1879)
);

INVxp67_ASAP7_75t_L g1880 ( 
.A(n_1747),
.Y(n_1880)
);

OA21x2_ASAP7_75t_L g1881 ( 
.A1(n_1739),
.A2(n_624),
.B(n_623),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1719),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1668),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1666),
.A2(n_1415),
.B(n_1413),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1686),
.B(n_628),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1703),
.Y(n_1886)
);

INVx4_ASAP7_75t_L g1887 ( 
.A(n_1703),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1733),
.A2(n_1389),
.B(n_1372),
.Y(n_1888)
);

BUFx8_ASAP7_75t_L g1889 ( 
.A(n_1693),
.Y(n_1889)
);

NAND2x1p5_ASAP7_75t_L g1890 ( 
.A(n_1678),
.B(n_1389),
.Y(n_1890)
);

AOI21x1_ASAP7_75t_L g1891 ( 
.A1(n_1673),
.A2(n_634),
.B(n_633),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1686),
.B(n_1415),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1668),
.Y(n_1893)
);

NAND2x1p5_ASAP7_75t_L g1894 ( 
.A(n_1678),
.B(n_1389),
.Y(n_1894)
);

INVx3_ASAP7_75t_L g1895 ( 
.A(n_1696),
.Y(n_1895)
);

AO31x2_ASAP7_75t_L g1896 ( 
.A1(n_1710),
.A2(n_634),
.A3(n_641),
.B(n_633),
.Y(n_1896)
);

OAI21x1_ASAP7_75t_L g1897 ( 
.A1(n_1666),
.A2(n_1434),
.B(n_1427),
.Y(n_1897)
);

OAI21x1_ASAP7_75t_L g1898 ( 
.A1(n_1666),
.A2(n_1434),
.B(n_1427),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1854),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1808),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1847),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1871),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1847),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1760),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1788),
.B(n_641),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1763),
.B(n_644),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1855),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1765),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1804),
.B(n_644),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1855),
.Y(n_1910)
);

INVx3_ASAP7_75t_L g1911 ( 
.A(n_1757),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1769),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1883),
.Y(n_1913)
);

HB1xp67_ASAP7_75t_L g1914 ( 
.A(n_1791),
.Y(n_1914)
);

OAI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1880),
.A2(n_646),
.B(n_645),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1893),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1803),
.B(n_645),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1803),
.B(n_1768),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1775),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1786),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1793),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1779),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1776),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_1844),
.Y(n_1924)
);

BUFx8_ASAP7_75t_SL g1925 ( 
.A(n_1792),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1832),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1810),
.B(n_646),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1848),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1806),
.A2(n_658),
.B(n_657),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1785),
.Y(n_1930)
);

HB1xp67_ASAP7_75t_L g1931 ( 
.A(n_1780),
.Y(n_1931)
);

AO21x2_ASAP7_75t_L g1932 ( 
.A1(n_1806),
.A2(n_658),
.B(n_657),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1866),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1843),
.B(n_662),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1783),
.Y(n_1935)
);

INVx3_ASAP7_75t_L g1936 ( 
.A(n_1757),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1821),
.B(n_662),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1822),
.B(n_674),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1783),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1868),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1880),
.B(n_674),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1808),
.B(n_694),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1813),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1896),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1896),
.Y(n_1945)
);

AO21x2_ASAP7_75t_L g1946 ( 
.A1(n_1823),
.A2(n_694),
.B(n_1446),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1825),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1813),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1851),
.B(n_1818),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1808),
.B(n_690),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1896),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1859),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1859),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1859),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1837),
.Y(n_1955)
);

NAND2x1p5_ASAP7_75t_L g1956 ( 
.A(n_1809),
.B(n_1759),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1757),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1860),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1889),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1841),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1757),
.Y(n_1961)
);

HB1xp67_ASAP7_75t_L g1962 ( 
.A(n_1816),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1764),
.B(n_580),
.Y(n_1963)
);

AOI22xp33_ASAP7_75t_SL g1964 ( 
.A1(n_1857),
.A2(n_619),
.B1(n_589),
.B2(n_629),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1816),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1754),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1771),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1771),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1771),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1752),
.B(n_0),
.Y(n_1970)
);

OAI21xp5_ASAP7_75t_L g1971 ( 
.A1(n_1891),
.A2(n_1287),
.B(n_1315),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1771),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1812),
.Y(n_1973)
);

INVx3_ASAP7_75t_L g1974 ( 
.A(n_1829),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1823),
.B(n_1),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1797),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1752),
.B(n_1),
.Y(n_1977)
);

HB1xp67_ASAP7_75t_L g1978 ( 
.A(n_1797),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1800),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1829),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1814),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1814),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1800),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1809),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1862),
.B(n_2),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1772),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1782),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1796),
.B(n_586),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1787),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1759),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1876),
.B(n_2),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1772),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1830),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1830),
.Y(n_1994)
);

BUFx6f_ASAP7_75t_L g1995 ( 
.A(n_1831),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1773),
.A2(n_1466),
.B(n_1454),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1885),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1782),
.Y(n_1998)
);

INVx2_ASAP7_75t_L g1999 ( 
.A(n_1861),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1861),
.Y(n_2000)
);

OAI21x1_ASAP7_75t_L g2001 ( 
.A1(n_1790),
.A2(n_1473),
.B(n_1426),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1869),
.Y(n_2002)
);

BUFx3_ASAP7_75t_L g2003 ( 
.A(n_1889),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1754),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1869),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1787),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1875),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1875),
.Y(n_2008)
);

AND2x4_ASAP7_75t_L g2009 ( 
.A(n_1849),
.B(n_203),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1756),
.Y(n_2010)
);

INVx4_ASAP7_75t_L g2011 ( 
.A(n_1849),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1890),
.Y(n_2012)
);

OA21x2_ASAP7_75t_L g2013 ( 
.A1(n_1790),
.A2(n_885),
.B(n_879),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1811),
.B(n_3),
.Y(n_2014)
);

INVxp67_ASAP7_75t_SL g2015 ( 
.A(n_1890),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1875),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1758),
.Y(n_2017)
);

AOI21xp5_ASAP7_75t_L g2018 ( 
.A1(n_1888),
.A2(n_1426),
.B(n_1417),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1811),
.B(n_3),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1758),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1894),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1756),
.Y(n_2022)
);

INVx3_ASAP7_75t_SL g2023 ( 
.A(n_1767),
.Y(n_2023)
);

INVx2_ASAP7_75t_SL g2024 ( 
.A(n_1831),
.Y(n_2024)
);

BUFx2_ASAP7_75t_L g2025 ( 
.A(n_1761),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1762),
.B(n_7),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1894),
.Y(n_2027)
);

OAI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1857),
.A2(n_1287),
.B(n_1315),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1845),
.B(n_587),
.Y(n_2029)
);

OAI21x1_ASAP7_75t_L g2030 ( 
.A1(n_1870),
.A2(n_1426),
.B(n_1417),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1820),
.B(n_7),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1849),
.B(n_207),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1798),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1820),
.B(n_10),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1766),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1831),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1766),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1850),
.B(n_591),
.Y(n_2038)
);

HB1xp67_ASAP7_75t_L g2039 ( 
.A(n_1761),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1798),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1827),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1856),
.B(n_1795),
.Y(n_2042)
);

OA21x2_ASAP7_75t_L g2043 ( 
.A1(n_1789),
.A2(n_885),
.B(n_879),
.Y(n_2043)
);

CKINVDCx20_ASAP7_75t_R g2044 ( 
.A(n_1925),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1904),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1971),
.A2(n_1774),
.B(n_1833),
.Y(n_2046)
);

NAND3xp33_ASAP7_75t_L g2047 ( 
.A(n_1964),
.B(n_1819),
.C(n_1846),
.Y(n_2047)
);

NAND2xp33_ASAP7_75t_L g2048 ( 
.A(n_2023),
.B(n_1767),
.Y(n_2048)
);

BUFx12f_ASAP7_75t_L g2049 ( 
.A(n_1959),
.Y(n_2049)
);

OAI21x1_ASAP7_75t_L g2050 ( 
.A1(n_1974),
.A2(n_1817),
.B(n_1794),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2028),
.A2(n_1840),
.B1(n_1877),
.B2(n_1878),
.Y(n_2051)
);

OAI33xp33_ASAP7_75t_L g2052 ( 
.A1(n_1941),
.A2(n_612),
.A3(n_603),
.B1(n_616),
.B2(n_604),
.B3(n_600),
.Y(n_2052)
);

OA21x2_ASAP7_75t_L g2053 ( 
.A1(n_1980),
.A2(n_2005),
.B(n_1999),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1928),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1915),
.A2(n_1778),
.B1(n_1807),
.B2(n_1774),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1947),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1922),
.B(n_1815),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1978),
.B(n_1784),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1959),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1922),
.B(n_1767),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1904),
.Y(n_2061)
);

AOI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1931),
.A2(n_1882),
.B1(n_1879),
.B2(n_1840),
.Y(n_2062)
);

INVx2_ASAP7_75t_SL g2063 ( 
.A(n_2023),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_L g2064 ( 
.A1(n_1985),
.A2(n_1879),
.B1(n_1778),
.B2(n_1819),
.Y(n_2064)
);

AOI22xp33_ASAP7_75t_L g2065 ( 
.A1(n_1985),
.A2(n_1836),
.B1(n_1807),
.B2(n_1881),
.Y(n_2065)
);

HB1xp67_ASAP7_75t_L g2066 ( 
.A(n_1914),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_2023),
.B(n_1826),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1918),
.B(n_1853),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1975),
.A2(n_1755),
.B1(n_1846),
.B2(n_1881),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1928),
.Y(n_2070)
);

OAI21x1_ASAP7_75t_L g2071 ( 
.A1(n_1974),
.A2(n_1789),
.B(n_1834),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_1921),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1918),
.B(n_1824),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1908),
.Y(n_2074)
);

OAI21x1_ASAP7_75t_L g2075 ( 
.A1(n_1974),
.A2(n_1770),
.B(n_1777),
.Y(n_2075)
);

INVx3_ASAP7_75t_SL g2076 ( 
.A(n_1959),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1908),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1902),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1912),
.Y(n_2079)
);

AOI22xp33_ASAP7_75t_L g2080 ( 
.A1(n_1973),
.A2(n_1836),
.B1(n_1887),
.B2(n_1886),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1947),
.B(n_1824),
.Y(n_2081)
);

OAI22xp5_ASAP7_75t_L g2082 ( 
.A1(n_1975),
.A2(n_1755),
.B1(n_1792),
.B2(n_1863),
.Y(n_2082)
);

OR2x2_ASAP7_75t_SL g2083 ( 
.A(n_1990),
.B(n_1799),
.Y(n_2083)
);

OAI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_2026),
.A2(n_1886),
.B1(n_1887),
.B2(n_1805),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1947),
.B(n_1842),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1928),
.Y(n_2086)
);

BUFx8_ASAP7_75t_L g2087 ( 
.A(n_2003),
.Y(n_2087)
);

OAI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_2026),
.A2(n_1805),
.B1(n_1799),
.B2(n_1835),
.Y(n_2088)
);

INVx3_ASAP7_75t_L g2089 ( 
.A(n_1955),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1912),
.Y(n_2090)
);

AOI22xp5_ASAP7_75t_L g2091 ( 
.A1(n_1942),
.A2(n_1835),
.B1(n_1784),
.B2(n_1781),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1913),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_L g2093 ( 
.A1(n_1949),
.A2(n_1942),
.B1(n_1900),
.B2(n_1997),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_1900),
.A2(n_1799),
.B1(n_619),
.B2(n_589),
.Y(n_2094)
);

OAI211xp5_ASAP7_75t_L g2095 ( 
.A1(n_2017),
.A2(n_1867),
.B(n_620),
.C(n_622),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1955),
.B(n_1842),
.Y(n_2096)
);

AOI22xp33_ASAP7_75t_L g2097 ( 
.A1(n_1997),
.A2(n_1827),
.B1(n_1892),
.B2(n_629),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_1929),
.A2(n_1888),
.B(n_1753),
.Y(n_2098)
);

AOI221xp5_ASAP7_75t_L g2099 ( 
.A1(n_1934),
.A2(n_639),
.B1(n_642),
.B2(n_637),
.C(n_618),
.Y(n_2099)
);

AO21x2_ASAP7_75t_L g2100 ( 
.A1(n_1929),
.A2(n_1762),
.B(n_1753),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1976),
.B(n_1864),
.Y(n_2101)
);

INVx5_ASAP7_75t_SL g2102 ( 
.A(n_2009),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1913),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1916),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1976),
.B(n_1864),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_2003),
.Y(n_2106)
);

OR2x6_ASAP7_75t_L g2107 ( 
.A(n_1956),
.B(n_1801),
.Y(n_2107)
);

AOI22xp33_ASAP7_75t_L g2108 ( 
.A1(n_2042),
.A2(n_1892),
.B1(n_1315),
.B2(n_1795),
.Y(n_2108)
);

INVxp67_ASAP7_75t_SL g2109 ( 
.A(n_1962),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1955),
.B(n_1872),
.Y(n_2110)
);

AOI222xp33_ASAP7_75t_L g2111 ( 
.A1(n_1988),
.A2(n_659),
.B1(n_647),
.B2(n_660),
.C1(n_656),
.C2(n_643),
.Y(n_2111)
);

AO21x2_ASAP7_75t_L g2112 ( 
.A1(n_1929),
.A2(n_1897),
.B(n_1884),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1916),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1919),
.Y(n_2114)
);

AOI222xp33_ASAP7_75t_L g2115 ( 
.A1(n_2029),
.A2(n_671),
.B1(n_668),
.B2(n_672),
.C1(n_670),
.C2(n_663),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2010),
.B(n_1872),
.Y(n_2116)
);

OAI21x1_ASAP7_75t_L g2117 ( 
.A1(n_1974),
.A2(n_1898),
.B(n_1802),
.Y(n_2117)
);

OA21x2_ASAP7_75t_L g2118 ( 
.A1(n_1980),
.A2(n_1828),
.B(n_1839),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_1929),
.A2(n_1802),
.B(n_1852),
.Y(n_2119)
);

AOI22xp33_ASAP7_75t_L g2120 ( 
.A1(n_2042),
.A2(n_2020),
.B1(n_2035),
.B2(n_2017),
.Y(n_2120)
);

OAI22xp5_ASAP7_75t_L g2121 ( 
.A1(n_2003),
.A2(n_1801),
.B1(n_1852),
.B2(n_1865),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_1966),
.Y(n_2122)
);

AO21x2_ASAP7_75t_L g2123 ( 
.A1(n_1932),
.A2(n_1858),
.B(n_1873),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2020),
.A2(n_1315),
.B1(n_1865),
.B2(n_1838),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1993),
.B(n_1895),
.Y(n_2125)
);

BUFx2_ASAP7_75t_L g2126 ( 
.A(n_1966),
.Y(n_2126)
);

OAI211xp5_ASAP7_75t_L g2127 ( 
.A1(n_2035),
.A2(n_678),
.B(n_684),
.C(n_673),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2039),
.B(n_1895),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1923),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2004),
.B(n_1838),
.Y(n_2130)
);

AOI22xp33_ASAP7_75t_L g2131 ( 
.A1(n_2037),
.A2(n_1222),
.B1(n_1204),
.B2(n_687),
.Y(n_2131)
);

BUFx12f_ASAP7_75t_L g2132 ( 
.A(n_1917),
.Y(n_2132)
);

AOI22xp33_ASAP7_75t_L g2133 ( 
.A1(n_2037),
.A2(n_1222),
.B1(n_1204),
.B2(n_688),
.Y(n_2133)
);

AOI22xp33_ASAP7_75t_L g2134 ( 
.A1(n_1965),
.A2(n_1222),
.B1(n_1204),
.B2(n_691),
.Y(n_2134)
);

NAND3xp33_ASAP7_75t_L g2135 ( 
.A(n_1993),
.B(n_692),
.C(n_686),
.Y(n_2135)
);

BUFx4f_ASAP7_75t_SL g2136 ( 
.A(n_1995),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_1924),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_1901),
.B(n_1874),
.Y(n_2138)
);

BUFx2_ASAP7_75t_L g2139 ( 
.A(n_2004),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_1917),
.A2(n_1204),
.B1(n_1222),
.B2(n_693),
.Y(n_2140)
);

AOI221xp5_ASAP7_75t_L g2141 ( 
.A1(n_2038),
.A2(n_493),
.B1(n_498),
.B2(n_490),
.C(n_489),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1923),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1919),
.Y(n_2143)
);

AOI221xp5_ASAP7_75t_L g2144 ( 
.A1(n_1905),
.A2(n_506),
.B1(n_515),
.B2(n_505),
.C(n_500),
.Y(n_2144)
);

AOI22xp33_ASAP7_75t_L g2145 ( 
.A1(n_1994),
.A2(n_1222),
.B1(n_1204),
.B2(n_528),
.Y(n_2145)
);

INVx3_ASAP7_75t_L g2146 ( 
.A(n_2010),
.Y(n_2146)
);

AOI22xp33_ASAP7_75t_L g2147 ( 
.A1(n_1994),
.A2(n_530),
.B1(n_535),
.B2(n_516),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1935),
.B(n_12),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_1950),
.A2(n_542),
.B1(n_545),
.B2(n_540),
.Y(n_2149)
);

NAND2x1_ASAP7_75t_L g2150 ( 
.A(n_2010),
.B(n_1417),
.Y(n_2150)
);

NOR2xp67_ASAP7_75t_L g2151 ( 
.A(n_1960),
.B(n_14),
.Y(n_2151)
);

OAI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1956),
.A2(n_556),
.B1(n_557),
.B2(n_551),
.Y(n_2152)
);

OR2x6_ASAP7_75t_L g2153 ( 
.A(n_1956),
.B(n_892),
.Y(n_2153)
);

OAI22xp33_ASAP7_75t_L g2154 ( 
.A1(n_2011),
.A2(n_564),
.B1(n_566),
.B2(n_561),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1950),
.A2(n_584),
.B1(n_585),
.B2(n_577),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_1919),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1930),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1930),
.Y(n_2158)
);

AND2x4_ASAP7_75t_L g2159 ( 
.A(n_2010),
.B(n_14),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2009),
.A2(n_609),
.B1(n_610),
.B2(n_593),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1920),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_1901),
.B(n_1903),
.Y(n_2162)
);

AOI31xp33_ASAP7_75t_L g2163 ( 
.A1(n_2014),
.A2(n_2031),
.A3(n_2034),
.B(n_2019),
.Y(n_2163)
);

AOI33xp33_ASAP7_75t_L g2164 ( 
.A1(n_1905),
.A2(n_15),
.A3(n_16),
.B1(n_17),
.B2(n_18),
.B3(n_19),
.Y(n_2164)
);

AOI22xp33_ASAP7_75t_SL g2165 ( 
.A1(n_1932),
.A2(n_615),
.B1(n_617),
.B2(n_614),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1920),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1958),
.Y(n_2167)
);

AOI21xp5_ASAP7_75t_L g2168 ( 
.A1(n_1932),
.A2(n_2018),
.B(n_2015),
.Y(n_2168)
);

AOI22xp33_ASAP7_75t_L g2169 ( 
.A1(n_1932),
.A2(n_2032),
.B1(n_2009),
.B2(n_1983),
.Y(n_2169)
);

AOI22xp33_ASAP7_75t_L g2170 ( 
.A1(n_2009),
.A2(n_2032),
.B1(n_1983),
.B2(n_1979),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_1963),
.A2(n_631),
.B1(n_636),
.B2(n_630),
.C(n_621),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1958),
.Y(n_2172)
);

AOI22xp33_ASAP7_75t_SL g2173 ( 
.A1(n_2014),
.A2(n_652),
.B1(n_655),
.B2(n_648),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_2032),
.A2(n_665),
.B1(n_666),
.B2(n_664),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1899),
.Y(n_2175)
);

NAND2x1_ASAP7_75t_L g2176 ( 
.A(n_2022),
.B(n_1435),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_2032),
.A2(n_669),
.B1(n_677),
.B2(n_667),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_1935),
.B(n_15),
.Y(n_2178)
);

AOI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_1979),
.A2(n_695),
.B1(n_696),
.B2(n_680),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_1986),
.A2(n_895),
.B1(n_897),
.B2(n_892),
.Y(n_2180)
);

NOR2x1_ASAP7_75t_SL g2181 ( 
.A(n_1946),
.B(n_1184),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_1986),
.A2(n_897),
.B1(n_902),
.B2(n_895),
.Y(n_2182)
);

AOI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_1992),
.A2(n_1970),
.B1(n_1977),
.B2(n_2019),
.Y(n_2183)
);

BUFx2_ASAP7_75t_L g2184 ( 
.A(n_2025),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1920),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1899),
.Y(n_2186)
);

AO31x2_ASAP7_75t_L g2187 ( 
.A1(n_1967),
.A2(n_905),
.A3(n_908),
.B(n_902),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_1946),
.A2(n_1442),
.B(n_1435),
.Y(n_2188)
);

AOI22xp33_ASAP7_75t_SL g2189 ( 
.A1(n_2031),
.A2(n_1184),
.B1(n_18),
.B2(n_16),
.Y(n_2189)
);

AOI222xp33_ASAP7_75t_L g2190 ( 
.A1(n_1970),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.C1(n_21),
.C2(n_22),
.Y(n_2190)
);

AOI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_1977),
.A2(n_908),
.B1(n_905),
.B2(n_1297),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_1906),
.Y(n_2192)
);

O2A1O1Ixp5_ASAP7_75t_L g2193 ( 
.A1(n_1960),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_2193)
);

AOI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_1992),
.A2(n_917),
.B1(n_866),
.B2(n_877),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2034),
.A2(n_917),
.B1(n_866),
.B2(n_877),
.Y(n_2195)
);

OAI221xp5_ASAP7_75t_L g2196 ( 
.A1(n_1909),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.C(n_27),
.Y(n_2196)
);

AOI21xp5_ASAP7_75t_L g2197 ( 
.A1(n_2013),
.A2(n_2043),
.B(n_2001),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2126),
.B(n_2139),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2184),
.B(n_2025),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2053),
.Y(n_2200)
);

OR2x2_ASAP7_75t_L g2201 ( 
.A(n_2058),
.B(n_1999),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2053),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2054),
.Y(n_2203)
);

INVx1_ASAP7_75t_SL g2204 ( 
.A(n_2044),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2070),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2107),
.B(n_1999),
.Y(n_2206)
);

AND2x2_ASAP7_75t_L g2207 ( 
.A(n_2056),
.B(n_1989),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2058),
.B(n_2005),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2109),
.B(n_1927),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_2066),
.Y(n_2210)
);

HB1xp67_ASAP7_75t_L g2211 ( 
.A(n_2137),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2120),
.B(n_2192),
.Y(n_2212)
);

NAND2x1_ASAP7_75t_L g2213 ( 
.A(n_2107),
.B(n_1989),
.Y(n_2213)
);

AND2x4_ASAP7_75t_L g2214 ( 
.A(n_2107),
.B(n_2005),
.Y(n_2214)
);

CKINVDCx5p33_ASAP7_75t_R g2215 ( 
.A(n_2049),
.Y(n_2215)
);

OAI21xp5_ASAP7_75t_L g2216 ( 
.A1(n_2047),
.A2(n_1991),
.B(n_1937),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2086),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2167),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2172),
.Y(n_2219)
);

INVxp67_ASAP7_75t_SL g2220 ( 
.A(n_2072),
.Y(n_2220)
);

INVxp33_ASAP7_75t_SL g2221 ( 
.A(n_2067),
.Y(n_2221)
);

INVx2_ASAP7_75t_SL g2222 ( 
.A(n_2059),
.Y(n_2222)
);

AND2x2_ASAP7_75t_L g2223 ( 
.A(n_2056),
.B(n_1989),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2045),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2083),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_2162),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2089),
.B(n_1989),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2089),
.B(n_2057),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2130),
.B(n_2022),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2175),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2186),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2061),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2114),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2073),
.B(n_2022),
.Y(n_2234)
);

INVx1_ASAP7_75t_SL g2235 ( 
.A(n_2076),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2074),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2143),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2122),
.B(n_2022),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2077),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_2146),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2156),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2122),
.B(n_2006),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2079),
.Y(n_2243)
);

AOI22xp33_ASAP7_75t_L g2244 ( 
.A1(n_2055),
.A2(n_2007),
.B1(n_2016),
.B2(n_2008),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_2125),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2161),
.Y(n_2246)
);

BUFx2_ASAP7_75t_L g2247 ( 
.A(n_2132),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2068),
.B(n_2085),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2166),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2078),
.B(n_1927),
.Y(n_2250)
);

AOI22xp33_ASAP7_75t_L g2251 ( 
.A1(n_2055),
.A2(n_2007),
.B1(n_2016),
.B2(n_2008),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_2125),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_2101),
.B(n_2000),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2090),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2096),
.B(n_2006),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2081),
.B(n_2006),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2185),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_2101),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_2064),
.A2(n_1995),
.B1(n_2011),
.B2(n_1991),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2105),
.B(n_1937),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2146),
.B(n_2000),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2092),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2046),
.A2(n_1995),
.B1(n_2011),
.B2(n_1946),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2103),
.Y(n_2264)
);

INVx3_ASAP7_75t_L g2265 ( 
.A(n_2116),
.Y(n_2265)
);

AND2x4_ASAP7_75t_L g2266 ( 
.A(n_2063),
.B(n_2116),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2104),
.Y(n_2267)
);

OAI22xp5_ASAP7_75t_L g2268 ( 
.A1(n_2051),
.A2(n_2011),
.B1(n_1938),
.B2(n_1909),
.Y(n_2268)
);

HB1xp67_ASAP7_75t_L g2269 ( 
.A(n_2105),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2082),
.A2(n_1995),
.B1(n_1946),
.B2(n_2012),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2183),
.B(n_1938),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2113),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2138),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_2110),
.B(n_2002),
.Y(n_2274)
);

INVxp33_ASAP7_75t_L g2275 ( 
.A(n_2181),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2129),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2069),
.A2(n_2024),
.B1(n_2036),
.B2(n_1995),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2128),
.B(n_2002),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2110),
.B(n_1939),
.Y(n_2279)
);

INVxp67_ASAP7_75t_SL g2280 ( 
.A(n_2151),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2093),
.B(n_2091),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2060),
.B(n_1939),
.Y(n_2282)
);

INVxp67_ASAP7_75t_SL g2283 ( 
.A(n_2148),
.Y(n_2283)
);

INVx2_ASAP7_75t_SL g2284 ( 
.A(n_2059),
.Y(n_2284)
);

HB1xp67_ASAP7_75t_L g2285 ( 
.A(n_2142),
.Y(n_2285)
);

NAND3xp33_ASAP7_75t_L g2286 ( 
.A(n_2111),
.B(n_1945),
.C(n_1944),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2157),
.Y(n_2287)
);

INVx2_ASAP7_75t_L g2288 ( 
.A(n_2158),
.Y(n_2288)
);

CKINVDCx5p33_ASAP7_75t_R g2289 ( 
.A(n_2087),
.Y(n_2289)
);

INVxp67_ASAP7_75t_SL g2290 ( 
.A(n_2148),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2082),
.A2(n_1995),
.B1(n_2021),
.B2(n_2012),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2178),
.Y(n_2292)
);

BUFx2_ASAP7_75t_L g2293 ( 
.A(n_2087),
.Y(n_2293)
);

OAI21xp5_ASAP7_75t_SL g2294 ( 
.A1(n_2111),
.A2(n_2036),
.B(n_2024),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2106),
.B(n_1901),
.Y(n_2295)
);

INVxp67_ASAP7_75t_SL g2296 ( 
.A(n_2178),
.Y(n_2296)
);

BUFx3_ASAP7_75t_L g2297 ( 
.A(n_2059),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2170),
.B(n_1903),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2153),
.B(n_1903),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2088),
.B(n_1907),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2069),
.A2(n_2041),
.B1(n_2021),
.B2(n_2027),
.Y(n_2301)
);

OAI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2065),
.A2(n_2021),
.B1(n_2027),
.B2(n_2012),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2118),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2071),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2153),
.B(n_1907),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2169),
.A2(n_2027),
.B1(n_2041),
.B2(n_1945),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_2153),
.B(n_1926),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_SL g2308 ( 
.A1(n_2196),
.A2(n_2013),
.B1(n_1951),
.B2(n_1944),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2121),
.Y(n_2309)
);

OAI221xp5_ASAP7_75t_SL g2310 ( 
.A1(n_2164),
.A2(n_1951),
.B1(n_1952),
.B2(n_1954),
.C(n_1953),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2121),
.Y(n_2311)
);

INVxp67_ASAP7_75t_L g2312 ( 
.A(n_2159),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2163),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2102),
.B(n_1907),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2084),
.B(n_1910),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2080),
.B(n_1910),
.Y(n_2316)
);

INVxp67_ASAP7_75t_SL g2317 ( 
.A(n_2159),
.Y(n_2317)
);

HB1xp67_ASAP7_75t_L g2318 ( 
.A(n_2150),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2163),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_L g2320 ( 
.A1(n_2190),
.A2(n_1953),
.B1(n_1954),
.B2(n_1952),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_2136),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2190),
.A2(n_1982),
.B1(n_1981),
.B2(n_1972),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2118),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2232),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2200),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_L g2326 ( 
.A(n_2283),
.B(n_2062),
.Y(n_2326)
);

OR2x2_ASAP7_75t_L g2327 ( 
.A(n_2313),
.B(n_2168),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2290),
.B(n_2191),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2228),
.B(n_2256),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2200),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2232),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2236),
.Y(n_2332)
);

AND2x4_ASAP7_75t_L g2333 ( 
.A(n_2225),
.B(n_2050),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2296),
.B(n_2292),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2202),
.Y(n_2335)
);

AND2x4_ASAP7_75t_L g2336 ( 
.A(n_2225),
.B(n_1926),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2236),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2202),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2221),
.B(n_2052),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2303),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2210),
.B(n_2102),
.Y(n_2341)
);

NOR2xp67_ASAP7_75t_L g2342 ( 
.A(n_2319),
.B(n_2098),
.Y(n_2342)
);

OR2x2_ASAP7_75t_L g2343 ( 
.A(n_2316),
.B(n_1910),
.Y(n_2343)
);

OAI21xp33_ASAP7_75t_SL g2344 ( 
.A1(n_2280),
.A2(n_2152),
.B(n_2094),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2221),
.B(n_2127),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2228),
.B(n_2256),
.Y(n_2346)
);

BUFx3_ASAP7_75t_L g2347 ( 
.A(n_2293),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2266),
.B(n_2102),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2239),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2239),
.Y(n_2350)
);

INVxp67_ASAP7_75t_SL g2351 ( 
.A(n_2323),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2266),
.B(n_2048),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2272),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2265),
.B(n_1926),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2266),
.B(n_2234),
.Y(n_2355)
);

INVx3_ASAP7_75t_L g2356 ( 
.A(n_2213),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2285),
.Y(n_2357)
);

OAI21xp33_ASAP7_75t_L g2358 ( 
.A1(n_2244),
.A2(n_2196),
.B(n_2115),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2272),
.Y(n_2359)
);

AND2x2_ASAP7_75t_L g2360 ( 
.A(n_2234),
.B(n_2108),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2287),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2260),
.B(n_2100),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2248),
.B(n_2124),
.Y(n_2363)
);

BUFx2_ASAP7_75t_L g2364 ( 
.A(n_2293),
.Y(n_2364)
);

INVxp67_ASAP7_75t_SL g2365 ( 
.A(n_2323),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2303),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2287),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2218),
.Y(n_2368)
);

HB1xp67_ASAP7_75t_L g2369 ( 
.A(n_2211),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2251),
.B(n_2152),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2212),
.B(n_2097),
.Y(n_2371)
);

BUFx2_ASAP7_75t_SL g2372 ( 
.A(n_2235),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2220),
.B(n_2119),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2219),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2224),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2243),
.Y(n_2376)
);

OAI221xp5_ASAP7_75t_L g2377 ( 
.A1(n_2294),
.A2(n_2189),
.B1(n_2115),
.B2(n_2099),
.C(n_2171),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2300),
.B(n_2100),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2248),
.B(n_1933),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2222),
.B(n_2284),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2254),
.Y(n_2381)
);

NAND3xp33_ASAP7_75t_L g2382 ( 
.A(n_2270),
.B(n_2165),
.C(n_2099),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2309),
.B(n_1933),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2265),
.B(n_1933),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_2261),
.Y(n_2385)
);

INVx2_ASAP7_75t_SL g2386 ( 
.A(n_2289),
.Y(n_2386)
);

HB1xp67_ASAP7_75t_L g2387 ( 
.A(n_2276),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2271),
.B(n_2245),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2311),
.B(n_1940),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2209),
.B(n_1940),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2252),
.B(n_2135),
.Y(n_2391)
);

OR2x2_ASAP7_75t_L g2392 ( 
.A(n_2315),
.B(n_1940),
.Y(n_2392)
);

HB1xp67_ASAP7_75t_L g2393 ( 
.A(n_2276),
.Y(n_2393)
);

INVxp67_ASAP7_75t_SL g2394 ( 
.A(n_2201),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2282),
.B(n_1899),
.Y(n_2395)
);

OR2x2_ASAP7_75t_L g2396 ( 
.A(n_2250),
.B(n_1967),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2261),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2282),
.B(n_2176),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2262),
.Y(n_2399)
);

AND2x6_ASAP7_75t_SL g2400 ( 
.A(n_2281),
.B(n_2173),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2297),
.B(n_2095),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2264),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2255),
.B(n_1972),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2255),
.B(n_2075),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2267),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2288),
.Y(n_2406)
);

OR2x2_ASAP7_75t_L g2407 ( 
.A(n_2302),
.B(n_2187),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2258),
.B(n_2195),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_2265),
.B(n_1911),
.Y(n_2409)
);

AND2x4_ASAP7_75t_L g2410 ( 
.A(n_2274),
.B(n_1911),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2269),
.B(n_2317),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2216),
.B(n_1981),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2288),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2203),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2298),
.B(n_2312),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2279),
.B(n_1984),
.Y(n_2416)
);

BUFx2_ASAP7_75t_SL g2417 ( 
.A(n_2247),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2298),
.B(n_1981),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_2203),
.Y(n_2419)
);

NAND4xp25_ASAP7_75t_L g2420 ( 
.A(n_2310),
.B(n_2193),
.C(n_2141),
.D(n_2171),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2230),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2230),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2279),
.B(n_1984),
.Y(n_2423)
);

INVxp67_ASAP7_75t_L g2424 ( 
.A(n_2286),
.Y(n_2424)
);

INVx1_ASAP7_75t_SL g2425 ( 
.A(n_2289),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2222),
.B(n_2284),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2231),
.Y(n_2427)
);

AND2x4_ASAP7_75t_SL g2428 ( 
.A(n_2198),
.B(n_2160),
.Y(n_2428)
);

NAND3xp33_ASAP7_75t_L g2429 ( 
.A(n_2301),
.B(n_2141),
.C(n_2144),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2205),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2263),
.B(n_1982),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2231),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2229),
.B(n_1984),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2205),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2217),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2217),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2357),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2347),
.Y(n_2438)
);

NAND2x1p5_ASAP7_75t_L g2439 ( 
.A(n_2356),
.B(n_2213),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2358),
.A2(n_2291),
.B1(n_2275),
.B2(n_2268),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2424),
.B(n_2226),
.Y(n_2441)
);

BUFx6f_ASAP7_75t_L g2442 ( 
.A(n_2347),
.Y(n_2442)
);

AOI22xp33_ASAP7_75t_L g2443 ( 
.A1(n_2424),
.A2(n_2275),
.B1(n_2277),
.B2(n_2308),
.Y(n_2443)
);

OAI221xp5_ASAP7_75t_L g2444 ( 
.A1(n_2344),
.A2(n_2377),
.B1(n_2429),
.B2(n_2420),
.C(n_2370),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2364),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2357),
.Y(n_2446)
);

OAI31xp33_ASAP7_75t_SL g2447 ( 
.A1(n_2377),
.A2(n_2306),
.A3(n_2204),
.B(n_2144),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2369),
.B(n_2226),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2369),
.B(n_2253),
.Y(n_2449)
);

AOI221xp5_ASAP7_75t_L g2450 ( 
.A1(n_2382),
.A2(n_2320),
.B1(n_2322),
.B2(n_2259),
.C(n_2304),
.Y(n_2450)
);

AOI22xp5_ASAP7_75t_L g2451 ( 
.A1(n_2417),
.A2(n_2247),
.B1(n_2321),
.B2(n_2297),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2355),
.Y(n_2452)
);

OR2x2_ASAP7_75t_L g2453 ( 
.A(n_2415),
.B(n_2253),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2352),
.B(n_2314),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2380),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2324),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_2380),
.B(n_2321),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2331),
.Y(n_2458)
);

AOI221xp5_ASAP7_75t_SL g2459 ( 
.A1(n_2371),
.A2(n_2304),
.B1(n_2238),
.B2(n_2198),
.C(n_2314),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_2387),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2332),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2411),
.B(n_2388),
.Y(n_2462)
);

BUFx2_ASAP7_75t_L g2463 ( 
.A(n_2401),
.Y(n_2463)
);

AND2x4_ASAP7_75t_L g2464 ( 
.A(n_2348),
.B(n_2318),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_2372),
.B(n_2207),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2337),
.Y(n_2466)
);

INVx5_ASAP7_75t_L g2467 ( 
.A(n_2386),
.Y(n_2467)
);

AOI22xp33_ASAP7_75t_L g2468 ( 
.A1(n_2345),
.A2(n_2273),
.B1(n_2274),
.B2(n_2215),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2425),
.B(n_2215),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2345),
.A2(n_2273),
.B1(n_2274),
.B2(n_2214),
.Y(n_2470)
);

OAI31xp33_ASAP7_75t_L g2471 ( 
.A1(n_2339),
.A2(n_2154),
.A3(n_2155),
.B(n_2149),
.Y(n_2471)
);

O2A1O1Ixp33_ASAP7_75t_L g2472 ( 
.A1(n_2339),
.A2(n_2208),
.B(n_2201),
.C(n_2206),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2356),
.Y(n_2473)
);

INVx1_ASAP7_75t_SL g2474 ( 
.A(n_2428),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2329),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2349),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2350),
.Y(n_2477)
);

BUFx3_ASAP7_75t_L g2478 ( 
.A(n_2426),
.Y(n_2478)
);

AOI221xp5_ASAP7_75t_L g2479 ( 
.A1(n_2373),
.A2(n_2214),
.B1(n_2206),
.B2(n_2305),
.C(n_2299),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2346),
.B(n_2207),
.Y(n_2480)
);

NAND3xp33_ASAP7_75t_L g2481 ( 
.A(n_2391),
.B(n_2147),
.C(n_2179),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2334),
.B(n_2233),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2336),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2325),
.Y(n_2484)
);

OAI31xp33_ASAP7_75t_SL g2485 ( 
.A1(n_2400),
.A2(n_2206),
.A3(n_2214),
.B(n_2199),
.Y(n_2485)
);

OAI22xp5_ASAP7_75t_L g2486 ( 
.A1(n_2326),
.A2(n_2177),
.B1(n_2174),
.B2(n_2199),
.Y(n_2486)
);

OAI33xp33_ASAP7_75t_L g2487 ( 
.A1(n_2378),
.A2(n_2208),
.A3(n_2249),
.B1(n_2246),
.B2(n_2233),
.B3(n_2237),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2353),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2360),
.B(n_2223),
.Y(n_2489)
);

NAND2x1p5_ASAP7_75t_L g2490 ( 
.A(n_2333),
.B(n_2307),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2363),
.B(n_2223),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2359),
.Y(n_2492)
);

AO221x2_ASAP7_75t_L g2493 ( 
.A1(n_2341),
.A2(n_2246),
.B1(n_2249),
.B2(n_2241),
.C(n_2237),
.Y(n_2493)
);

BUFx6f_ASAP7_75t_L g2494 ( 
.A(n_2336),
.Y(n_2494)
);

AOI22xp33_ASAP7_75t_L g2495 ( 
.A1(n_2342),
.A2(n_2227),
.B1(n_2305),
.B2(n_2299),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2325),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2330),
.Y(n_2497)
);

INVx3_ASAP7_75t_SL g2498 ( 
.A(n_2428),
.Y(n_2498)
);

AND2x2_ASAP7_75t_L g2499 ( 
.A(n_2398),
.B(n_2227),
.Y(n_2499)
);

AOI21xp33_ASAP7_75t_L g2500 ( 
.A1(n_2327),
.A2(n_2140),
.B(n_2134),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2379),
.B(n_2229),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2361),
.Y(n_2502)
);

OAI33xp33_ASAP7_75t_L g2503 ( 
.A1(n_2367),
.A2(n_2257),
.A3(n_2241),
.B1(n_1957),
.B2(n_1961),
.B3(n_1968),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2432),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2432),
.Y(n_2505)
);

INVx3_ASAP7_75t_L g2506 ( 
.A(n_2336),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2328),
.B(n_2295),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2383),
.B(n_2295),
.Y(n_2508)
);

NOR3xp33_ASAP7_75t_L g2509 ( 
.A(n_2408),
.B(n_2240),
.C(n_2238),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2389),
.B(n_2278),
.Y(n_2510)
);

OR2x2_ASAP7_75t_L g2511 ( 
.A(n_2412),
.B(n_2257),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2368),
.Y(n_2512)
);

OAI31xp33_ASAP7_75t_L g2513 ( 
.A1(n_2431),
.A2(n_2242),
.A3(n_2307),
.B(n_2131),
.Y(n_2513)
);

OAI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2394),
.A2(n_2307),
.B1(n_2278),
.B2(n_2242),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_2354),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2374),
.B(n_2240),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2375),
.B(n_2240),
.Y(n_2517)
);

AOI221xp5_ASAP7_75t_L g2518 ( 
.A1(n_2394),
.A2(n_2133),
.B1(n_2145),
.B2(n_2182),
.C(n_2180),
.Y(n_2518)
);

AOI22xp33_ASAP7_75t_SL g2519 ( 
.A1(n_2333),
.A2(n_2013),
.B1(n_1936),
.B2(n_1911),
.Y(n_2519)
);

NAND4xp25_ASAP7_75t_L g2520 ( 
.A(n_2362),
.B(n_2194),
.C(n_2188),
.D(n_2197),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2376),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2330),
.Y(n_2522)
);

OR2x2_ASAP7_75t_L g2523 ( 
.A(n_2343),
.B(n_2187),
.Y(n_2523)
);

OR2x2_ASAP7_75t_L g2524 ( 
.A(n_2390),
.B(n_2187),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2460),
.Y(n_2525)
);

INVx1_ASAP7_75t_SL g2526 ( 
.A(n_2498),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2445),
.B(n_2447),
.Y(n_2527)
);

OR2x6_ASAP7_75t_L g2528 ( 
.A(n_2463),
.B(n_2333),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2465),
.B(n_2416),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2467),
.B(n_2423),
.Y(n_2530)
);

AND2x2_ASAP7_75t_L g2531 ( 
.A(n_2467),
.B(n_2454),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2474),
.B(n_2385),
.Y(n_2532)
);

AND2x4_ASAP7_75t_L g2533 ( 
.A(n_2467),
.B(n_2351),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2504),
.Y(n_2534)
);

NOR3xp33_ASAP7_75t_L g2535 ( 
.A(n_2444),
.B(n_2365),
.C(n_2351),
.Y(n_2535)
);

AND2x2_ASAP7_75t_L g2536 ( 
.A(n_2474),
.B(n_2385),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2505),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2437),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2442),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2457),
.B(n_2397),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2457),
.B(n_2397),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2442),
.Y(n_2542)
);

INVxp67_ASAP7_75t_L g2543 ( 
.A(n_2442),
.Y(n_2543)
);

AOI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2450),
.A2(n_2407),
.B1(n_2365),
.B2(n_2392),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2455),
.B(n_2421),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2494),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2438),
.B(n_2491),
.Y(n_2547)
);

INVx1_ASAP7_75t_SL g2548 ( 
.A(n_2464),
.Y(n_2548)
);

INVx6_ASAP7_75t_L g2549 ( 
.A(n_2494),
.Y(n_2549)
);

AND2x2_ASAP7_75t_L g2550 ( 
.A(n_2489),
.B(n_2410),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2494),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_2441),
.B(n_2396),
.Y(n_2552)
);

INVx1_ASAP7_75t_SL g2553 ( 
.A(n_2464),
.Y(n_2553)
);

OAI31xp33_ASAP7_75t_L g2554 ( 
.A1(n_2443),
.A2(n_2418),
.A3(n_2381),
.B(n_2402),
.Y(n_2554)
);

OR2x2_ASAP7_75t_L g2555 ( 
.A(n_2441),
.B(n_2399),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2506),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2451),
.B(n_2410),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2452),
.B(n_2395),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2446),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2456),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2447),
.B(n_2405),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2478),
.B(n_2433),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2458),
.Y(n_2563)
);

OR2x2_ASAP7_75t_L g2564 ( 
.A(n_2462),
.B(n_2434),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2475),
.B(n_2404),
.Y(n_2565)
);

INVx4_ASAP7_75t_L g2566 ( 
.A(n_2473),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2468),
.B(n_2403),
.Y(n_2567)
);

AND2x4_ASAP7_75t_L g2568 ( 
.A(n_2483),
.B(n_2422),
.Y(n_2568)
);

AND2x2_ASAP7_75t_L g2569 ( 
.A(n_2470),
.B(n_2427),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2480),
.B(n_2406),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2506),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2461),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2499),
.B(n_2413),
.Y(n_2573)
);

OAI221xp5_ASAP7_75t_L g2574 ( 
.A1(n_2485),
.A2(n_2436),
.B1(n_2387),
.B2(n_2393),
.C(n_2419),
.Y(n_2574)
);

AND4x1_ASAP7_75t_L g2575 ( 
.A(n_2485),
.B(n_2197),
.C(n_29),
.D(n_26),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2510),
.B(n_2410),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_SL g2577 ( 
.A(n_2513),
.B(n_2440),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2453),
.B(n_2414),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2466),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2473),
.B(n_2335),
.Y(n_2580)
);

NOR2xp67_ASAP7_75t_SL g2581 ( 
.A(n_2481),
.B(n_2335),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2476),
.Y(n_2582)
);

INVxp67_ASAP7_75t_L g2583 ( 
.A(n_2469),
.Y(n_2583)
);

OR2x2_ASAP7_75t_L g2584 ( 
.A(n_2507),
.B(n_2414),
.Y(n_2584)
);

INVx2_ASAP7_75t_SL g2585 ( 
.A(n_2490),
.Y(n_2585)
);

INVxp67_ASAP7_75t_L g2586 ( 
.A(n_2448),
.Y(n_2586)
);

OR2x2_ASAP7_75t_L g2587 ( 
.A(n_2448),
.B(n_2419),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2477),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2490),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2508),
.B(n_2430),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2515),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2488),
.Y(n_2592)
);

OR2x2_ASAP7_75t_L g2593 ( 
.A(n_2482),
.B(n_2430),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2492),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2481),
.A2(n_2338),
.B1(n_2366),
.B2(n_2340),
.Y(n_2595)
);

OR2x2_ASAP7_75t_L g2596 ( 
.A(n_2482),
.B(n_2435),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2509),
.B(n_2435),
.Y(n_2597)
);

NAND2xp33_ASAP7_75t_L g2598 ( 
.A(n_2486),
.B(n_2393),
.Y(n_2598)
);

OR2x2_ASAP7_75t_L g2599 ( 
.A(n_2449),
.B(n_2338),
.Y(n_2599)
);

NAND5xp2_ASAP7_75t_L g2600 ( 
.A(n_2459),
.B(n_2366),
.C(n_2340),
.D(n_2409),
.E(n_30),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2515),
.B(n_2354),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2502),
.Y(n_2602)
);

NOR2x1p5_ASAP7_75t_L g2603 ( 
.A(n_2449),
.B(n_2354),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2439),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2486),
.B(n_2384),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_2513),
.B(n_2384),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2532),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2526),
.B(n_2495),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2532),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2531),
.B(n_2459),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2536),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2536),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2543),
.B(n_2472),
.Y(n_2613)
);

INVxp67_ASAP7_75t_L g2614 ( 
.A(n_2581),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2525),
.Y(n_2615)
);

OR2x2_ASAP7_75t_L g2616 ( 
.A(n_2599),
.B(n_2587),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2533),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2543),
.B(n_2512),
.Y(n_2618)
);

OR2x2_ASAP7_75t_L g2619 ( 
.A(n_2552),
.B(n_2484),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2555),
.B(n_2586),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2530),
.B(n_2493),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2548),
.B(n_2493),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2553),
.B(n_2439),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2539),
.B(n_2521),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2533),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2539),
.B(n_2542),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2547),
.B(n_2501),
.Y(n_2627)
);

OR2x2_ASAP7_75t_L g2628 ( 
.A(n_2586),
.B(n_2496),
.Y(n_2628)
);

AND2x2_ASAP7_75t_L g2629 ( 
.A(n_2547),
.B(n_2479),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2533),
.Y(n_2630)
);

INVx1_ASAP7_75t_SL g2631 ( 
.A(n_2549),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2538),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2559),
.Y(n_2633)
);

AND2x2_ASAP7_75t_L g2634 ( 
.A(n_2550),
.B(n_2497),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2534),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2542),
.B(n_2517),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2583),
.B(n_2487),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2537),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2560),
.Y(n_2639)
);

INVx1_ASAP7_75t_SL g2640 ( 
.A(n_2549),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2550),
.B(n_2522),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2541),
.B(n_2516),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2541),
.B(n_2516),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2544),
.A2(n_2577),
.B1(n_2527),
.B2(n_2561),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2540),
.B(n_2514),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2557),
.B(n_2514),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2549),
.Y(n_2647)
);

OR2x6_ASAP7_75t_L g2648 ( 
.A(n_2583),
.B(n_2511),
.Y(n_2648)
);

AND2x2_ASAP7_75t_L g2649 ( 
.A(n_2557),
.B(n_2384),
.Y(n_2649)
);

AND2x4_ASAP7_75t_L g2650 ( 
.A(n_2566),
.B(n_2409),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2546),
.B(n_2409),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2535),
.B(n_2500),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2566),
.B(n_2524),
.Y(n_2653)
);

INVx1_ASAP7_75t_SL g2654 ( 
.A(n_2598),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2546),
.B(n_2551),
.Y(n_2655)
);

NAND2x1p5_ASAP7_75t_L g2656 ( 
.A(n_2575),
.B(n_2013),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_2535),
.B(n_2500),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2528),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2551),
.B(n_2523),
.Y(n_2659)
);

NOR2x1_ASAP7_75t_L g2660 ( 
.A(n_2598),
.B(n_2520),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2563),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2562),
.B(n_2585),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2577),
.B(n_2544),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2585),
.B(n_2519),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2572),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2528),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2566),
.B(n_28),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2528),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2644),
.A2(n_2574),
.B1(n_2606),
.B2(n_2605),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2607),
.Y(n_2670)
);

NAND2xp5_ASAP7_75t_L g2671 ( 
.A(n_2654),
.B(n_2554),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2609),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2663),
.B(n_2579),
.Y(n_2673)
);

AND2x4_ASAP7_75t_L g2674 ( 
.A(n_2617),
.B(n_2568),
.Y(n_2674)
);

INVx1_ASAP7_75t_SL g2675 ( 
.A(n_2631),
.Y(n_2675)
);

OAI22xp33_ASAP7_75t_SL g2676 ( 
.A1(n_2660),
.A2(n_2657),
.B1(n_2614),
.B2(n_2652),
.Y(n_2676)
);

OAI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2656),
.A2(n_2606),
.B1(n_2589),
.B2(n_2605),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2617),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2627),
.B(n_2569),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2650),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2611),
.Y(n_2681)
);

AOI22xp5_ASAP7_75t_L g2682 ( 
.A1(n_2637),
.A2(n_2567),
.B1(n_2589),
.B2(n_2603),
.Y(n_2682)
);

AOI21xp5_ASAP7_75t_L g2683 ( 
.A1(n_2613),
.A2(n_2600),
.B(n_2595),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2640),
.B(n_2556),
.Y(n_2684)
);

A2O1A1Ixp33_ASAP7_75t_L g2685 ( 
.A1(n_2610),
.A2(n_2595),
.B(n_2471),
.C(n_2597),
.Y(n_2685)
);

INVx2_ASAP7_75t_SL g2686 ( 
.A(n_2650),
.Y(n_2686)
);

OR2x2_ASAP7_75t_L g2687 ( 
.A(n_2612),
.B(n_2564),
.Y(n_2687)
);

AOI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2610),
.A2(n_2592),
.B1(n_2594),
.B2(n_2588),
.C(n_2582),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2650),
.Y(n_2689)
);

INVx1_ASAP7_75t_SL g2690 ( 
.A(n_2667),
.Y(n_2690)
);

NOR2x1p5_ASAP7_75t_L g2691 ( 
.A(n_2626),
.B(n_2647),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2655),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2655),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2630),
.B(n_2602),
.Y(n_2694)
);

AND2x2_ASAP7_75t_L g2695 ( 
.A(n_2627),
.B(n_2576),
.Y(n_2695)
);

AOI32xp33_ASAP7_75t_L g2696 ( 
.A1(n_2629),
.A2(n_2568),
.A3(n_2604),
.B1(n_2571),
.B2(n_2556),
.Y(n_2696)
);

INVx2_ASAP7_75t_L g2697 ( 
.A(n_2630),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2628),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2628),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2619),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2619),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2615),
.B(n_2545),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2618),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2625),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2648),
.B(n_2584),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2616),
.Y(n_2706)
);

NOR2xp33_ASAP7_75t_L g2707 ( 
.A(n_2608),
.B(n_2578),
.Y(n_2707)
);

AO21x1_ASAP7_75t_L g2708 ( 
.A1(n_2667),
.A2(n_2568),
.B(n_2571),
.Y(n_2708)
);

AOI221xp5_ASAP7_75t_L g2709 ( 
.A1(n_2622),
.A2(n_2591),
.B1(n_2545),
.B2(n_2503),
.C(n_2604),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2647),
.B(n_2545),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2616),
.Y(n_2711)
);

O2A1O1Ixp33_ASAP7_75t_L g2712 ( 
.A1(n_2648),
.A2(n_2471),
.B(n_2591),
.C(n_2593),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2662),
.B(n_2576),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2662),
.B(n_2573),
.Y(n_2714)
);

INVx2_ASAP7_75t_L g2715 ( 
.A(n_2658),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2678),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_SL g2717 ( 
.A(n_2676),
.B(n_2656),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2674),
.Y(n_2718)
);

OAI21xp5_ASAP7_75t_SL g2719 ( 
.A1(n_2669),
.A2(n_2608),
.B(n_2656),
.Y(n_2719)
);

AND2x4_ASAP7_75t_L g2720 ( 
.A(n_2674),
.B(n_2658),
.Y(n_2720)
);

AOI21xp33_ASAP7_75t_L g2721 ( 
.A1(n_2676),
.A2(n_2648),
.B(n_2620),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2692),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2685),
.A2(n_2648),
.B1(n_2620),
.B2(n_2622),
.Y(n_2723)
);

AOI22xp33_ASAP7_75t_L g2724 ( 
.A1(n_2683),
.A2(n_2629),
.B1(n_2646),
.B2(n_2645),
.Y(n_2724)
);

OAI221xp5_ASAP7_75t_L g2725 ( 
.A1(n_2682),
.A2(n_2666),
.B1(n_2668),
.B2(n_2636),
.C(n_2621),
.Y(n_2725)
);

OAI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2671),
.A2(n_2677),
.B1(n_2712),
.B2(n_2675),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2675),
.A2(n_2646),
.B1(n_2621),
.B2(n_2666),
.Y(n_2727)
);

O2A1O1Ixp33_ASAP7_75t_L g2728 ( 
.A1(n_2708),
.A2(n_2668),
.B(n_2633),
.C(n_2635),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2693),
.Y(n_2729)
);

NOR2xp33_ASAP7_75t_L g2730 ( 
.A(n_2707),
.B(n_2624),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2697),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2686),
.Y(n_2732)
);

AOI221xp5_ASAP7_75t_L g2733 ( 
.A1(n_2688),
.A2(n_2696),
.B1(n_2673),
.B2(n_2709),
.C(n_2706),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2690),
.B(n_2667),
.Y(n_2734)
);

INVx2_ASAP7_75t_SL g2735 ( 
.A(n_2689),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2673),
.A2(n_2623),
.B(n_2632),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2704),
.Y(n_2737)
);

OR2x2_ASAP7_75t_L g2738 ( 
.A(n_2690),
.B(n_2642),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2715),
.B(n_2632),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2711),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2713),
.B(n_2623),
.Y(n_2741)
);

OAI22xp5_ASAP7_75t_L g2742 ( 
.A1(n_2705),
.A2(n_2645),
.B1(n_2633),
.B2(n_2638),
.Y(n_2742)
);

AOI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2695),
.A2(n_2649),
.B1(n_2641),
.B2(n_2634),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2679),
.B(n_2634),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2680),
.B(n_2642),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2691),
.B(n_2641),
.Y(n_2746)
);

A2O1A1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2700),
.A2(n_2664),
.B(n_2635),
.C(n_2638),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2698),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2687),
.Y(n_2749)
);

AND2x2_ASAP7_75t_L g2750 ( 
.A(n_2714),
.B(n_2643),
.Y(n_2750)
);

AOI22xp33_ASAP7_75t_L g2751 ( 
.A1(n_2703),
.A2(n_2701),
.B1(n_2664),
.B2(n_2649),
.Y(n_2751)
);

A2O1A1Ixp33_ASAP7_75t_L g2752 ( 
.A1(n_2699),
.A2(n_2643),
.B(n_2661),
.C(n_2639),
.Y(n_2752)
);

OAI21xp33_ASAP7_75t_L g2753 ( 
.A1(n_2684),
.A2(n_2651),
.B(n_2659),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2720),
.B(n_2670),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2720),
.B(n_2672),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2741),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_2718),
.Y(n_2757)
);

AOI221xp5_ASAP7_75t_L g2758 ( 
.A1(n_2723),
.A2(n_2726),
.B1(n_2721),
.B2(n_2733),
.C(n_2717),
.Y(n_2758)
);

NAND3xp33_ASAP7_75t_L g2759 ( 
.A(n_2721),
.B(n_2694),
.C(n_2681),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2744),
.B(n_2710),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2734),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2726),
.A2(n_2651),
.B1(n_2659),
.B2(n_2653),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2735),
.B(n_2724),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2746),
.B(n_2702),
.Y(n_2764)
);

INVx2_ASAP7_75t_SL g2765 ( 
.A(n_2738),
.Y(n_2765)
);

INVx3_ASAP7_75t_L g2766 ( 
.A(n_2732),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2745),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2739),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2739),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2749),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2740),
.Y(n_2771)
);

OAI31xp33_ASAP7_75t_L g2772 ( 
.A1(n_2723),
.A2(n_2702),
.A3(n_2694),
.B(n_2665),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2728),
.A2(n_2653),
.B(n_2580),
.Y(n_2773)
);

AOI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2719),
.A2(n_2653),
.B1(n_2601),
.B2(n_2570),
.Y(n_2774)
);

OAI211xp5_ASAP7_75t_L g2775 ( 
.A1(n_2725),
.A2(n_2596),
.B(n_2520),
.C(n_2518),
.Y(n_2775)
);

AOI221xp5_ASAP7_75t_L g2776 ( 
.A1(n_2727),
.A2(n_2580),
.B1(n_2601),
.B2(n_2590),
.C(n_2565),
.Y(n_2776)
);

OR2x2_ASAP7_75t_L g2777 ( 
.A(n_2727),
.B(n_2558),
.Y(n_2777)
);

INVx2_ASAP7_75t_SL g2778 ( 
.A(n_2748),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2742),
.Y(n_2779)
);

A2O1A1Ixp33_ASAP7_75t_L g2780 ( 
.A1(n_2736),
.A2(n_2730),
.B(n_2747),
.C(n_2753),
.Y(n_2780)
);

INVx1_ASAP7_75t_SL g2781 ( 
.A(n_2750),
.Y(n_2781)
);

OAI21xp5_ASAP7_75t_L g2782 ( 
.A1(n_2743),
.A2(n_2580),
.B(n_2601),
.Y(n_2782)
);

OAI221xp5_ASAP7_75t_L g2783 ( 
.A1(n_2751),
.A2(n_2529),
.B1(n_1982),
.B2(n_1936),
.C(n_1911),
.Y(n_2783)
);

INVx1_ASAP7_75t_SL g2784 ( 
.A(n_2742),
.Y(n_2784)
);

A2O1A1Ixp33_ASAP7_75t_L g2785 ( 
.A1(n_2752),
.A2(n_2001),
.B(n_2117),
.C(n_1936),
.Y(n_2785)
);

AOI21xp33_ASAP7_75t_L g2786 ( 
.A1(n_2772),
.A2(n_2731),
.B(n_2716),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2754),
.Y(n_2787)
);

AOI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2758),
.A2(n_2729),
.B1(n_2722),
.B2(n_2737),
.Y(n_2788)
);

NOR3xp33_ASAP7_75t_L g2789 ( 
.A(n_2780),
.B(n_29),
.C(n_30),
.Y(n_2789)
);

OAI21xp5_ASAP7_75t_SL g2790 ( 
.A1(n_2772),
.A2(n_31),
.B(n_33),
.Y(n_2790)
);

OAI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2759),
.A2(n_2030),
.B(n_1996),
.Y(n_2791)
);

AOI22xp5_ASAP7_75t_L g2792 ( 
.A1(n_2775),
.A2(n_1936),
.B1(n_1961),
.B2(n_1957),
.Y(n_2792)
);

OAI211xp5_ASAP7_75t_L g2793 ( 
.A1(n_2784),
.A2(n_37),
.B(n_33),
.C(n_35),
.Y(n_2793)
);

NOR2xp33_ASAP7_75t_L g2794 ( 
.A(n_2781),
.B(n_37),
.Y(n_2794)
);

AOI211xp5_ASAP7_75t_L g2795 ( 
.A1(n_2759),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_2795)
);

AOI221xp5_ASAP7_75t_SL g2796 ( 
.A1(n_2773),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.C(n_42),
.Y(n_2796)
);

OAI211xp5_ASAP7_75t_SL g2797 ( 
.A1(n_2763),
.A2(n_44),
.B(n_41),
.C(n_43),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_SL g2798 ( 
.A1(n_2765),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_2798)
);

AOI211xp5_ASAP7_75t_L g2799 ( 
.A1(n_2782),
.A2(n_48),
.B(n_46),
.C(n_47),
.Y(n_2799)
);

NAND3xp33_ASAP7_75t_L g2800 ( 
.A(n_2762),
.B(n_49),
.C(n_50),
.Y(n_2800)
);

NAND4xp25_ASAP7_75t_L g2801 ( 
.A(n_2774),
.B(n_54),
.C(n_51),
.D(n_52),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2755),
.Y(n_2802)
);

OAI31xp33_ASAP7_75t_L g2803 ( 
.A1(n_2779),
.A2(n_55),
.A3(n_51),
.B(n_54),
.Y(n_2803)
);

OAI22xp33_ASAP7_75t_SL g2804 ( 
.A1(n_2777),
.A2(n_1961),
.B1(n_1968),
.B2(n_1957),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2756),
.B(n_2766),
.Y(n_2805)
);

AOI221xp5_ASAP7_75t_L g2806 ( 
.A1(n_2776),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_60),
.Y(n_2806)
);

OAI21xp5_ASAP7_75t_SL g2807 ( 
.A1(n_2760),
.A2(n_57),
.B(n_58),
.Y(n_2807)
);

NOR3xp33_ASAP7_75t_L g2808 ( 
.A(n_2764),
.B(n_60),
.C(n_63),
.Y(n_2808)
);

INVxp33_ASAP7_75t_SL g2809 ( 
.A(n_2770),
.Y(n_2809)
);

AOI211xp5_ASAP7_75t_L g2810 ( 
.A1(n_2761),
.A2(n_68),
.B(n_63),
.C(n_66),
.Y(n_2810)
);

AOI222xp33_ASAP7_75t_L g2811 ( 
.A1(n_2790),
.A2(n_2769),
.B1(n_2768),
.B2(n_2771),
.C1(n_2767),
.C2(n_2778),
.Y(n_2811)
);

AOI21xp33_ASAP7_75t_L g2812 ( 
.A1(n_2805),
.A2(n_2757),
.B(n_2766),
.Y(n_2812)
);

NOR4xp25_ASAP7_75t_L g2813 ( 
.A(n_2786),
.B(n_2783),
.C(n_2785),
.D(n_75),
.Y(n_2813)
);

O2A1O1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2797),
.A2(n_75),
.B(n_71),
.C(n_73),
.Y(n_2814)
);

AOI321xp33_ASAP7_75t_L g2815 ( 
.A1(n_2789),
.A2(n_2787),
.A3(n_2802),
.B1(n_2788),
.B2(n_2799),
.C(n_2806),
.Y(n_2815)
);

AOI22x1_ASAP7_75t_L g2816 ( 
.A1(n_2796),
.A2(n_78),
.B1(n_73),
.B2(n_76),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2798),
.Y(n_2817)
);

AOI21xp5_ASAP7_75t_L g2818 ( 
.A1(n_2809),
.A2(n_79),
.B(n_80),
.Y(n_2818)
);

OAI321xp33_ASAP7_75t_L g2819 ( 
.A1(n_2801),
.A2(n_81),
.A3(n_82),
.B1(n_85),
.B2(n_86),
.C(n_87),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2794),
.Y(n_2820)
);

AOI221xp5_ASAP7_75t_L g2821 ( 
.A1(n_2800),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.C(n_90),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2793),
.Y(n_2822)
);

AOI221xp5_ASAP7_75t_L g2823 ( 
.A1(n_2795),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.C(n_95),
.Y(n_2823)
);

O2A1O1Ixp33_ASAP7_75t_L g2824 ( 
.A1(n_2808),
.A2(n_96),
.B(n_92),
.C(n_94),
.Y(n_2824)
);

OAI211xp5_ASAP7_75t_L g2825 ( 
.A1(n_2807),
.A2(n_98),
.B(n_96),
.C(n_97),
.Y(n_2825)
);

OAI22xp5_ASAP7_75t_L g2826 ( 
.A1(n_2810),
.A2(n_1969),
.B1(n_1968),
.B2(n_1948),
.Y(n_2826)
);

O2A1O1Ixp33_ASAP7_75t_L g2827 ( 
.A1(n_2803),
.A2(n_102),
.B(n_97),
.C(n_99),
.Y(n_2827)
);

OAI211xp5_ASAP7_75t_L g2828 ( 
.A1(n_2792),
.A2(n_104),
.B(n_99),
.C(n_103),
.Y(n_2828)
);

NAND2xp33_ASAP7_75t_L g2829 ( 
.A(n_2791),
.B(n_103),
.Y(n_2829)
);

AOI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2817),
.A2(n_2804),
.B1(n_1969),
.B2(n_1943),
.Y(n_2830)
);

INVx3_ASAP7_75t_L g2831 ( 
.A(n_2820),
.Y(n_2831)
);

AOI22xp5_ASAP7_75t_L g2832 ( 
.A1(n_2822),
.A2(n_1969),
.B1(n_1943),
.B2(n_1948),
.Y(n_2832)
);

AOI221xp5_ASAP7_75t_L g2833 ( 
.A1(n_2813),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.C(n_108),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2816),
.Y(n_2834)
);

OAI21xp33_ASAP7_75t_SL g2835 ( 
.A1(n_2812),
.A2(n_1948),
.B(n_1943),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_L g2836 ( 
.A(n_2827),
.B(n_106),
.C(n_108),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2825),
.Y(n_2837)
);

OAI211xp5_ASAP7_75t_SL g2838 ( 
.A1(n_2811),
.A2(n_112),
.B(n_109),
.C(n_111),
.Y(n_2838)
);

OR2x2_ASAP7_75t_L g2839 ( 
.A(n_2828),
.B(n_111),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2824),
.Y(n_2840)
);

O2A1O1Ixp33_ASAP7_75t_L g2841 ( 
.A1(n_2814),
.A2(n_117),
.B(n_113),
.C(n_114),
.Y(n_2841)
);

AOI21xp5_ASAP7_75t_L g2842 ( 
.A1(n_2829),
.A2(n_2818),
.B(n_2819),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2839),
.Y(n_2843)
);

XNOR2xp5_ASAP7_75t_L g2844 ( 
.A(n_2834),
.B(n_2837),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2831),
.Y(n_2845)
);

AOI22xp33_ASAP7_75t_L g2846 ( 
.A1(n_2838),
.A2(n_2826),
.B1(n_2823),
.B2(n_2821),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2836),
.B(n_2815),
.Y(n_2847)
);

INVx2_ASAP7_75t_L g2848 ( 
.A(n_2840),
.Y(n_2848)
);

AOI322xp5_ASAP7_75t_L g2849 ( 
.A1(n_2833),
.A2(n_113),
.A3(n_118),
.B1(n_119),
.B2(n_121),
.C1(n_122),
.C2(n_123),
.Y(n_2849)
);

OAI211xp5_ASAP7_75t_L g2850 ( 
.A1(n_2842),
.A2(n_124),
.B(n_118),
.C(n_122),
.Y(n_2850)
);

O2A1O1Ixp33_ASAP7_75t_L g2851 ( 
.A1(n_2841),
.A2(n_126),
.B(n_124),
.C(n_125),
.Y(n_2851)
);

A2O1A1Ixp33_ASAP7_75t_L g2852 ( 
.A1(n_2835),
.A2(n_130),
.B(n_126),
.C(n_129),
.Y(n_2852)
);

AOI21xp5_ASAP7_75t_L g2853 ( 
.A1(n_2830),
.A2(n_129),
.B(n_131),
.Y(n_2853)
);

OAI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2832),
.A2(n_132),
.B(n_133),
.Y(n_2854)
);

AOI221xp5_ASAP7_75t_L g2855 ( 
.A1(n_2838),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.C(n_140),
.Y(n_2855)
);

BUFx2_ASAP7_75t_L g2856 ( 
.A(n_2845),
.Y(n_2856)
);

AND2x4_ASAP7_75t_L g2857 ( 
.A(n_2848),
.B(n_140),
.Y(n_2857)
);

AO22x2_ASAP7_75t_SL g2858 ( 
.A1(n_2843),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2844),
.Y(n_2859)
);

AND2x4_ASAP7_75t_L g2860 ( 
.A(n_2847),
.B(n_145),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2850),
.Y(n_2861)
);

NOR2x1_ASAP7_75t_L g2862 ( 
.A(n_2851),
.B(n_146),
.Y(n_2862)
);

INVxp67_ASAP7_75t_SL g2863 ( 
.A(n_2855),
.Y(n_2863)
);

NOR2x1_ASAP7_75t_L g2864 ( 
.A(n_2854),
.B(n_146),
.Y(n_2864)
);

AOI22xp5_ASAP7_75t_L g2865 ( 
.A1(n_2846),
.A2(n_2123),
.B1(n_2112),
.B2(n_1987),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2852),
.Y(n_2866)
);

INVx1_ASAP7_75t_SL g2867 ( 
.A(n_2853),
.Y(n_2867)
);

AO22x1_ASAP7_75t_L g2868 ( 
.A1(n_2849),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_2868)
);

AOI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2845),
.A2(n_2123),
.B1(n_2112),
.B2(n_1987),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2850),
.B(n_147),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2844),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2845),
.Y(n_2872)
);

OAI221xp5_ASAP7_75t_SL g2873 ( 
.A1(n_2861),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.C(n_151),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2858),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2871),
.A2(n_1987),
.B1(n_1998),
.B2(n_2040),
.Y(n_2875)
);

INVxp67_ASAP7_75t_L g2876 ( 
.A(n_2870),
.Y(n_2876)
);

HB1xp67_ASAP7_75t_L g2877 ( 
.A(n_2857),
.Y(n_2877)
);

NOR2x1_ASAP7_75t_L g2878 ( 
.A(n_2856),
.B(n_151),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2856),
.B(n_152),
.Y(n_2879)
);

XNOR2xp5_ASAP7_75t_L g2880 ( 
.A(n_2859),
.B(n_153),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2860),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2868),
.B(n_154),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2862),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2872),
.Y(n_2884)
);

AOI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2863),
.A2(n_154),
.B(n_155),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2866),
.B(n_155),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2867),
.B(n_156),
.Y(n_2887)
);

OAI221xp5_ASAP7_75t_R g2888 ( 
.A1(n_2880),
.A2(n_2865),
.B1(n_2869),
.B2(n_2864),
.C(n_160),
.Y(n_2888)
);

NAND4xp25_ASAP7_75t_L g2889 ( 
.A(n_2874),
.B(n_157),
.C(n_158),
.D(n_159),
.Y(n_2889)
);

OAI311xp33_ASAP7_75t_L g2890 ( 
.A1(n_2883),
.A2(n_157),
.A3(n_160),
.B1(n_161),
.C1(n_162),
.Y(n_2890)
);

AOI22xp5_ASAP7_75t_L g2891 ( 
.A1(n_2884),
.A2(n_1998),
.B1(n_2040),
.B2(n_2033),
.Y(n_2891)
);

O2A1O1Ixp5_ASAP7_75t_SL g2892 ( 
.A1(n_2876),
.A2(n_161),
.B(n_162),
.C(n_163),
.Y(n_2892)
);

OA22x2_ASAP7_75t_L g2893 ( 
.A1(n_2879),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_2893)
);

AOI222xp33_ASAP7_75t_L g2894 ( 
.A1(n_2881),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.C1(n_170),
.C2(n_171),
.Y(n_2894)
);

OA22x2_ASAP7_75t_L g2895 ( 
.A1(n_2882),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_2895)
);

NAND4xp25_ASAP7_75t_L g2896 ( 
.A(n_2887),
.B(n_172),
.C(n_173),
.D(n_174),
.Y(n_2896)
);

OR2x6_ASAP7_75t_L g2897 ( 
.A(n_2878),
.B(n_172),
.Y(n_2897)
);

NOR4xp25_ASAP7_75t_L g2898 ( 
.A(n_2886),
.B(n_173),
.C(n_175),
.D(n_177),
.Y(n_2898)
);

OAI211xp5_ASAP7_75t_SL g2899 ( 
.A1(n_2877),
.A2(n_2885),
.B(n_2875),
.C(n_2873),
.Y(n_2899)
);

OR2x2_ASAP7_75t_L g2900 ( 
.A(n_2898),
.B(n_175),
.Y(n_2900)
);

OAI22xp33_ASAP7_75t_L g2901 ( 
.A1(n_2897),
.A2(n_177),
.B1(n_178),
.B2(n_181),
.Y(n_2901)
);

INVx2_ASAP7_75t_L g2902 ( 
.A(n_2893),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2895),
.Y(n_2903)
);

NAND3xp33_ASAP7_75t_L g2904 ( 
.A(n_2892),
.B(n_178),
.C(n_181),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2894),
.B(n_182),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2889),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2896),
.B(n_182),
.Y(n_2907)
);

OAI21xp33_ASAP7_75t_L g2908 ( 
.A1(n_2899),
.A2(n_183),
.B(n_184),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2891),
.Y(n_2909)
);

XNOR2x1_ASAP7_75t_L g2910 ( 
.A(n_2890),
.B(n_187),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2902),
.B(n_2903),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2910),
.Y(n_2912)
);

XNOR2xp5_ASAP7_75t_L g2913 ( 
.A(n_2906),
.B(n_2888),
.Y(n_2913)
);

XNOR2x1_ASAP7_75t_L g2914 ( 
.A(n_2900),
.B(n_188),
.Y(n_2914)
);

INVx1_ASAP7_75t_SL g2915 ( 
.A(n_2905),
.Y(n_2915)
);

AND2x4_ASAP7_75t_L g2916 ( 
.A(n_2909),
.B(n_188),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2907),
.Y(n_2917)
);

OAI22xp5_ASAP7_75t_SL g2918 ( 
.A1(n_2904),
.A2(n_2908),
.B1(n_2901),
.B2(n_191),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2910),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2900),
.Y(n_2920)
);

XNOR2xp5_ASAP7_75t_L g2921 ( 
.A(n_2910),
.B(n_189),
.Y(n_2921)
);

INVx4_ASAP7_75t_L g2922 ( 
.A(n_2902),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2910),
.Y(n_2923)
);

INVx3_ASAP7_75t_L g2924 ( 
.A(n_2916),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2921),
.Y(n_2925)
);

AOI22xp5_ASAP7_75t_L g2926 ( 
.A1(n_2911),
.A2(n_189),
.B1(n_190),
.B2(n_192),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2921),
.Y(n_2927)
);

INVxp33_ASAP7_75t_L g2928 ( 
.A(n_2914),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2918),
.Y(n_2929)
);

INVx1_ASAP7_75t_SL g2930 ( 
.A(n_2915),
.Y(n_2930)
);

BUFx2_ASAP7_75t_L g2931 ( 
.A(n_2912),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2919),
.Y(n_2932)
);

OAI21x1_ASAP7_75t_SL g2933 ( 
.A1(n_2932),
.A2(n_2913),
.B(n_2920),
.Y(n_2933)
);

OA21x2_ASAP7_75t_L g2934 ( 
.A1(n_2931),
.A2(n_2923),
.B(n_2917),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2930),
.A2(n_2922),
.B1(n_193),
.B2(n_194),
.Y(n_2935)
);

OAI21xp5_ASAP7_75t_L g2936 ( 
.A1(n_2928),
.A2(n_192),
.B(n_194),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2924),
.B(n_195),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2925),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2926),
.B(n_196),
.Y(n_2939)
);

OAI21xp33_ASAP7_75t_L g2940 ( 
.A1(n_2927),
.A2(n_196),
.B(n_197),
.Y(n_2940)
);

HB1xp67_ASAP7_75t_L g2941 ( 
.A(n_2929),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2931),
.Y(n_2942)
);

HB1xp67_ASAP7_75t_L g2943 ( 
.A(n_2931),
.Y(n_2943)
);

OAI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2932),
.A2(n_198),
.B1(n_199),
.B2(n_200),
.Y(n_2944)
);

AO22x2_ASAP7_75t_L g2945 ( 
.A1(n_2932),
.A2(n_199),
.B1(n_201),
.B2(n_210),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2932),
.A2(n_864),
.B(n_863),
.Y(n_2946)
);

OA22x2_ASAP7_75t_L g2947 ( 
.A1(n_2932),
.A2(n_1998),
.B1(n_2040),
.B2(n_2033),
.Y(n_2947)
);

OAI22xp5_ASAP7_75t_L g2948 ( 
.A1(n_2932),
.A2(n_2033),
.B1(n_864),
.B2(n_2043),
.Y(n_2948)
);

INVx2_ASAP7_75t_SL g2949 ( 
.A(n_2931),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2931),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2931),
.B(n_217),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2931),
.Y(n_2952)
);

OAI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2949),
.A2(n_1464),
.B1(n_1442),
.B2(n_1435),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2937),
.Y(n_2954)
);

AOI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2942),
.A2(n_863),
.B1(n_874),
.B2(n_1322),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2935),
.B(n_220),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2943),
.Y(n_2957)
);

CKINVDCx20_ASAP7_75t_R g2958 ( 
.A(n_2941),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2950),
.Y(n_2959)
);

OAI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2952),
.A2(n_2951),
.B1(n_2938),
.B2(n_2939),
.Y(n_2960)
);

OAI22xp5_ASAP7_75t_SL g2961 ( 
.A1(n_2934),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_2961)
);

NAND4xp25_ASAP7_75t_L g2962 ( 
.A(n_2936),
.B(n_225),
.C(n_227),
.D(n_231),
.Y(n_2962)
);

AO22x2_ASAP7_75t_L g2963 ( 
.A1(n_2933),
.A2(n_2944),
.B1(n_2946),
.B2(n_2940),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2945),
.Y(n_2964)
);

AO22x2_ASAP7_75t_L g2965 ( 
.A1(n_2945),
.A2(n_233),
.B1(n_235),
.B2(n_237),
.Y(n_2965)
);

BUFx2_ASAP7_75t_L g2966 ( 
.A(n_2947),
.Y(n_2966)
);

AOI21xp5_ASAP7_75t_L g2967 ( 
.A1(n_2948),
.A2(n_917),
.B(n_893),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2937),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_L g2969 ( 
.A1(n_2949),
.A2(n_917),
.B1(n_863),
.B2(n_874),
.Y(n_2969)
);

OAI22xp5_ASAP7_75t_SL g2970 ( 
.A1(n_2942),
.A2(n_239),
.B1(n_242),
.B2(n_245),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2937),
.Y(n_2971)
);

INVx1_ASAP7_75t_L g2972 ( 
.A(n_2937),
.Y(n_2972)
);

CKINVDCx20_ASAP7_75t_R g2973 ( 
.A(n_2943),
.Y(n_2973)
);

INVxp67_ASAP7_75t_L g2974 ( 
.A(n_2937),
.Y(n_2974)
);

OAI22xp5_ASAP7_75t_L g2975 ( 
.A1(n_2949),
.A2(n_1299),
.B1(n_1302),
.B2(n_1298),
.Y(n_2975)
);

OAI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2949),
.A2(n_1305),
.B1(n_1306),
.B2(n_851),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_2957),
.B(n_917),
.Y(n_2977)
);

OAI21xp5_ASAP7_75t_SL g2978 ( 
.A1(n_2959),
.A2(n_247),
.B(n_250),
.Y(n_2978)
);

AOI221xp5_ASAP7_75t_L g2979 ( 
.A1(n_2964),
.A2(n_884),
.B1(n_888),
.B2(n_893),
.C(n_1324),
.Y(n_2979)
);

OAI22xp5_ASAP7_75t_L g2980 ( 
.A1(n_2973),
.A2(n_851),
.B1(n_1322),
.B2(n_1324),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2954),
.B(n_251),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2968),
.B(n_252),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2958),
.Y(n_2983)
);

OAI21x1_ASAP7_75t_L g2984 ( 
.A1(n_2956),
.A2(n_2030),
.B(n_1324),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_2971),
.A2(n_874),
.B1(n_863),
.B2(n_851),
.Y(n_2985)
);

AOI221xp5_ASAP7_75t_L g2986 ( 
.A1(n_2960),
.A2(n_2966),
.B1(n_2965),
.B2(n_2953),
.C(n_2963),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2974),
.A2(n_893),
.B(n_888),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2963),
.Y(n_2988)
);

OAI22xp5_ASAP7_75t_SL g2989 ( 
.A1(n_2961),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2972),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2970),
.Y(n_2991)
);

OAI22xp33_ASAP7_75t_L g2992 ( 
.A1(n_2962),
.A2(n_1464),
.B1(n_1442),
.B2(n_1322),
.Y(n_2992)
);

OAI21xp5_ASAP7_75t_L g2993 ( 
.A1(n_2967),
.A2(n_863),
.B(n_874),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2976),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2975),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2955),
.B(n_257),
.Y(n_2996)
);

OAI21xp5_ASAP7_75t_L g2997 ( 
.A1(n_2969),
.A2(n_874),
.B(n_884),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2957),
.B(n_260),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2957),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2998),
.Y(n_3000)
);

AOI222xp33_ASAP7_75t_L g3001 ( 
.A1(n_2999),
.A2(n_874),
.B1(n_264),
.B2(n_268),
.C1(n_269),
.C2(n_272),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_L g3002 ( 
.A1(n_2983),
.A2(n_851),
.B1(n_884),
.B2(n_888),
.Y(n_3002)
);

AOI21xp33_ASAP7_75t_L g3003 ( 
.A1(n_2988),
.A2(n_262),
.B(n_274),
.Y(n_3003)
);

OAI22xp33_ASAP7_75t_L g3004 ( 
.A1(n_2981),
.A2(n_1464),
.B1(n_1283),
.B2(n_280),
.Y(n_3004)
);

OAI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2982),
.A2(n_277),
.B1(n_278),
.B2(n_281),
.Y(n_3005)
);

OAI21xp5_ASAP7_75t_L g3006 ( 
.A1(n_2990),
.A2(n_282),
.B(n_287),
.Y(n_3006)
);

OAI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2991),
.A2(n_1312),
.B1(n_1304),
.B2(n_1293),
.Y(n_3007)
);

AOI21xp5_ASAP7_75t_L g3008 ( 
.A1(n_2986),
.A2(n_873),
.B(n_857),
.Y(n_3008)
);

AO21x2_ASAP7_75t_L g3009 ( 
.A1(n_2977),
.A2(n_2987),
.B(n_2997),
.Y(n_3009)
);

OAI21xp33_ASAP7_75t_SL g3010 ( 
.A1(n_2996),
.A2(n_292),
.B(n_294),
.Y(n_3010)
);

OAI22xp5_ASAP7_75t_L g3011 ( 
.A1(n_2989),
.A2(n_1312),
.B1(n_1304),
.B2(n_1293),
.Y(n_3011)
);

AOI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_3000),
.A2(n_2978),
.B1(n_2992),
.B2(n_2995),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_3010),
.A2(n_2994),
.B1(n_2980),
.B2(n_2979),
.Y(n_3013)
);

AOI222xp33_ASAP7_75t_L g3014 ( 
.A1(n_3007),
.A2(n_2993),
.B1(n_2984),
.B2(n_2985),
.C1(n_303),
.C2(n_306),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_L g3015 ( 
.A1(n_3004),
.A2(n_3009),
.B1(n_3008),
.B2(n_3001),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_3011),
.Y(n_3016)
);

AOI222xp33_ASAP7_75t_L g3017 ( 
.A1(n_3006),
.A2(n_296),
.B1(n_301),
.B2(n_302),
.C1(n_308),
.C2(n_311),
.Y(n_3017)
);

AOI22xp5_ASAP7_75t_L g3018 ( 
.A1(n_3005),
.A2(n_1288),
.B1(n_1284),
.B2(n_1229),
.Y(n_3018)
);

AOI21xp33_ASAP7_75t_SL g3019 ( 
.A1(n_3003),
.A2(n_313),
.B(n_316),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_3012),
.A2(n_3002),
.B1(n_1288),
.B2(n_1284),
.Y(n_3020)
);

AOI22xp5_ASAP7_75t_L g3021 ( 
.A1(n_3013),
.A2(n_3014),
.B1(n_3017),
.B2(n_3015),
.Y(n_3021)
);

AOI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_3016),
.A2(n_3018),
.B1(n_3019),
.B2(n_1229),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_3016),
.A2(n_880),
.B1(n_881),
.B2(n_883),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_3012),
.A2(n_1229),
.B1(n_1207),
.B2(n_1195),
.Y(n_3024)
);

AOI22xp5_ASAP7_75t_L g3025 ( 
.A1(n_3012),
.A2(n_1207),
.B1(n_1195),
.B2(n_883),
.Y(n_3025)
);

NAND2x1p5_ASAP7_75t_L g3026 ( 
.A(n_3021),
.B(n_873),
.Y(n_3026)
);

OA22x2_ASAP7_75t_L g3027 ( 
.A1(n_3022),
.A2(n_333),
.B1(n_337),
.B2(n_338),
.Y(n_3027)
);

AOI21xp5_ASAP7_75t_L g3028 ( 
.A1(n_3026),
.A2(n_3020),
.B(n_3025),
.Y(n_3028)
);

AOI211xp5_ASAP7_75t_L g3029 ( 
.A1(n_3028),
.A2(n_3024),
.B(n_3027),
.C(n_3023),
.Y(n_3029)
);


endmodule