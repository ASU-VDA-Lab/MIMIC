module fake_jpeg_116_n_360 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_7),
.B(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_12),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_56),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_24),
.Y(n_48)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_0),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_53),
.B(n_75),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_25),
.B(n_14),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_18),
.B(n_10),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_61),
.B(n_77),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_76),
.Y(n_100)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_89),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_22),
.B(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_85),
.B(n_117),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_22),
.B1(n_26),
.B2(n_32),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_86),
.A2(n_91),
.B1(n_121),
.B2(n_1),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_17),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_58),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_90),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_33),
.B1(n_32),
.B2(n_41),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_96),
.B(n_128),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_33),
.B1(n_32),
.B2(n_41),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_103),
.A2(n_110),
.B1(n_54),
.B2(n_44),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_52),
.A2(n_33),
.B1(n_17),
.B2(n_41),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_51),
.B(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_122),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_65),
.A2(n_33),
.B1(n_35),
.B2(n_27),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_30),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_70),
.A2(n_34),
.B1(n_35),
.B2(n_29),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_16),
.B1(n_27),
.B2(n_28),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_75),
.B(n_38),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_131),
.B1(n_154),
.B2(n_165),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_112),
.B1(n_110),
.B2(n_49),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_130),
.A2(n_113),
.B1(n_104),
.B2(n_7),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_115),
.B1(n_81),
.B2(n_105),
.Y(n_131)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_133),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_135),
.A2(n_140),
.B(n_155),
.Y(n_191)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_142),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_84),
.A2(n_76),
.B1(n_78),
.B2(n_108),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_161),
.B1(n_164),
.B2(n_124),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_106),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_147),
.A2(n_148),
.B(n_159),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_59),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_87),
.B(n_59),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_80),
.A2(n_71),
.B1(n_55),
.B2(n_54),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_44),
.B1(n_23),
.B2(n_2),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_157),
.B(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_93),
.B(n_0),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_82),
.B(n_1),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_105),
.A2(n_23),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_170),
.Y(n_175)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_98),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_166),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_92),
.B(n_11),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_169),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_97),
.A2(n_11),
.B1(n_10),
.B2(n_6),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_120),
.B1(n_109),
.B2(n_10),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_102),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_109),
.A2(n_1),
.B(n_4),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_4),
.B(n_6),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_99),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_172),
.B(n_184),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_98),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_99),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_165),
.A2(n_118),
.B1(n_80),
.B2(n_124),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_183),
.A2(n_190),
.B1(n_195),
.B2(n_203),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_134),
.B(n_101),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_99),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_186),
.B(n_174),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_147),
.B(n_130),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_192),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_158),
.B(n_118),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_196),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_120),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_147),
.A2(n_113),
.B1(n_104),
.B2(n_7),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_199),
.A2(n_205),
.B1(n_136),
.B2(n_152),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_171),
.B(n_170),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_154),
.B1(n_150),
.B2(n_159),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_7),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_153),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_187),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_226),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_210),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_192),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_217),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_220),
.Y(n_243)
);

OR2x2_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_198),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_219),
.B(n_222),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_139),
.C(n_157),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_139),
.B(n_169),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_237),
.B(n_195),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_151),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_184),
.B(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_227),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_160),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_148),
.C(n_166),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_231),
.B1(n_182),
.B2(n_173),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_185),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_175),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_239),
.Y(n_250)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_183),
.A2(n_133),
.B1(n_148),
.B2(n_166),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_204),
.A2(n_156),
.B(n_146),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_236),
.B(n_188),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_132),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_189),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_149),
.B(n_142),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_205),
.A2(n_138),
.B(n_133),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_SL g238 ( 
.A(n_199),
.B(n_8),
.C(n_9),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_191),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_173),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_182),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_252),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_SL g281 ( 
.A1(n_244),
.A2(n_253),
.B(n_260),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_225),
.B1(n_212),
.B2(n_236),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_247),
.A2(n_264),
.B(n_218),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_251),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_219),
.Y(n_252)
);

CKINVDCx12_ASAP7_75t_R g255 ( 
.A(n_226),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_188),
.B1(n_208),
.B2(n_202),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_230),
.B1(n_232),
.B2(n_194),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_265),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_262),
.B(n_266),
.Y(n_276)
);

OR2x4_ASAP7_75t_L g264 ( 
.A(n_216),
.B(n_211),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_209),
.B(n_206),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_212),
.B(n_208),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_213),
.C(n_216),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_269),
.C(n_272),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_211),
.B1(n_224),
.B2(n_221),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_255),
.B1(n_245),
.B2(n_242),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_217),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_273),
.B1(n_274),
.B2(n_279),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_217),
.C(n_223),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_246),
.A2(n_225),
.B1(n_220),
.B2(n_237),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_241),
.A2(n_231),
.B1(n_228),
.B2(n_233),
.Y(n_274)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_258),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_253),
.A2(n_210),
.B1(n_234),
.B2(n_235),
.Y(n_279)
);

OAI21xp33_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_258),
.B(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_223),
.B1(n_229),
.B2(n_214),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_282),
.A2(n_284),
.B1(n_286),
.B2(n_265),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_247),
.A2(n_229),
.B1(n_189),
.B2(n_238),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_251),
.A2(n_202),
.B1(n_200),
.B2(n_179),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_304),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_276),
.Y(n_292)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_293),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_297),
.B1(n_303),
.B2(n_268),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_259),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_302),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_245),
.B(n_250),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_296),
.A2(n_300),
.B(n_277),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_287),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_299),
.Y(n_320)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_271),
.B(n_250),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_278),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_269),
.B(n_243),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_243),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_262),
.C(n_248),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_297),
.B1(n_298),
.B2(n_270),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_306),
.B(n_310),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_272),
.C(n_267),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_307),
.B(n_311),
.C(n_304),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_308),
.A2(n_320),
.B(n_318),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_282),
.C(n_285),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_279),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_311),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_271),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_296),
.B1(n_294),
.B2(n_292),
.Y(n_317)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_330),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_305),
.B(n_299),
.C(n_281),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_308),
.B(n_306),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_326),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_331),
.C(n_330),
.Y(n_337)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_327),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_284),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_274),
.Y(n_331)
);

OAI21x1_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_326),
.B(n_323),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_324),
.B(n_307),
.C(n_309),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_337),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_315),
.B1(n_290),
.B2(n_316),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_340),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_327),
.A2(n_316),
.B(n_290),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_338),
.A2(n_286),
.B(n_275),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_314),
.C(n_273),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_336),
.Y(n_342)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_342),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_333),
.B(n_331),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_344),
.B(n_345),
.C(n_334),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_339),
.A2(n_328),
.B1(n_322),
.B2(n_340),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_346),
.A2(n_347),
.B(n_339),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_350),
.Y(n_352)
);

AOI322xp5_ASAP7_75t_L g351 ( 
.A1(n_341),
.A2(n_244),
.A3(n_334),
.B1(n_248),
.B2(n_263),
.C1(n_206),
.C2(n_174),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_351),
.B(n_341),
.C(n_263),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_353),
.B(n_179),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_343),
.B(n_349),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_355),
.Y(n_357)
);

AOI322xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_356),
.A3(n_352),
.B1(n_244),
.B2(n_200),
.C1(n_194),
.C2(n_201),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_358),
.A2(n_197),
.B(n_201),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_359),
.B(n_197),
.Y(n_360)
);


endmodule