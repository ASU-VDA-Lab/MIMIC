module real_jpeg_10254_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_3),
.A2(n_67),
.B1(n_73),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_90),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_90),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_90),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_SL g35 ( 
.A1(n_6),
.A2(n_36),
.B(n_38),
.C(n_39),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_6),
.B(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_7),
.Y(n_60)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_9),
.A2(n_67),
.B1(n_73),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_9),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_107),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_107),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_107),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_62),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_12),
.A2(n_67),
.B1(n_73),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_12),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_76),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_12),
.A2(n_36),
.B1(n_37),
.B2(n_76),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_76),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_15),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_15),
.A2(n_57),
.B(n_69),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_15),
.A2(n_67),
.B1(n_73),
.B2(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_15),
.B(n_133),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_15),
.A2(n_36),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_15),
.B(n_36),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_15),
.A2(n_26),
.B1(n_31),
.B2(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_15),
.A2(n_56),
.B(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_15),
.B(n_56),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_17),
.A2(n_67),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_17),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_17),
.A2(n_56),
.B1(n_57),
.B2(n_74),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_74),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_17),
.A2(n_36),
.B1(n_37),
.B2(n_74),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_118),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_94),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_21),
.B(n_94),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_46),
.B1(n_78),
.B2(n_79),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_23),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_45),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_26),
.A2(n_31),
.B1(n_49),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_26),
.A2(n_31),
.B1(n_83),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_26),
.A2(n_31),
.B1(n_169),
.B2(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_26),
.A2(n_31),
.B1(n_171),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_26),
.A2(n_31),
.B1(n_202),
.B2(n_218),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_27),
.A2(n_28),
.B1(n_115),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_27),
.A2(n_28),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_28),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_29),
.B(n_40),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_29),
.B(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_30),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_31),
.B(n_111),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_39),
.B1(n_41),
.B2(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_35),
.A2(n_39),
.B1(n_51),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_35),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_35),
.A2(n_39),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_35),
.A2(n_39),
.B1(n_177),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_35),
.A2(n_39),
.B1(n_200),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_35),
.A2(n_39),
.B1(n_136),
.B2(n_208),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_36),
.B(n_60),
.Y(n_215)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_37),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_38),
.Y(n_181)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_39),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_39),
.B(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_53),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_48),
.B(n_50),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_64),
.B1(n_65),
.B2(n_77),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_59),
.B1(n_61),
.B2(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_59),
.B1(n_93),
.B2(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_55),
.A2(n_59),
.B1(n_102),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_55),
.A2(n_59),
.B1(n_129),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_55),
.A2(n_59),
.B1(n_155),
.B2(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_56),
.A2(n_57),
.B1(n_68),
.B2(n_69),
.Y(n_71)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_58),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_59),
.B(n_111),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_71),
.B1(n_72),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_71),
.B1(n_89),
.B2(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_70),
.C(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_68),
.B(n_111),
.C(n_112),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_71),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.C(n_91),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_84),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_86),
.A2(n_135),
.B1(n_137),
.B2(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_99),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_103),
.C(n_108),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_108),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_160),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_142),
.B(n_159),
.Y(n_120)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_121),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_139),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_139),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.C(n_126),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_134),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_128),
.B1(n_134),
.B2(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_143),
.B(n_145),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_146),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_149),
.A2(n_151),
.B1(n_152),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_149),
.Y(n_238)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_153),
.A2(n_154),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_156),
.B(n_157),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_240),
.C(n_241),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_234),
.B(n_239),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_220),
.B(n_233),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_204),
.B(n_219),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_194),
.B(n_203),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_183),
.B(n_193),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_167),
.B(n_172),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_178),
.B2(n_182),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_173),
.B(n_182),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_176),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_178),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_188),
.B(n_192),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_196),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_199),
.C(n_201),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_205),
.B(n_206),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.CI(n_212),
.CON(n_206),
.SN(n_206)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_211),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_217),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_221),
.B(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_230),
.C(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_230),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_235),
.B(n_236),
.Y(n_239)
);


endmodule