module real_aes_18158_n_15 (n_13, n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_15);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_15;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_33;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_16;
wire n_37;
wire n_51;
wire n_35;
wire n_42;
wire n_45;
wire n_39;
wire n_27;
wire n_50;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_52;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_53;
wire n_36;
INVx2_ASAP7_75t_L g32 ( .A(n_0), .Y(n_32) );
AOI322xp5_ASAP7_75t_R g44 ( .A1(n_1), .A2(n_5), .A3(n_9), .B1(n_18), .B2(n_45), .C1(n_47), .C2(n_50), .Y(n_44) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_2), .B(n_8), .C(n_21), .Y(n_20) );
NOR5xp2_ASAP7_75t_SL g18 ( .A(n_3), .B(n_12), .C(n_19), .D(n_23), .E(n_24), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g37 ( .A(n_3), .Y(n_37) );
NAND2xp33_ASAP7_75t_R g26 ( .A(n_4), .B(n_7), .Y(n_26) );
NOR2xp33_ASAP7_75t_R g43 ( .A(n_4), .B(n_7), .Y(n_43) );
NOR2xp33_ASAP7_75t_R g45 ( .A(n_4), .B(n_46), .Y(n_45) );
CKINVDCx5p33_ASAP7_75t_R g53 ( .A(n_4), .Y(n_53) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_6), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g46 ( .A(n_7), .Y(n_46) );
NOR2xp33_ASAP7_75t_R g52 ( .A(n_7), .B(n_53), .Y(n_52) );
CKINVDCx5p33_ASAP7_75t_R g24 ( .A(n_10), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_11), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g42 ( .A(n_12), .Y(n_42) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_13), .Y(n_23) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_14), .Y(n_21) );
OAI221xp5_ASAP7_75t_R g15 ( .A1(n_16), .A2(n_17), .B1(n_27), .B2(n_33), .C(n_44), .Y(n_15) );
NAND2xp33_ASAP7_75t_R g17 ( .A(n_18), .B(n_25), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g49 ( .A(n_18), .Y(n_49) );
CKINVDCx5p33_ASAP7_75t_R g41 ( .A(n_19), .Y(n_41) );
NAND2xp33_ASAP7_75t_R g19 ( .A(n_20), .B(n_22), .Y(n_19) );
NAND2xp33_ASAP7_75t_R g38 ( .A(n_23), .B(n_39), .Y(n_38) );
NAND2xp33_ASAP7_75t_R g40 ( .A(n_24), .B(n_41), .Y(n_40) );
CKINVDCx16_ASAP7_75t_R g25 ( .A(n_26), .Y(n_25) );
INVx1_ASAP7_75t_SL g27 ( .A(n_28), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
BUFx2_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
NAND2xp33_ASAP7_75t_R g33 ( .A(n_34), .B(n_43), .Y(n_33) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_35), .Y(n_34) );
NAND2xp33_ASAP7_75t_R g35 ( .A(n_36), .B(n_42), .Y(n_35) );
NOR2xp33_ASAP7_75t_R g36 ( .A(n_37), .B(n_38), .Y(n_36) );
CKINVDCx5p33_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
CKINVDCx5p33_ASAP7_75t_R g48 ( .A(n_43), .Y(n_48) );
NOR2xp33_ASAP7_75t_R g47 ( .A(n_48), .B(n_49), .Y(n_47) );
NOR2xp33_ASAP7_75t_R g50 ( .A(n_49), .B(n_51), .Y(n_50) );
CKINVDCx5p33_ASAP7_75t_R g51 ( .A(n_52), .Y(n_51) );
endmodule