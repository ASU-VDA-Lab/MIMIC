module real_jpeg_5012_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_1),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_2),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_2),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_2),
.B(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_2),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_2),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_2),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_3),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_3),
.B(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_3),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_4),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_4),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_4),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_4),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_4),
.B(n_35),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_4),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_4),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_4),
.B(n_486),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_5),
.B(n_161),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_5),
.A2(n_65),
.B(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_5),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_5),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_5),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_5),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_5),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_5),
.B(n_388),
.Y(n_415)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_7),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_7),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_7),
.B(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_7),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_7),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_7),
.B(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_8),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_8),
.Y(n_325)
);

BUFx5_ASAP7_75t_L g388 ( 
.A(n_8),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_9),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_9),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_9),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_9),
.B(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_9),
.B(n_377),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_9),
.B(n_412),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_10),
.Y(n_319)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_12),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_12),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_12),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_12),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_12),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_12),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_12),
.B(n_429),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_13),
.Y(n_95)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_13),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_13),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_13),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_14),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_14),
.Y(n_377)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_14),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_15),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_15),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_15),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_15),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_15),
.B(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_468),
.Y(n_16)
);

OAI21xp33_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_225),
.B(n_465),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_182),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_SL g465 ( 
.A1(n_19),
.A2(n_466),
.B(n_467),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_140),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_20),
.B(n_140),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_103),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_21),
.B(n_104),
.C(n_118),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_67),
.C(n_84),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_22),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_49),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_23),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_37),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_28),
.A2(n_33),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_28),
.B(n_209),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_28),
.A2(n_33),
.B1(n_208),
.B2(n_209),
.Y(n_433)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_31),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.C(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_34),
.A2(n_37),
.B1(n_112),
.B2(n_115),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_34),
.B(n_277),
.C(n_281),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_34),
.A2(n_37),
.B1(n_281),
.B2(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_37),
.B(n_107),
.C(n_112),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_38),
.B(n_49),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_39),
.A2(n_122),
.B1(n_123),
.B2(n_130),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_39),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_39),
.A2(n_44),
.B1(n_130),
.B2(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_43),
.Y(n_331)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_46),
.Y(n_216)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_47),
.Y(n_350)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_48),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_48),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_61),
.B2(n_62),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_54),
.Y(n_249)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_54),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_55),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_55),
.B(n_59),
.C(n_62),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_55),
.B(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_60),
.B(n_195),
.C(n_200),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_61),
.A2(n_62),
.B1(n_477),
.B2(n_478),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_66),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_67),
.A2(n_84),
.B1(n_85),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_73),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_78),
.C(n_82),
.Y(n_120)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_72),
.Y(n_220)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_78),
.B1(n_82),
.B2(n_83),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_74),
.B(n_88),
.C(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_74),
.A2(n_82),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_77),
.Y(n_177)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_96),
.C(n_100),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_86),
.A2(n_87),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.C(n_94),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_88),
.A2(n_94),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_88),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_88),
.A2(n_164),
.B1(n_170),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_88),
.A2(n_164),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_88),
.B(n_392),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_90),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_90),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_90),
.B(n_247),
.C(n_250),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_90),
.A2(n_166),
.B1(n_247),
.B2(n_314),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_94),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_96),
.A2(n_100),
.B1(n_101),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_99),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_99),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_100),
.A2(n_101),
.B1(n_173),
.B2(n_223),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_169),
.C(n_173),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_118),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_116),
.C(n_117),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_107),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_106),
.B(n_235),
.C(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_106),
.A2(n_107),
.B1(n_235),
.B2(n_236),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_107),
.B(n_124),
.C(n_130),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_112),
.Y(n_115)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_117),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_131),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_120),
.B(n_121),
.C(n_131),
.Y(n_472)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_124),
.A2(n_125),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_124),
.A2(n_125),
.B1(n_153),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_125),
.B(n_208),
.C(n_214),
.Y(n_207)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_129),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_132),
.B(n_136),
.C(n_138),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_141),
.B(n_144),
.CI(n_146),
.CON(n_224),
.SN(n_224)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_168),
.C(n_178),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.C(n_162),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_148),
.B(n_152),
.Y(n_298)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.C(n_158),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_153),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_153),
.Y(n_479)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_158),
.Y(n_205)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_160),
.Y(n_486)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_162),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_178),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_170),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_170),
.A2(n_193),
.B1(n_285),
.B2(n_286),
.Y(n_357)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_171),
.Y(n_384)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_171),
.Y(n_406)
);

BUFx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_172),
.Y(n_414)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_177),
.Y(n_282)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_179),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_224),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_183),
.B(n_224),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_184),
.B(n_186),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_188),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_206),
.C(n_221),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_189),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.C(n_204),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_190),
.Y(n_270)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_194),
.B(n_204),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_206),
.B(n_221),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_215),
.C(n_217),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_207),
.B(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_208),
.A2(n_209),
.B1(n_214),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_213),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_214),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_224),
.Y(n_490)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_363),
.B1(n_458),
.B2(n_463),
.C(n_464),
.Y(n_225)
);

NOR3xp33_ASAP7_75t_SL g226 ( 
.A(n_227),
.B(n_302),
.C(n_306),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_227),
.A2(n_459),
.B(n_462),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_295),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_228),
.B(n_295),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_269),
.C(n_272),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_229),
.B(n_269),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_254),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_255),
.C(n_266),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.C(n_245),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_232),
.B(n_246),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_234),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_240),
.B(n_275),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g391 ( 
.A(n_244),
.Y(n_391)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_247),
.Y(n_314)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_250),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_266),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_261),
.C(n_264),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_256),
.A2(n_257),
.B(n_316),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_264),
.Y(n_294)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_263),
.B(n_317),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_289),
.C(n_293),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_273),
.B(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.C(n_283),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_274),
.B(n_359),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_276),
.A2(n_283),
.B1(n_284),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_277),
.B(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_301),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_299),
.C(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_302),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_303),
.B(n_304),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_336),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_307),
.A2(n_460),
.B(n_461),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_334),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_308),
.B(n_334),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.C(n_332),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_309),
.B(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_311),
.B(n_332),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_315),
.C(n_320),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_315),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.C(n_326),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_321),
.A2(n_322),
.B1(n_446),
.B2(n_447),
.Y(n_445)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_323),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_446)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_361),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_337),
.B(n_361),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.C(n_358),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_338),
.B(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_340),
.B(n_358),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_356),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_341),
.B(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_344),
.A2(n_356),
.B1(n_357),
.B2(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_344),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_348),
.C(n_351),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_345),
.A2(n_346),
.B1(n_351),
.B2(n_352),
.Y(n_438)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_348),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_453),
.B(n_457),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_440),
.B(n_452),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_424),
.B(n_439),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_400),
.B(n_423),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_368),
.B(n_393),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_393),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_380),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_369),
.B(n_381),
.C(n_389),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_376),
.C(n_378),
.Y(n_436)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_389),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_385),
.Y(n_394)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_390),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.C(n_396),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_395),
.Y(n_421)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_417),
.B(n_422),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_410),
.B(n_416),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_409),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_409),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_407),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_407),
.Y(n_418)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_415),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_413),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_419),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_426),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_435),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_427),
.A2(n_443),
.B1(n_444),
.B2(n_445),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_436),
.C(n_437),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_433),
.CI(n_434),
.CON(n_427),
.SN(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_451),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_441),
.B(n_451),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_448),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_443),
.B(n_445),
.C(n_448),
.Y(n_454)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_446),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_454),
.B(n_455),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_488),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_471),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_475),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_480),
.B1(n_481),
.B2(n_487),
.Y(n_475)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_476),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_482),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_483),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_485),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);


endmodule