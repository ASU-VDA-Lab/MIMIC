module fake_jpeg_31129_n_135 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_135);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_33),
.B(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_0),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_65),
.Y(n_71)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_56),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_56),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_66),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_72),
.B1(n_80),
.B2(n_18),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_46),
.B1(n_50),
.B2(n_49),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_24),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_64),
.A2(n_51),
.B1(n_47),
.B2(n_48),
.Y(n_75)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_52),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_3),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_19),
.B1(n_41),
.B2(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_71),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_85),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_84),
.B(n_5),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_3),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_94),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_23),
.C(n_39),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.C(n_6),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_4),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_97),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_108),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_109),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_8),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_14),
.B1(n_17),
.B2(n_26),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_121),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_29),
.C(n_31),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_122),
.B(n_35),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_SL g124 ( 
.A1(n_115),
.A2(n_99),
.A3(n_109),
.B1(n_107),
.B2(n_113),
.C1(n_103),
.C2(n_105),
.Y(n_124)
);

OAI322xp33_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_117),
.A3(n_116),
.B1(n_38),
.B2(n_42),
.C1(n_36),
.C2(n_37),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_123),
.A2(n_103),
.B(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_126),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_118),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_129),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_127),
.C(n_100),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_101),
.C(n_120),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_121),
.Y(n_135)
);


endmodule