module real_jpeg_18957_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_0),
.B(n_2),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_10),
.Y(n_9)
);

OR2x4_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_10),
.Y(n_21)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_13),
.Y(n_12)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_5),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_3),
.B(n_16),
.Y(n_15)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_7),
.B(n_23),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_11),
.B1(n_21),
.B2(n_22),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_9),
.Y(n_8)
);

AND2x4_ASAP7_75t_L g25 ( 
.A(n_10),
.B(n_26),
.Y(n_25)
);

OR2x4_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_18),
.Y(n_11)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_15),
.C(n_17),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_19),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2x1p5_ASAP7_75t_R g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);


endmodule