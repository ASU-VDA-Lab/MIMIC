module fake_netlist_5_2568_n_171 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_171);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_171;

wire n_137;
wire n_168;
wire n_164;
wire n_91;
wire n_122;
wire n_82;
wire n_142;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_146;
wire n_143;
wire n_132;
wire n_83;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_165;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_167;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_163;
wire n_95;
wire n_119;
wire n_169;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_162;
wire n_170;
wire n_77;
wire n_102;
wire n_106;
wire n_64;
wire n_161;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_141;
wire n_166;
wire n_97;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx2_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_0),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVxp67_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_0),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_32),
.B(n_1),
.C(n_2),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_37),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_35),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g74 ( 
.A(n_34),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_L g75 ( 
.A(n_33),
.B(n_5),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_56),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_47),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_58),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_44),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_73),
.A2(n_48),
.B1(n_46),
.B2(n_40),
.Y(n_92)
);

NOR2xp67_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_6),
.Y(n_93)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_60),
.B(n_65),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_59),
.B(n_71),
.Y(n_95)
);

OAI21x1_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_56),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_68),
.Y(n_97)
);

AOI21x1_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_59),
.B(n_66),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AO31x2_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_60),
.A3(n_65),
.B(n_69),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_68),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_90),
.A2(n_59),
.B(n_56),
.Y(n_102)
);

AOI221xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_76),
.B1(n_72),
.B2(n_62),
.C(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_90),
.A2(n_59),
.B(n_63),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_79),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_104),
.B(n_79),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_72),
.B1(n_92),
.B2(n_77),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_75),
.B(n_62),
.C(n_88),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_79),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_75),
.B(n_86),
.C(n_69),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_88),
.Y(n_111)
);

AND2x4_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_109),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_100),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_111),
.Y(n_119)
);

NOR2xp67_ASAP7_75t_L g120 ( 
.A(n_118),
.B(n_87),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_111),
.Y(n_123)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_119),
.A2(n_107),
.B1(n_113),
.B2(n_115),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

OAI31xp33_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_114),
.A3(n_108),
.B(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_113),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_118),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_105),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_74),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g138 ( 
.A1(n_128),
.A2(n_38),
.A3(n_40),
.B1(n_70),
.B2(n_61),
.C1(n_53),
.C2(n_69),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_74),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_64),
.A3(n_133),
.B1(n_65),
.B2(n_134),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_138),
.A2(n_93),
.B(n_126),
.Y(n_141)
);

NAND4xp25_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_93),
.C(n_70),
.D(n_110),
.Y(n_142)
);

NOR4xp25_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_110),
.C(n_136),
.D(n_135),
.Y(n_143)
);

AOI222xp33_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_61),
.B1(n_64),
.B2(n_124),
.C1(n_106),
.C2(n_130),
.Y(n_144)
);

OAI221xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_74),
.B1(n_126),
.B2(n_133),
.C(n_134),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_124),
.B1(n_130),
.B2(n_66),
.C(n_79),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_130),
.C(n_134),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g148 ( 
.A1(n_139),
.A2(n_131),
.B1(n_130),
.B2(n_116),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_141),
.B(n_131),
.Y(n_149)
);

OAI221xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_66),
.B1(n_116),
.B2(n_94),
.C(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_66),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_148),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_66),
.B(n_112),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_100),
.Y(n_156)
);

NAND4xp25_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_117),
.Y(n_159)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_11),
.Y(n_160)
);

NOR2x1_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_155),
.Y(n_161)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.C(n_83),
.Y(n_162)
);

AOI211xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_117),
.B(n_112),
.C(n_83),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_117),
.A3(n_112),
.B1(n_81),
.B2(n_80),
.C1(n_98),
.C2(n_20),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_162),
.A2(n_117),
.A3(n_112),
.B1(n_80),
.B2(n_21),
.C1(n_25),
.C2(n_24),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_158),
.A2(n_112),
.A3(n_82),
.B1(n_68),
.B2(n_85),
.C1(n_100),
.C2(n_84),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_160),
.B1(n_159),
.B2(n_94),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_94),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_164),
.B(n_166),
.Y(n_169)
);

AOI222xp33_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_168),
.B1(n_68),
.B2(n_84),
.C1(n_101),
.C2(n_97),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_170),
.A2(n_68),
.B1(n_84),
.B2(n_99),
.Y(n_171)
);


endmodule