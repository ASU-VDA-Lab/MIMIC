module fake_jpeg_23817_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_27),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_55),
.Y(n_70)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_15),
.Y(n_56)
);

HAxp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_57),
.CON(n_83),
.SN(n_83)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_15),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_15),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_25),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_66),
.Y(n_90)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_30),
.B1(n_28),
.B2(n_41),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_73),
.B1(n_78),
.B2(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_75),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_28),
.B1(n_41),
.B2(n_30),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_20),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

CKINVDCx12_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_77),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_28),
.B1(n_30),
.B2(n_26),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_82),
.Y(n_111)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVxp33_ASAP7_75t_SL g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_100),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_48),
.C(n_49),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_92),
.C(n_94),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_72),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_99),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_57),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_22),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_87),
.B(n_36),
.Y(n_118)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_30),
.B1(n_52),
.B2(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_127),
.C(n_129),
.Y(n_139)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_83),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_130),
.C(n_107),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_21),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_121),
.Y(n_152)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_126),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_56),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_136),
.Y(n_147)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_65),
.C(n_40),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_128),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_65),
.C(n_40),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_81),
.Y(n_143)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_137),
.Y(n_160)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_61),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_64),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_142),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_101),
.B1(n_88),
.B2(n_108),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_159),
.B1(n_120),
.B2(n_71),
.Y(n_168)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_145),
.Y(n_177)
);

AOI32xp33_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_103),
.A3(n_111),
.B1(n_55),
.B2(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_114),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_149),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_158),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_153),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_164),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_113),
.A2(n_55),
.B1(n_66),
.B2(n_84),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_156),
.A2(n_150),
.B1(n_123),
.B2(n_98),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

INVx6_ASAP7_75t_SL g185 ( 
.A(n_157),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_112),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_130),
.A2(n_82),
.B1(n_50),
.B2(n_69),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_110),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_34),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_116),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_162),
.Y(n_183)
);

NOR2x1_ASAP7_75t_R g164 ( 
.A(n_118),
.B(n_22),
.Y(n_164)
);

CKINVDCx12_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_171),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_129),
.C(n_117),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_176),
.C(n_19),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_22),
.B1(n_42),
.B2(n_45),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_168),
.A2(n_173),
.B(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_156),
.B1(n_161),
.B2(n_144),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_178),
.B1(n_188),
.B2(n_190),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_64),
.B1(n_134),
.B2(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_22),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_50),
.C(n_96),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_152),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_182),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_153),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_142),
.A2(n_126),
.B(n_122),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_131),
.B1(n_69),
.B2(n_62),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_147),
.A2(n_36),
.B1(n_22),
.B2(n_21),
.Y(n_190)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_162),
.B(n_147),
.C(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_140),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_197),
.C(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_22),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_34),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_195),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_187),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_210),
.B1(n_189),
.B2(n_184),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_17),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_33),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_176),
.C(n_170),
.Y(n_217)
);

NAND2xp33_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_10),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_204),
.A2(n_207),
.B1(n_175),
.B2(n_25),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_183),
.B(n_16),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_211),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_20),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_36),
.B(n_19),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_23),
.B(n_19),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_34),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_131),
.Y(n_214)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_214),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_199),
.C(n_198),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_218),
.A2(n_23),
.B1(n_29),
.B2(n_16),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_174),
.CI(n_180),
.CON(n_219),
.SN(n_219)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_20),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_167),
.B1(n_180),
.B2(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_182),
.B1(n_173),
.B2(n_62),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_198),
.A2(n_173),
.B(n_29),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_33),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_34),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_33),
.Y(n_244)
);

AOI21xp33_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_8),
.B(n_13),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_232),
.B(n_211),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_191),
.B1(n_201),
.B2(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_236),
.B(n_248),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_252),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_192),
.C(n_203),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_242),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_209),
.C(n_193),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_222),
.A2(n_206),
.B1(n_210),
.B2(n_62),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_251),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_221),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_250),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_102),
.C(n_45),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_39),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_39),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_226),
.C(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_229),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_17),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_242),
.B(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_250),
.A2(n_234),
.B(n_223),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_258),
.A2(n_259),
.B(n_16),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_219),
.B(n_224),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_224),
.C(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_266),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_45),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_239),
.A2(n_246),
.B1(n_237),
.B2(n_240),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_18),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_251),
.B1(n_80),
.B2(n_29),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_278),
.B1(n_269),
.B2(n_9),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_255),
.A2(n_261),
.B(n_260),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_39),
.C(n_37),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_281),
.C(n_283),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_11),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_SL g279 ( 
.A(n_263),
.B(n_9),
.C(n_13),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_9),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_39),
.C(n_37),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_284),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_37),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_18),
.Y(n_284)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_289),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_267),
.B1(n_24),
.B2(n_17),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_7),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_291),
.B(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_24),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_37),
.C(n_24),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_12),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_0),
.B(n_1),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_24),
.B1(n_17),
.B2(n_2),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_277),
.B1(n_272),
.B2(n_24),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_281),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_299),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_310)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_11),
.C(n_7),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_300),
.A2(n_303),
.B(n_1),
.Y(n_311)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_0),
.B(n_1),
.Y(n_305)
);

OA21x2_ASAP7_75t_SL g307 ( 
.A1(n_305),
.A2(n_1),
.B(n_2),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_292),
.B(n_285),
.Y(n_306)
);

OAI321xp33_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_307),
.A3(n_311),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_293),
.C(n_296),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_3),
.B(n_5),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_304),
.Y(n_312)
);

OAI22xp33_ASAP7_75t_L g315 ( 
.A1(n_312),
.A2(n_313),
.B1(n_314),
.B2(n_5),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_5),
.B(n_6),
.Y(n_316)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_306),
.C(n_6),
.Y(n_317)
);

AOI32xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_6),
.A3(n_18),
.B1(n_308),
.B2(n_286),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_6),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_18),
.Y(n_320)
);


endmodule