module real_jpeg_8785_n_21 (n_17, n_8, n_0, n_95, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_94, n_1, n_20, n_19, n_96, n_16, n_15, n_13, n_21);

input n_17;
input n_8;
input n_0;
input n_95;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_94;
input n_1;
input n_20;
input n_19;
input n_96;
input n_16;
input n_15;
input n_13;

output n_21;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_0),
.B(n_14),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_8),
.Y(n_47)
);

OAI221xp5_ASAP7_75t_L g43 ( 
.A1(n_2),
.A2(n_8),
.B1(n_31),
.B2(n_44),
.C(n_45),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_3),
.B(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_3),
.B(n_5),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_7),
.A2(n_8),
.B1(n_31),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_SL g37 ( 
.A(n_8),
.B(n_26),
.C(n_38),
.Y(n_37)
);

OAI221xp5_ASAP7_75t_L g39 ( 
.A1(n_8),
.A2(n_10),
.B1(n_31),
.B2(n_40),
.C(n_41),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_8),
.A2(n_16),
.B1(n_31),
.B2(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_19),
.B1(n_31),
.B2(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_8),
.A2(n_47),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_9),
.A2(n_23),
.B1(n_50),
.B2(n_51),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_51),
.B1(n_81),
.B2(n_91),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_12),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_13),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_15),
.A2(n_53),
.B1(n_60),
.B2(n_71),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_94),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_95),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_96),
.Y(n_66)
);

AOI221xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_52),
.B1(n_75),
.B2(n_80),
.C(n_92),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

NOR5xp2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.C(n_39),
.D(n_43),
.E(n_47),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_32),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_87),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_31),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_30),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_32),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_34),
.B(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR4xp25_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_83),
.C(n_89),
.D(n_90),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_77),
.B(n_79),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_72),
.B(n_74),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_72),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_67),
.B(n_70),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);


endmodule