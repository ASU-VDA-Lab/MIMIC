module real_jpeg_5776_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_1),
.A2(n_113),
.B1(n_116),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_1),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_1),
.A2(n_116),
.B1(n_289),
.B2(n_292),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_1),
.A2(n_49),
.B1(n_116),
.B2(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_1),
.A2(n_116),
.B1(n_358),
.B2(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_2),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_2),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_2),
.A2(n_35),
.B1(n_132),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_2),
.A2(n_132),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_2),
.A2(n_86),
.B1(n_132),
.B2(n_173),
.Y(n_391)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_4),
.A2(n_121),
.B1(n_123),
.B2(n_124),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_4),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_4),
.A2(n_123),
.B1(n_133),
.B2(n_216),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_4),
.A2(n_123),
.B1(n_296),
.B2(n_298),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_4),
.A2(n_123),
.B1(n_365),
.B2(n_366),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_5),
.A2(n_37),
.B1(n_172),
.B2(n_175),
.Y(n_171)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_7),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_7),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_8),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_8),
.A2(n_85),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_8),
.A2(n_85),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_9),
.A2(n_115),
.B1(n_243),
.B2(n_246),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_9),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_9),
.A2(n_86),
.B1(n_246),
.B2(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_9),
.A2(n_246),
.B1(n_316),
.B2(n_318),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_9),
.A2(n_155),
.B1(n_246),
.B2(n_360),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_10),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_10),
.Y(n_106)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_11),
.Y(n_104)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_12),
.Y(n_98)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_12),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_12),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_12),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_12),
.Y(n_245)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_47),
.B1(n_75),
.B2(n_79),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_14),
.A2(n_47),
.B1(n_146),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_15),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_15),
.B(n_265),
.C(n_269),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_15),
.A2(n_275),
.B1(n_276),
.B2(n_279),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_15),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_15),
.B(n_152),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_15),
.A2(n_24),
.B1(n_315),
.B2(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_15),
.B(n_204),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_15),
.A2(n_97),
.B(n_230),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_251),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_249),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_208),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_19),
.B(n_208),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_157),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_89),
.C(n_127),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_22),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_23),
.B(n_51),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_33),
.B(n_41),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_24),
.A2(n_161),
.B(n_165),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_24),
.B(n_43),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_24),
.A2(n_33),
.B1(n_234),
.B2(n_239),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_24),
.A2(n_184),
.B(n_295),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_24),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_24),
.A2(n_305),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_24),
.A2(n_41),
.B(n_165),
.Y(n_353)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_25),
.Y(n_306)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_27),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_29),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_42),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_30),
.A2(n_183),
.B(n_235),
.Y(n_381)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_32),
.Y(n_327)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_35),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_35),
.Y(n_238)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_36),
.Y(n_300)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_36),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_40),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_46),
.Y(n_168)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_73),
.B1(n_82),
.B2(n_88),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_52),
.A2(n_170),
.B(n_176),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_52),
.A2(n_388),
.B(n_389),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_52),
.A2(n_176),
.B(n_391),
.Y(n_404)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_53),
.A2(n_171),
.B1(n_177),
.B2(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_53),
.A2(n_177),
.B1(n_274),
.B2(n_280),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_53),
.A2(n_177),
.B1(n_280),
.B2(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_53),
.A2(n_177),
.B1(n_288),
.B2(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_66),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_61),
.B2(n_64),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_57),
.Y(n_279)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_57),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_57),
.Y(n_292)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_57),
.Y(n_352)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_63),
.Y(n_268)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_74),
.B(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_80),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_81),
.Y(n_174)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_81),
.Y(n_263)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_81),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_81),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_82),
.Y(n_189)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_87),
.A2(n_138),
.B1(n_139),
.B2(n_142),
.Y(n_137)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_87),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g177 ( 
.A(n_88),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_88),
.B(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_88),
.B(n_391),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_89),
.A2(n_90),
.B1(n_127),
.B2(n_128),
.Y(n_210)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_112),
.B1(n_120),
.B2(n_126),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_91),
.A2(n_120),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_91),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_91),
.A2(n_126),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_97),
.B2(n_99),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_107),
.B2(n_110),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_104),
.Y(n_222)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_109),
.Y(n_217)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_111),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_112),
.Y(n_248)
);

OAI32xp33_ASAP7_75t_L g220 ( 
.A1(n_113),
.A2(n_221),
.A3(n_223),
.B1(n_225),
.B2(n_229),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_124),
.Y(n_203)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_135),
.B(n_151),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_129),
.B(n_137),
.Y(n_218)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_131),
.Y(n_146)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_135),
.A2(n_137),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_135),
.A2(n_137),
.B1(n_376),
.B2(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_136),
.B(n_153),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_136),
.A2(n_215),
.B(n_218),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_136),
.A2(n_152),
.B1(n_356),
.B2(n_359),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_145),
.Y(n_136)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_137),
.A2(n_192),
.B(n_196),
.Y(n_191)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_141),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_141),
.Y(n_348)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_150),
.Y(n_145)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_149),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_149),
.Y(n_362)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_150),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_155),
.A2(n_340),
.A3(n_342),
.B1(n_343),
.B2(n_346),
.Y(n_339)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_179),
.B1(n_206),
.B2(n_207),
.Y(n_157)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_169),
.B2(n_178),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_161),
.Y(n_309)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_181),
.A2(n_187),
.B1(n_188),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_197),
.B1(n_198),
.B2(n_205),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_204),
.Y(n_199)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_204),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.C(n_213),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_209),
.B(n_211),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_213),
.B(n_417),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.C(n_241),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_214),
.B(n_241),
.Y(n_413)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_215),
.Y(n_403)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_219),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_233),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_220),
.B(n_233),
.Y(n_399)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_242),
.Y(n_407)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_409),
.B(n_422),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_395),
.B(n_408),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_369),
.B(n_394),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_335),
.B(n_368),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_301),
.B(n_334),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_283),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_258),
.B(n_283),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_273),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_259),
.B(n_273),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_275),
.B(n_344),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_SL g356 ( 
.A1(n_275),
.A2(n_343),
.B(n_357),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_294),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_293),
.C(n_294),
.Y(n_336)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_287),
.Y(n_293)
);

INVx4_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_311),
.B(n_333),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_310),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_310),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_312),
.A2(n_321),
.B(n_332),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_313),
.B(n_314),
.Y(n_332)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_319),
.Y(n_324)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_337),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_354),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_355),
.C(n_363),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_353),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_353),
.Y(n_386)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_351),
.Y(n_365)
);

INVx4_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_363),
.Y(n_354)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_359),
.Y(n_375)
);

INVx5_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_362),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_364),
.Y(n_388)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_370),
.B(n_371),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_384),
.B2(n_385),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_387),
.C(n_392),
.Y(n_396)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_379),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_380),
.C(n_383),
.Y(n_400)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_382),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_392),
.B2(n_393),
.Y(n_385)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_386),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_387),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_397),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_401),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_400),
.C(n_401),
.Y(n_419)
);

BUFx24_ASAP7_75t_SL g426 ( 
.A(n_401),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_404),
.CI(n_405),
.CON(n_401),
.SN(n_401)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_418),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_410),
.A2(n_423),
.B(n_424),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_416),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_411),
.B(n_416),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.C(n_415),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_414),
.B(n_415),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_420),
.Y(n_423)
);


endmodule