module real_aes_1842_n_350 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_350);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_350;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_980;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_963;
wire n_865;
wire n_666;
wire n_551;
wire n_537;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_889;
wire n_696;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_892;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_872;
wire n_636;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_680;
wire n_595;
wire n_726;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_860;
wire n_748;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_936;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_947;
wire n_561;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_756;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_831;
wire n_487;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_359;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_371;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_842;
wire n_849;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_0), .A2(n_301), .B1(n_545), .B2(n_581), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_1), .A2(n_199), .B1(n_551), .B2(n_552), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g738 ( .A1(n_2), .A2(n_249), .B1(n_412), .B2(n_416), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g627 ( .A1(n_3), .A2(n_147), .B1(n_459), .B2(n_460), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_4), .A2(n_111), .B1(n_435), .B2(n_438), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_5), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g517 ( .A1(n_6), .A2(n_177), .B1(n_472), .B2(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_7), .B(n_631), .Y(n_921) );
AOI22xp33_ASAP7_75t_SL g689 ( .A1(n_8), .A2(n_229), .B1(n_545), .B2(n_581), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_9), .A2(n_299), .B1(n_426), .B2(n_666), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_10), .A2(n_171), .B1(n_481), .B2(n_524), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_11), .A2(n_254), .B1(n_422), .B2(n_425), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_12), .A2(n_335), .B1(n_614), .B2(n_615), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_13), .A2(n_184), .B1(n_547), .B2(n_548), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_14), .A2(n_78), .B1(n_439), .B2(n_524), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g574 ( .A1(n_15), .A2(n_80), .B1(n_540), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_16), .A2(n_226), .B1(n_539), .B2(n_661), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_17), .A2(n_296), .B1(n_429), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_18), .A2(n_174), .B1(n_403), .B2(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_19), .A2(n_167), .B1(n_771), .B2(n_915), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_20), .A2(n_201), .B1(n_536), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_21), .A2(n_160), .B1(n_441), .B2(n_445), .Y(n_440) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_22), .A2(n_158), .B1(n_552), .B2(n_555), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_23), .A2(n_324), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_24), .A2(n_131), .B1(n_398), .B2(n_467), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_25), .A2(n_60), .B1(n_412), .B2(n_658), .Y(n_657) );
AO222x2_ASAP7_75t_L g809 ( .A1(n_26), .A2(n_126), .B1(n_215), .B2(n_530), .C1(n_532), .C2(n_533), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_27), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_28), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_29), .A2(n_310), .B1(n_536), .B2(n_537), .Y(n_812) );
INVx1_ASAP7_75t_SL g380 ( .A(n_30), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g944 ( .A(n_30), .B(n_44), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_31), .A2(n_318), .B1(n_429), .B2(n_432), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_32), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g857 ( .A1(n_33), .A2(n_155), .B1(n_722), .B2(n_754), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_34), .A2(n_117), .B1(n_459), .B2(n_506), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_35), .B(n_464), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_36), .A2(n_265), .B1(n_547), .B2(n_548), .Y(n_933) );
AOI22x1_ASAP7_75t_L g584 ( .A1(n_37), .A2(n_179), .B1(n_547), .B2(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_38), .A2(n_105), .B1(n_536), .B2(n_537), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_39), .A2(n_198), .B1(n_639), .B2(n_773), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_40), .A2(n_195), .B1(n_467), .B2(n_615), .Y(n_761) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_41), .A2(n_351), .B(n_360), .C(n_945), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_42), .A2(n_170), .B1(n_575), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_43), .A2(n_300), .B1(n_476), .B2(n_477), .Y(n_602) );
AO22x2_ASAP7_75t_L g382 ( .A1(n_44), .A2(n_329), .B1(n_379), .B2(n_383), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_45), .A2(n_154), .B1(n_781), .B2(n_915), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_46), .A2(n_191), .B1(n_425), .B2(n_600), .Y(n_950) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_47), .A2(n_54), .B1(n_412), .B2(n_416), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_48), .A2(n_298), .B1(n_425), .B2(n_600), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_49), .A2(n_163), .B1(n_407), .B2(n_498), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_50), .A2(n_255), .B1(n_476), .B2(n_667), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_51), .B(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g381 ( .A(n_52), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_53), .A2(n_281), .B1(n_548), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_55), .A2(n_278), .B1(n_547), .B2(n_554), .Y(n_690) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_56), .A2(n_287), .B1(n_476), .B2(n_637), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g770 ( .A1(n_57), .A2(n_125), .B1(n_671), .B2(n_771), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_58), .A2(n_326), .B1(n_771), .B2(n_835), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_59), .A2(n_273), .B1(n_601), .B2(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_61), .A2(n_222), .B1(n_403), .B2(n_456), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_62), .A2(n_323), .B1(n_480), .B2(n_609), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_63), .A2(n_193), .B1(n_480), .B2(n_481), .Y(n_479) );
AO22x2_ASAP7_75t_L g389 ( .A1(n_64), .A2(n_176), .B1(n_379), .B2(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_65), .A2(n_282), .B1(n_425), .B2(n_441), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_66), .A2(n_139), .B1(n_552), .B2(n_694), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_67), .A2(n_124), .B1(n_548), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_68), .A2(n_214), .B1(n_429), .B2(n_639), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_69), .A2(n_128), .B1(n_637), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_70), .A2(n_99), .B1(n_572), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_71), .A2(n_144), .B1(n_540), .B2(n_575), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_72), .A2(n_148), .B1(n_548), .B2(n_554), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_73), .A2(n_293), .B1(n_585), .B2(n_878), .Y(n_911) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_74), .A2(n_182), .B1(n_476), .B2(n_477), .Y(n_475) );
AOI22xp33_ASAP7_75t_SL g772 ( .A1(n_75), .A2(n_303), .B1(n_773), .B2(n_775), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_76), .A2(n_136), .B1(n_585), .B2(n_915), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_77), .A2(n_103), .B1(n_545), .B2(n_581), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_79), .A2(n_260), .B1(n_554), .B2(n_555), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_81), .A2(n_225), .B1(n_532), .B2(n_572), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_82), .B(n_502), .Y(n_501) );
XOR2xp5_ASAP7_75t_L g766 ( .A(n_83), .B(n_767), .Y(n_766) );
OAI22x1_ASAP7_75t_L g799 ( .A1(n_83), .A2(n_767), .B1(n_800), .B2(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_83), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_84), .A2(n_213), .B1(n_600), .B2(n_601), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_85), .A2(n_340), .B1(n_403), .B2(n_407), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g957 ( .A1(n_86), .A2(n_275), .B1(n_614), .B2(n_710), .Y(n_957) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_87), .A2(n_252), .B1(n_473), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_88), .A2(n_118), .B1(n_483), .B2(n_484), .Y(n_482) );
AO222x2_ASAP7_75t_L g683 ( .A1(n_89), .A2(n_190), .B1(n_332), .B2(n_530), .C1(n_540), .C2(n_577), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_90), .A2(n_112), .B1(n_724), .B2(n_726), .Y(n_723) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_91), .A2(n_211), .B1(n_577), .B2(n_925), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_92), .A2(n_212), .B1(n_498), .B2(n_500), .Y(n_497) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_93), .A2(n_232), .B1(n_532), .B2(n_572), .Y(n_686) );
AOI222xp33_ASAP7_75t_L g958 ( .A1(n_94), .A2(n_156), .B1(n_316), .B2(n_407), .C1(n_760), .C2(n_959), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_95), .A2(n_138), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_96), .A2(n_122), .B1(n_412), .B2(n_459), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_97), .A2(n_116), .B1(n_779), .B2(n_780), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_98), .A2(n_192), .B1(n_794), .B2(n_795), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_100), .A2(n_307), .B1(n_667), .B2(n_835), .Y(n_913) );
AO22x2_ASAP7_75t_L g386 ( .A1(n_101), .A2(n_258), .B1(n_379), .B2(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_102), .A2(n_272), .B1(n_392), .B2(n_398), .Y(n_391) );
OAI22x1_ASAP7_75t_L g654 ( .A1(n_104), .A2(n_655), .B1(n_674), .B2(n_675), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g675 ( .A(n_104), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_106), .A2(n_134), .B1(n_392), .B2(n_468), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_107), .A2(n_345), .B1(n_722), .B2(n_835), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_108), .A2(n_242), .B1(n_435), .B2(n_438), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_109), .A2(n_218), .B1(n_459), .B2(n_460), .Y(n_612) );
XOR2xp5_ASAP7_75t_L g946 ( .A(n_110), .B(n_947), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_113), .A2(n_322), .B1(n_544), .B2(n_545), .Y(n_543) );
OA22x2_ASAP7_75t_L g491 ( .A1(n_114), .A2(n_492), .B1(n_493), .B2(n_494), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_114), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_115), .A2(n_186), .B1(n_551), .B2(n_552), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_119), .A2(n_153), .B1(n_521), .B2(n_522), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g934 ( .A(n_120), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_121), .A2(n_245), .B1(n_403), .B2(n_407), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_123), .A2(n_207), .B1(n_435), .B2(n_756), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_127), .A2(n_151), .B1(n_467), .B2(n_468), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_129), .A2(n_135), .B1(n_554), .B2(n_555), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_130), .A2(n_305), .B1(n_459), .B2(n_460), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_132), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_133), .A2(n_217), .B1(n_403), .B2(n_500), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_137), .A2(n_202), .B1(n_666), .B2(n_667), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_140), .A2(n_346), .B1(n_477), .B2(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_141), .B(n_502), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_142), .A2(n_261), .B1(n_432), .B2(n_472), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_143), .A2(n_337), .B1(n_710), .B2(n_711), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_145), .B(n_372), .Y(n_371) );
AOI22xp33_ASAP7_75t_SL g910 ( .A1(n_146), .A2(n_291), .B1(n_429), .B2(n_431), .Y(n_910) );
OA22x2_ASAP7_75t_L g966 ( .A1(n_149), .A2(n_967), .B1(n_979), .B2(n_980), .Y(n_966) );
INVx1_ASAP7_75t_L g979 ( .A(n_149), .Y(n_979) );
AOI22xp33_ASAP7_75t_SL g638 ( .A1(n_150), .A2(n_274), .B1(n_429), .B2(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g621 ( .A(n_152), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_157), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_159), .A2(n_317), .B1(n_585), .B2(n_671), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_161), .B(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g891 ( .A1(n_162), .A2(n_347), .B1(n_785), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_164), .A2(n_189), .B1(n_412), .B2(n_459), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_165), .A2(n_233), .B1(n_412), .B2(n_416), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_166), .A2(n_239), .B1(n_412), .B2(n_416), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_168), .A2(n_302), .B1(n_484), .B2(n_702), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_169), .A2(n_262), .B1(n_500), .B2(n_786), .Y(n_971) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_172), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_173), .A2(n_284), .B1(n_441), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_175), .A2(n_227), .B1(n_831), .B2(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g943 ( .A(n_176), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_178), .A2(n_210), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_180), .A2(n_234), .B1(n_545), .B2(n_581), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_181), .A2(n_283), .B1(n_710), .B2(n_798), .Y(n_797) );
XNOR2xp5_ASAP7_75t_L g562 ( .A(n_183), .B(n_563), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_185), .A2(n_330), .B1(n_412), .B2(n_658), .Y(n_829) );
INVx1_ASAP7_75t_L g733 ( .A(n_187), .Y(n_733) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_188), .A2(n_290), .B1(n_536), .B2(n_539), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_194), .A2(n_251), .B1(n_875), .B2(n_876), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_196), .A2(n_286), .B1(n_756), .B2(n_878), .Y(n_877) );
OA22x2_ASAP7_75t_L g595 ( .A1(n_197), .A2(n_596), .B1(n_597), .B2(n_618), .Y(n_595) );
INVxp67_ASAP7_75t_L g618 ( .A(n_197), .Y(n_618) );
INVx2_ASAP7_75t_L g357 ( .A(n_200), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_203), .A2(n_341), .B1(n_552), .B2(n_694), .Y(n_818) );
OA22x2_ASAP7_75t_L g451 ( .A1(n_204), .A2(n_452), .B1(n_486), .B2(n_487), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_204), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g859 ( .A1(n_205), .A2(n_246), .B1(n_435), .B2(n_860), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_206), .A2(n_219), .B1(n_480), .B2(n_781), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g787 ( .A(n_208), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_209), .A2(n_228), .B1(n_459), .B2(n_506), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_216), .A2(n_253), .B1(n_472), .B2(n_473), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g556 ( .A(n_220), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_221), .A2(n_717), .B1(n_718), .B2(n_740), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_221), .Y(n_717) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_223), .A2(n_680), .B1(n_681), .B2(n_695), .Y(n_679) );
INVx1_ASAP7_75t_L g695 ( .A(n_223), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_224), .A2(n_315), .B1(n_711), .B2(n_907), .Y(n_906) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_230), .A2(n_311), .B1(n_532), .B2(n_533), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_231), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_235), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g848 ( .A1(n_236), .A2(n_243), .B1(n_403), .B2(n_407), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_237), .A2(n_256), .B1(n_539), .B2(n_540), .Y(n_811) );
AO22x2_ASAP7_75t_L g749 ( .A1(n_238), .A2(n_750), .B1(n_764), .B2(n_765), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_238), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_240), .A2(n_349), .B1(n_551), .B2(n_552), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_241), .A2(n_270), .B1(n_407), .B2(n_498), .Y(n_826) );
AOI22x1_ASAP7_75t_L g841 ( .A1(n_244), .A2(n_842), .B1(n_843), .B2(n_862), .Y(n_841) );
INVx1_ASAP7_75t_L g862 ( .A(n_244), .Y(n_862) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_247), .A2(n_328), .B1(n_601), .B2(n_671), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_248), .A2(n_325), .B1(n_431), .B2(n_472), .Y(n_705) );
OA22x2_ASAP7_75t_L g869 ( .A1(n_250), .A2(n_870), .B1(n_871), .B2(n_872), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_250), .Y(n_870) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_257), .A2(n_304), .B1(n_422), .B2(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_258), .B(n_942), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_259), .A2(n_327), .B1(n_403), .B2(n_500), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_263), .B(n_373), .Y(n_972) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_264), .A2(n_271), .B1(n_312), .B2(n_530), .C1(n_533), .C2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_266), .A2(n_314), .B1(n_552), .B2(n_694), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_267), .B(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_268), .A2(n_348), .B1(n_429), .B2(n_431), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_269), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_276), .Y(n_847) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_277), .A2(n_292), .B1(n_431), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_279), .A2(n_294), .B1(n_431), .B2(n_976), .Y(n_975) );
INVx3_ASAP7_75t_L g379 ( .A(n_280), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_285), .A2(n_295), .B1(n_552), .B2(n_694), .Y(n_932) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_288), .A2(n_336), .B1(n_393), .B2(n_615), .Y(n_628) );
OAI22x1_ASAP7_75t_L g368 ( .A1(n_289), .A2(n_369), .B1(n_448), .B2(n_449), .Y(n_368) );
INVx1_ASAP7_75t_L g449 ( .A(n_289), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g840 ( .A(n_297), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_306), .A2(n_333), .B1(n_658), .B2(n_889), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_308), .A2(n_338), .B1(n_425), .B2(n_476), .Y(n_752) );
XNOR2x1_ASAP7_75t_L g697 ( .A(n_309), .B(n_698), .Y(n_697) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_313), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_319), .Y(n_512) );
INVx1_ASAP7_75t_L g897 ( .A(n_320), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_321), .A2(n_344), .B1(n_467), .B2(n_831), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_331), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g939 ( .A(n_331), .Y(n_939) );
INVx1_ASAP7_75t_L g354 ( .A(n_334), .Y(n_354) );
AND2x2_ASAP7_75t_R g961 ( .A(n_334), .B(n_939), .Y(n_961) );
INVxp67_ASAP7_75t_L g359 ( .A(n_339), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_342), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_343), .B(n_502), .Y(n_707) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2x1_ASAP7_75t_R g352 ( .A(n_353), .B(n_355), .Y(n_352) );
OR2x2_ASAP7_75t_L g984 ( .A(n_353), .B(n_356), .Y(n_984) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_354), .B(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B1(n_647), .B2(n_935), .C(n_936), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_590), .B1(n_591), .B2(n_646), .Y(n_363) );
INVx1_ASAP7_75t_L g646 ( .A(n_364), .Y(n_646) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_489), .B(n_587), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g589 ( .A(n_366), .Y(n_589) );
AO22x2_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_450), .B2(n_451), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g448 ( .A(n_369), .Y(n_448) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_420), .Y(n_369) );
NAND4xp25_ASAP7_75t_L g370 ( .A(n_371), .B(n_391), .C(n_402), .D(n_411), .Y(n_370) );
INVx3_ASAP7_75t_L g734 ( .A(n_372), .Y(n_734) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g885 ( .A(n_373), .Y(n_885) );
INVx3_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVx3_ASAP7_75t_L g464 ( .A(n_374), .Y(n_464) );
INVx3_ASAP7_75t_L g502 ( .A(n_374), .Y(n_502) );
INVx4_ASAP7_75t_SL g631 ( .A(n_374), .Y(n_631) );
INVx4_ASAP7_75t_SL g760 ( .A(n_374), .Y(n_760) );
BUFx2_ASAP7_75t_L g788 ( .A(n_374), .Y(n_788) );
INVx6_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_384), .Y(n_375) );
AND2x4_ASAP7_75t_L g400 ( .A(n_376), .B(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g417 ( .A(n_376), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g530 ( .A(n_376), .B(n_384), .Y(n_530) );
AND2x2_ASAP7_75t_L g537 ( .A(n_376), .B(n_418), .Y(n_537) );
AND2x2_ASAP7_75t_L g540 ( .A(n_376), .B(n_401), .Y(n_540) );
AND2x2_ASAP7_75t_L g577 ( .A(n_376), .B(n_418), .Y(n_577) );
AND2x2_ASAP7_75t_L g661 ( .A(n_376), .B(n_401), .Y(n_661) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_382), .Y(n_376) );
INVx2_ASAP7_75t_L g397 ( .A(n_377), .Y(n_397) );
AND2x2_ASAP7_75t_L g405 ( .A(n_377), .B(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_377), .Y(n_410) );
OAI22x1_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_379), .B1(n_380), .B2(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g383 ( .A(n_379), .Y(n_383) );
INVx2_ASAP7_75t_L g387 ( .A(n_379), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_379), .Y(n_390) );
AND2x2_ASAP7_75t_L g396 ( .A(n_382), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g406 ( .A(n_382), .Y(n_406) );
BUFx2_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
AND2x2_ASAP7_75t_L g424 ( .A(n_384), .B(n_396), .Y(n_424) );
AND2x4_ASAP7_75t_L g437 ( .A(n_384), .B(n_405), .Y(n_437) );
AND2x4_ASAP7_75t_L g444 ( .A(n_384), .B(n_427), .Y(n_444) );
AND2x6_ASAP7_75t_L g547 ( .A(n_384), .B(n_396), .Y(n_547) );
AND2x2_ASAP7_75t_L g551 ( .A(n_384), .B(n_405), .Y(n_551) );
AND2x2_ASAP7_75t_L g554 ( .A(n_384), .B(n_427), .Y(n_554) );
AND2x2_ASAP7_75t_L g694 ( .A(n_384), .B(n_405), .Y(n_694) );
AND2x4_ASAP7_75t_L g384 ( .A(n_385), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g395 ( .A(n_386), .B(n_388), .Y(n_395) );
AND2x2_ASAP7_75t_L g409 ( .A(n_386), .B(n_389), .Y(n_409) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
INVxp67_ASAP7_75t_L g401 ( .A(n_388), .Y(n_401) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g414 ( .A(n_389), .B(n_415), .Y(n_414) );
BUFx4f_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g511 ( .A(n_393), .Y(n_511) );
BUFx2_ASAP7_75t_L g798 ( .A(n_393), .Y(n_798) );
BUFx2_ASAP7_75t_L g887 ( .A(n_393), .Y(n_887) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx3_ASAP7_75t_L g467 ( .A(n_394), .Y(n_467) );
BUFx2_ASAP7_75t_L g614 ( .A(n_394), .Y(n_614) );
BUFx2_ASAP7_75t_L g711 ( .A(n_394), .Y(n_711) );
AND2x4_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g404 ( .A(n_395), .B(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g426 ( .A(n_395), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g532 ( .A(n_395), .B(n_405), .Y(n_532) );
AND2x2_ASAP7_75t_L g539 ( .A(n_395), .B(n_396), .Y(n_539) );
AND2x2_ASAP7_75t_L g555 ( .A(n_395), .B(n_427), .Y(n_555) );
AND2x2_ASAP7_75t_L g575 ( .A(n_395), .B(n_396), .Y(n_575) );
AND2x2_ASAP7_75t_L g430 ( .A(n_396), .B(n_414), .Y(n_430) );
AND2x2_ASAP7_75t_L g544 ( .A(n_396), .B(n_414), .Y(n_544) );
AND2x2_ASAP7_75t_SL g581 ( .A(n_396), .B(n_414), .Y(n_581) );
AND2x4_ASAP7_75t_L g427 ( .A(n_397), .B(n_406), .Y(n_427) );
INVx2_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_SL g468 ( .A(n_399), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_399), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVx1_ASAP7_75t_L g615 ( .A(n_399), .Y(n_615) );
INVx2_ASAP7_75t_L g710 ( .A(n_399), .Y(n_710) );
INVx2_ASAP7_75t_L g831 ( .A(n_399), .Y(n_831) );
INVx2_ASAP7_75t_L g907 ( .A(n_399), .Y(n_907) );
INVx6_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx5_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g499 ( .A(n_404), .Y(n_499) );
BUFx3_ASAP7_75t_L g786 ( .A(n_404), .Y(n_786) );
AND2x2_ASAP7_75t_L g413 ( .A(n_405), .B(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g536 ( .A(n_405), .B(n_414), .Y(n_536) );
INVx2_ASAP7_75t_L g791 ( .A(n_407), .Y(n_791) );
BUFx3_ASAP7_75t_L g892 ( .A(n_407), .Y(n_892) );
BUFx12f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
AND2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
AND2x4_ASAP7_75t_L g432 ( .A(n_409), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g439 ( .A(n_409), .B(n_427), .Y(n_439) );
AND2x2_ASAP7_75t_SL g533 ( .A(n_409), .B(n_410), .Y(n_533) );
AND2x4_ASAP7_75t_L g545 ( .A(n_409), .B(n_433), .Y(n_545) );
AND2x4_ASAP7_75t_L g552 ( .A(n_409), .B(n_427), .Y(n_552) );
AND2x2_ASAP7_75t_SL g572 ( .A(n_409), .B(n_410), .Y(n_572) );
BUFx6f_ASAP7_75t_SL g794 ( .A(n_412), .Y(n_794) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx3_ASAP7_75t_L g461 ( .A(n_413), .Y(n_461) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_413), .Y(n_506) );
AND2x4_ASAP7_75t_L g447 ( .A(n_414), .B(n_427), .Y(n_447) );
AND2x6_ASAP7_75t_L g548 ( .A(n_414), .B(n_427), .Y(n_548) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_415), .Y(n_419) );
BUFx4f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_SL g459 ( .A(n_417), .Y(n_459) );
INVx2_ASAP7_75t_L g659 ( .A(n_417), .Y(n_659) );
INVx1_ASAP7_75t_L g796 ( .A(n_417), .Y(n_796) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g420 ( .A(n_421), .B(n_428), .C(n_434), .D(n_440), .Y(n_420) );
INVx2_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g483 ( .A(n_423), .Y(n_483) );
INVx2_ASAP7_75t_L g600 ( .A(n_423), .Y(n_600) );
INVx2_ASAP7_75t_SL g754 ( .A(n_423), .Y(n_754) );
INVx3_ASAP7_75t_L g835 ( .A(n_423), .Y(n_835) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx2_ASAP7_75t_L g516 ( .A(n_424), .Y(n_516) );
BUFx2_ASAP7_75t_L g666 ( .A(n_424), .Y(n_666) );
BUFx2_ASAP7_75t_L g876 ( .A(n_425), .Y(n_876) );
BUFx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g485 ( .A(n_426), .Y(n_485) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_426), .Y(n_585) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_426), .Y(n_601) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
INVx2_ASAP7_75t_L g606 ( .A(n_430), .Y(n_606) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx5_ASAP7_75t_SL g474 ( .A(n_432), .Y(n_474) );
BUFx3_ASAP7_75t_L g518 ( .A(n_432), .Y(n_518) );
BUFx2_ASAP7_75t_L g664 ( .A(n_432), .Y(n_664) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g480 ( .A(n_436), .Y(n_480) );
INVx3_ASAP7_75t_L g608 ( .A(n_436), .Y(n_608) );
INVx1_ASAP7_75t_SL g779 ( .A(n_436), .Y(n_779) );
INVx6_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx3_ASAP7_75t_L g524 ( .A(n_437), .Y(n_524) );
BUFx3_ASAP7_75t_L g878 ( .A(n_437), .Y(n_878) );
BUFx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
INVx2_ASAP7_75t_L g610 ( .A(n_439), .Y(n_610) );
BUFx3_ASAP7_75t_L g781 ( .A(n_439), .Y(n_781) );
BUFx2_ASAP7_75t_SL g860 ( .A(n_439), .Y(n_860) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_SL g476 ( .A(n_443), .Y(n_476) );
INVx2_ASAP7_75t_SL g521 ( .A(n_443), .Y(n_521) );
INVx2_ASAP7_75t_L g671 ( .A(n_443), .Y(n_671) );
INVx3_ASAP7_75t_SL g915 ( .A(n_443), .Y(n_915) );
INVx8_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
INVx1_ASAP7_75t_SL g637 ( .A(n_446), .Y(n_637) );
INVx2_ASAP7_75t_L g667 ( .A(n_446), .Y(n_667) );
INVx2_ASAP7_75t_SL g722 ( .A(n_446), .Y(n_722) );
INVx2_ASAP7_75t_SL g771 ( .A(n_446), .Y(n_771) );
INVx8_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AO22x2_ASAP7_75t_SL g619 ( .A1(n_450), .A2(n_451), .B1(n_620), .B2(n_644), .Y(n_619) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_469), .Y(n_452) );
NOR3xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_462), .C(n_465), .Y(n_453) );
NOR4xp25_ASAP7_75t_L g487 ( .A(n_454), .B(n_470), .C(n_478), .D(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_458), .Y(n_454) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g500 ( .A(n_457), .Y(n_500) );
INVx3_ASAP7_75t_L g736 ( .A(n_457), .Y(n_736) );
INVxp67_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g890 ( .A(n_461), .Y(n_890) );
INVx4_ASAP7_75t_L g925 ( .A(n_461), .Y(n_925) );
INVxp67_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_463), .B(n_466), .Y(n_488) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_478), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_475), .Y(n_470) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g639 ( .A(n_474), .Y(n_639) );
INVx2_ASAP7_75t_L g726 ( .A(n_474), .Y(n_726) );
INVx2_ASAP7_75t_L g775 ( .A(n_474), .Y(n_775) );
BUFx2_ASAP7_75t_L g875 ( .A(n_476), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_482), .Y(n_478) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g522 ( .A(n_485), .Y(n_522) );
INVx1_ASAP7_75t_L g729 ( .A(n_485), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_489), .B(n_588), .Y(n_587) );
XNOR2x1_ASAP7_75t_L g489 ( .A(n_490), .B(n_559), .Y(n_489) );
AO22x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_525), .B1(n_557), .B2(n_558), .Y(n_490) );
INVx1_ASAP7_75t_L g557 ( .A(n_491), .Y(n_557) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_513), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_503), .C(n_509), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g959 ( .A(n_499), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_507), .B2(n_508), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_519), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_517), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_523), .Y(n_519) );
INVx1_ASAP7_75t_L g558 ( .A(n_525), .Y(n_558) );
XOR2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_556), .Y(n_525) );
NAND2x1p5_ASAP7_75t_L g526 ( .A(n_527), .B(n_541), .Y(n_526) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx2_ASAP7_75t_SL g567 ( .A(n_530), .Y(n_567) );
INVx1_ASAP7_75t_SL g569 ( .A(n_532), .Y(n_569) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_532), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_549), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
INVx1_ASAP7_75t_L g703 ( .A(n_547), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_553), .Y(n_549) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g563 ( .A(n_564), .B(n_578), .Y(n_563) );
NOR2x1_ASAP7_75t_L g564 ( .A(n_565), .B(n_573), .Y(n_564) );
OAI222xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_568), .B2(n_569), .C1(n_570), .C2(n_571), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g900 ( .A1(n_567), .A2(n_901), .B(n_902), .Y(n_900) );
INVx1_ASAP7_75t_L g903 ( .A(n_569), .Y(n_903) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_583), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_582), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_619), .B(n_645), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_593), .B(n_619), .Y(n_645) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_611), .Y(n_597) );
NAND4xp25_ASAP7_75t_SL g598 ( .A(n_599), .B(n_602), .C(n_603), .D(n_607), .Y(n_598) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g725 ( .A(n_605), .Y(n_725) );
INVx1_ASAP7_75t_L g856 ( .A(n_605), .Y(n_856) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g774 ( .A(n_606), .Y(n_774) );
INVx1_ASAP7_75t_L g976 ( .A(n_606), .Y(n_976) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g756 ( .A(n_610), .Y(n_756) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .C(n_616), .D(n_617), .Y(n_611) );
INVx2_ASAP7_75t_L g644 ( .A(n_620), .Y(n_644) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_643), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_621), .B(n_624), .Y(n_643) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_634), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_629), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_628), .Y(n_626) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_632), .B(n_633), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_635), .B(n_640), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g935 ( .A(n_647), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_743), .B2(n_744), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AO22x1_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B1(n_713), .B2(n_741), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AO22x2_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_676), .B2(n_677), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND4xp25_ASAP7_75t_SL g655 ( .A(n_656), .B(n_662), .C(n_668), .D(n_672), .Y(n_655) );
AND4x1_ASAP7_75t_L g674 ( .A(n_656), .B(n_662), .C(n_668), .D(n_672), .Y(n_674) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OA22x2_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_679), .B1(n_696), .B2(n_697), .Y(n_677) );
INVx1_ASAP7_75t_L g715 ( .A(n_678), .Y(n_715) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_682), .B(n_687), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
NOR2x1_ASAP7_75t_L g698 ( .A(n_699), .B(n_706), .Y(n_698) );
NAND4xp25_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .C(n_704), .D(n_705), .Y(n_699) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND4xp25_ASAP7_75t_SL g706 ( .A(n_707), .B(n_708), .C(n_709), .D(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx3_ASAP7_75t_L g742 ( .A(n_714), .Y(n_742) );
XNOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
INVx1_ASAP7_75t_SL g740 ( .A(n_718), .Y(n_740) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_731), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_727), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_730), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_737), .Y(n_731) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_735), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_865), .B2(n_866), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_802), .B1(n_803), .B2(n_864), .Y(n_746) );
INVx1_ASAP7_75t_L g864 ( .A(n_747), .Y(n_864) );
OAI22xp5_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_749), .B1(n_766), .B2(n_799), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g765 ( .A(n_750), .Y(n_765) );
NOR2x1_ASAP7_75t_L g750 ( .A(n_751), .B(n_758), .Y(n_750) );
NAND4xp25_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .C(n_755), .D(n_757), .Y(n_751) );
NAND4xp25_ASAP7_75t_SL g758 ( .A(n_759), .B(n_761), .C(n_762), .D(n_763), .Y(n_758) );
INVx1_ASAP7_75t_L g846 ( .A(n_760), .Y(n_846) );
INVx2_ASAP7_75t_L g800 ( .A(n_767), .Y(n_800) );
AND2x4_ASAP7_75t_L g767 ( .A(n_768), .B(n_782), .Y(n_767) );
NOR2x1_ASAP7_75t_L g768 ( .A(n_769), .B(n_776), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_772), .Y(n_769) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
NOR2x1_ASAP7_75t_L g782 ( .A(n_783), .B(n_792), .Y(n_782) );
OAI222xp33_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_787), .B1(n_788), .B2(n_789), .C1(n_790), .C2(n_791), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
BUFx6f_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_797), .Y(n_792) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_820), .B1(n_821), .B2(n_863), .Y(n_803) );
INVx1_ASAP7_75t_L g863 ( .A(n_804), .Y(n_863) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
XNOR2x1_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_813), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_817), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_841), .Y(n_821) );
XOR2x2_ASAP7_75t_L g822 ( .A(n_823), .B(n_840), .Y(n_822) );
NAND2x1p5_ASAP7_75t_L g823 ( .A(n_824), .B(n_832), .Y(n_823) );
NOR2x1_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_826), .B(n_827), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
NOR2x1_ASAP7_75t_L g832 ( .A(n_833), .B(n_837), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_834), .B(n_836), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_844), .B(n_852), .Y(n_843) );
NOR2xp67_ASAP7_75t_L g844 ( .A(n_845), .B(n_849), .Y(n_844) );
OAI21xp5_ASAP7_75t_SL g845 ( .A1(n_846), .A2(n_847), .B(n_848), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NOR2x1_ASAP7_75t_L g852 ( .A(n_853), .B(n_858), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_854), .B(n_857), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_861), .Y(n_858) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OA22x2_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_893), .B2(n_894), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
NOR3x1_ASAP7_75t_SL g872 ( .A(n_873), .B(n_879), .C(n_882), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_877), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
NAND4xp25_ASAP7_75t_SL g882 ( .A(n_883), .B(n_886), .C(n_888), .D(n_891), .Y(n_882) );
INVx2_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
BUFx3_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_895), .A2(n_896), .B1(n_916), .B2(n_917), .Y(n_894) );
INVx2_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
XNOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
NAND2x1_ASAP7_75t_L g898 ( .A(n_899), .B(n_908), .Y(n_898) );
NOR2xp67_ASAP7_75t_L g899 ( .A(n_900), .B(n_904), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_905), .B(n_906), .Y(n_904) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_909), .B(n_912), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
INVx1_ASAP7_75t_SL g916 ( .A(n_917), .Y(n_916) );
XOR2x2_ASAP7_75t_L g917 ( .A(n_918), .B(n_934), .Y(n_917) );
NAND2xp5_ASAP7_75t_SL g918 ( .A(n_919), .B(n_927), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_923), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_926), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_928), .B(n_931), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_932), .B(n_933), .Y(n_931) );
INVx3_ASAP7_75t_SL g936 ( .A(n_937), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_938), .B(n_940), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_938), .B(n_941), .Y(n_983) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
OAI222xp33_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_960), .B1(n_962), .B2(n_979), .C1(n_981), .C2(n_984), .Y(n_945) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
NAND4xp75_ASAP7_75t_L g948 ( .A(n_949), .B(n_952), .C(n_955), .D(n_958), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_951), .Y(n_949) );
AND2x2_ASAP7_75t_L g952 ( .A(n_953), .B(n_954), .Y(n_952) );
AND2x2_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
INVx2_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx2_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g980 ( .A(n_967), .Y(n_980) );
NOR2x1_ASAP7_75t_L g967 ( .A(n_968), .B(n_973), .Y(n_967) );
NAND4xp25_ASAP7_75t_L g968 ( .A(n_969), .B(n_970), .C(n_971), .D(n_972), .Y(n_968) );
NAND4xp25_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .C(n_977), .D(n_978), .Y(n_973) );
INVx1_ASAP7_75t_SL g981 ( .A(n_982), .Y(n_981) );
CKINVDCx6p67_ASAP7_75t_R g982 ( .A(n_983), .Y(n_982) );
endmodule