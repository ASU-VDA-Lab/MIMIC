module fake_jpeg_10588_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_32),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_42),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_45),
.Y(n_52)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_29),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_28),
.B(n_20),
.Y(n_104)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_70),
.B1(n_34),
.B2(n_18),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_63),
.B1(n_43),
.B2(n_20),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_46),
.B1(n_27),
.B2(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_33),
.B1(n_27),
.B2(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_66),
.Y(n_79)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_27),
.B1(n_24),
.B2(n_16),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_77),
.A2(n_81),
.B1(n_86),
.B2(n_45),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_46),
.B1(n_45),
.B2(n_20),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_78),
.A2(n_83),
.B1(n_88),
.B2(n_105),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_64),
.B1(n_49),
.B2(n_54),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_95),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_92),
.Y(n_122)
);

NOR2xp67_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_1),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_28),
.B1(n_34),
.B2(n_24),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_18),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_4),
.C(n_5),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_96),
.Y(n_116)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_48),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_20),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_104),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_22),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_26),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_103),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_51),
.A2(n_19),
.B1(n_22),
.B2(n_3),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_1),
.B(n_4),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_68),
.B1(n_66),
.B2(n_19),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_107),
.A2(n_125),
.B1(n_135),
.B2(n_103),
.Y(n_161)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_115),
.B(n_74),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_121),
.A2(n_123),
.B1(n_92),
.B2(n_75),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_45),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_98),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_83),
.A2(n_45),
.B1(n_3),
.B2(n_4),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_126),
.A2(n_129),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_98),
.B(n_101),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_6),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_80),
.A2(n_45),
.B1(n_7),
.B2(n_8),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_149),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_73),
.C(n_72),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_153),
.C(n_136),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_145),
.B(n_151),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_78),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_156),
.C(n_118),
.Y(n_172)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_160),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_85),
.Y(n_143)
);

NAND2x1_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_136),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_93),
.B(n_80),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_126),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

OR2x4_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_95),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_152),
.B(n_154),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_96),
.B(n_94),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_119),
.B(n_74),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_157),
.B(n_158),
.Y(n_171)
);

OA21x2_ASAP7_75t_R g158 ( 
.A1(n_132),
.A2(n_8),
.B(n_9),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_161),
.B1(n_121),
.B2(n_132),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_116),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_115),
.B(n_8),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_133),
.C(n_130),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_159),
.B1(n_158),
.B2(n_112),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_182),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_166),
.A2(n_174),
.B(n_149),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_176),
.Y(n_190)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_175),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_178),
.C(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_118),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_117),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_184),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_127),
.C(n_111),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_156),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_183),
.C(n_152),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_112),
.C(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_184),
.B(n_179),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_188),
.A2(n_191),
.B(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_192),
.A2(n_198),
.B1(n_125),
.B2(n_157),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_139),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_201),
.C(n_181),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_167),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_195),
.B(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_202),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_144),
.Y(n_197)
);

AO21x2_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_150),
.B(n_153),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_161),
.B1(n_134),
.B2(n_131),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_190),
.C(n_193),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_206),
.C(n_212),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_172),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_205),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_176),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_198),
.A2(n_175),
.B1(n_107),
.B2(n_135),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_209),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_180),
.C(n_169),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_138),
.Y(n_213)
);

NOR4xp25_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_185),
.C(n_199),
.D(n_192),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_177),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_215),
.C(n_186),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_146),
.C(n_163),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_216),
.B(n_196),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_221),
.Y(n_235)
);

NOR3xp33_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_187),
.C(n_198),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_224),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_217),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_227),
.Y(n_230)
);

AOI31xp67_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_198),
.A3(n_202),
.B(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_191),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_210),
.B1(n_186),
.B2(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_236),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_206),
.B(n_110),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_237),
.C(n_233),
.Y(n_240)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_207),
.B(n_120),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_141),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_241),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_230),
.Y(n_246)
);

OAI221xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_229),
.B1(n_222),
.B2(n_223),
.C(n_220),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_223),
.B(n_220),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_230),
.B(n_123),
.C(n_116),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_243),
.B(n_246),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_244),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_9),
.B(n_12),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_204),
.B(n_75),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.C(n_10),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_251),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_12),
.C(n_13),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_14),
.Y(n_254)
);


endmodule