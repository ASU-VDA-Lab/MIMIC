module fake_jpeg_12624_n_184 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx6p67_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_23),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_43),
.A2(n_53),
.B1(n_0),
.B2(n_5),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_58),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_49),
.Y(n_66)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_26),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_13),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_21),
.C(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_8),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_30),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_17),
.B1(n_25),
.B2(n_13),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_89),
.B1(n_68),
.B2(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_34),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_29),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_37),
.B(n_24),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_51),
.B1(n_46),
.B2(n_38),
.Y(n_92)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_107),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_114),
.Y(n_117)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_45),
.B1(n_54),
.B2(n_71),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_108),
.B1(n_60),
.B2(n_84),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_74),
.B1(n_63),
.B2(n_78),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_110),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_66),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_113),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_88),
.B(n_79),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_130),
.B(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_82),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_85),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_124),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_85),
.Y(n_124)
);

NAND2xp33_ASAP7_75t_L g129 ( 
.A(n_94),
.B(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_100),
.B(n_106),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_77),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_90),
.C(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_84),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_106),
.A2(n_61),
.B1(n_62),
.B2(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_62),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_138),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_95),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_102),
.C(n_61),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_144),
.C(n_133),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_147),
.B(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

AND2x4_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVxp67_ASAP7_75t_SL g149 ( 
.A(n_146),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_132),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_150),
.A2(n_155),
.B(n_118),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_140),
.C(n_144),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_156),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_147),
.A2(n_118),
.B(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_131),
.B1(n_145),
.B2(n_118),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_141),
.A2(n_117),
.B(n_142),
.Y(n_155)
);

NOR4xp25_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_115),
.C(n_130),
.D(n_122),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_160),
.B(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_164),
.B1(n_166),
.B2(n_159),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_158),
.B(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_136),
.C(n_137),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_154),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_157),
.B1(n_154),
.B2(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_172),
.A2(n_163),
.B(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_134),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

AO21x2_ASAP7_75t_L g178 ( 
.A1(n_174),
.A2(n_172),
.B(n_167),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_179),
.B1(n_173),
.B2(n_166),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_170),
.B1(n_168),
.B2(n_166),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_181),
.B(n_178),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_128),
.B(n_120),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_126),
.B(n_182),
.Y(n_184)
);


endmodule