module real_aes_16569_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_889;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_502;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g117 ( .A(n_0), .B(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_1), .A2(n_533), .B1(n_534), .B2(n_536), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_1), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_2), .A2(n_35), .B1(n_160), .B2(n_252), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_3), .A2(n_12), .B1(n_565), .B2(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g118 ( .A(n_4), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_5), .Y(n_579) );
CKINVDCx5p33_ASAP7_75t_R g854 ( .A(n_6), .Y(n_854) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_7), .A2(n_13), .B1(n_566), .B2(n_602), .Y(n_601) );
XNOR2xp5_ASAP7_75t_L g534 ( .A(n_8), .B(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g121 ( .A(n_9), .Y(n_121) );
OR2x2_ASAP7_75t_L g139 ( .A(n_9), .B(n_31), .Y(n_139) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_10), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_11), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_14), .B(n_175), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_15), .A2(n_102), .B1(n_205), .B2(n_565), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_16), .A2(n_32), .B1(n_583), .B2(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_17), .B(n_175), .Y(n_580) );
OAI21x1_ASAP7_75t_L g155 ( .A1(n_18), .A2(n_48), .B(n_156), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_19), .B(n_256), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_20), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_20), .A2(n_95), .B1(n_638), .B2(n_873), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_21), .A2(n_39), .B1(n_212), .B2(n_227), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_22), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_23), .A2(n_45), .B1(n_227), .B2(n_565), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_24), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_25), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_26), .B(n_235), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_27), .Y(n_572) );
XNOR2x1_ASAP7_75t_L g535 ( .A(n_28), .B(n_40), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_29), .B(n_153), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_30), .Y(n_204) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_31), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_33), .A2(n_86), .B1(n_160), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_34), .A2(n_38), .B1(n_160), .B2(n_568), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_36), .A2(n_51), .B1(n_565), .B2(n_620), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_37), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_41), .B(n_175), .Y(n_223) );
INVx2_ASAP7_75t_L g134 ( .A(n_42), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_43), .B(n_208), .Y(n_250) );
INVx1_ASAP7_75t_L g113 ( .A(n_44), .Y(n_113) );
BUFx3_ASAP7_75t_L g137 ( .A(n_44), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_46), .B(n_194), .Y(n_258) );
XOR2x2_ASAP7_75t_L g142 ( .A(n_47), .B(n_143), .Y(n_142) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_47), .A2(n_875), .B1(n_876), .B2(n_879), .Y(n_874) );
INVx1_ASAP7_75t_L g879 ( .A(n_47), .Y(n_879) );
AND2x2_ASAP7_75t_L g286 ( .A(n_49), .B(n_194), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_50), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_52), .B(n_235), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g897 ( .A(n_53), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_54), .B(n_212), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_55), .A2(n_73), .B1(n_212), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_56), .A2(n_76), .B1(n_160), .B2(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_57), .B(n_316), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_58), .A2(n_164), .B(n_173), .C(n_279), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_59), .Y(n_891) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_60), .A2(n_99), .B1(n_565), .B2(n_566), .Y(n_564) );
INVx1_ASAP7_75t_L g156 ( .A(n_61), .Y(n_156) );
AND2x4_ASAP7_75t_L g178 ( .A(n_62), .B(n_179), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_63), .A2(n_64), .B1(n_227), .B2(n_239), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_65), .A2(n_83), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_65), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_66), .B(n_153), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_67), .B(n_194), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_68), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_69), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g179 ( .A(n_70), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_71), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_72), .B(n_153), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_74), .B(n_160), .Y(n_311) );
NAND3xp33_ASAP7_75t_L g251 ( .A(n_75), .B(n_208), .C(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_77), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g166 ( .A(n_78), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_79), .B(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_80), .B(n_175), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_81), .B(n_169), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_82), .A2(n_98), .B1(n_173), .B2(n_227), .Y(n_552) );
INVx1_ASAP7_75t_L g878 ( .A(n_83), .Y(n_878) );
CKINVDCx5p33_ASAP7_75t_R g623 ( .A(n_84), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_85), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_87), .A2(n_92), .B1(n_234), .B2(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_88), .B(n_175), .Y(n_207) );
NAND2xp33_ASAP7_75t_SL g192 ( .A(n_89), .B(n_163), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_90), .B(n_206), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_91), .B(n_153), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g605 ( .A(n_93), .Y(n_605) );
INVx1_ASAP7_75t_L g116 ( .A(n_94), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_94), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g873 ( .A(n_95), .Y(n_873) );
NAND2xp33_ASAP7_75t_L g584 ( .A(n_96), .B(n_175), .Y(n_584) );
NAND2xp33_ASAP7_75t_L g162 ( .A(n_97), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_100), .B(n_194), .Y(n_318) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_101), .B(n_163), .C(n_187), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_103), .B(n_160), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_104), .B(n_235), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_124), .B(n_896), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx11_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx10_ASAP7_75t_R g898 ( .A(n_109), .Y(n_898) );
OR2x6_ASAP7_75t_L g109 ( .A(n_110), .B(n_119), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2x1p5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
AND3x2_ASAP7_75t_L g885 ( .A(n_112), .B(n_115), .C(n_138), .Y(n_885) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g890 ( .A(n_113), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_117), .Y(n_114) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_115), .Y(n_864) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g130 ( .A(n_116), .Y(n_130) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
INVxp33_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_886), .Y(n_124) );
OAI211xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_140), .B(n_537), .C(n_865), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
NOR2xp67_ASAP7_75t_SL g127 ( .A(n_128), .B(n_131), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g859 ( .A(n_130), .B(n_860), .Y(n_859) );
NOR2x1_ASAP7_75t_R g863 ( .A(n_131), .B(n_864), .Y(n_863) );
INVx5_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x6_ASAP7_75t_SL g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_134), .B(n_858), .Y(n_857) );
INVx3_ASAP7_75t_L g868 ( .A(n_134), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2x1_ASAP7_75t_L g860 ( .A(n_137), .B(n_139), .Y(n_860) );
AND2x6_ASAP7_75t_SL g888 ( .A(n_138), .B(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B1(n_531), .B2(n_532), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVxp67_ASAP7_75t_SL g882 ( .A(n_143), .Y(n_882) );
OR2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_463), .Y(n_143) );
NAND4xp25_ASAP7_75t_L g144 ( .A(n_145), .B(n_338), .C(n_378), .D(n_427), .Y(n_144) );
NOR2xp67_ASAP7_75t_L g145 ( .A(n_146), .B(n_287), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_197), .B1(n_259), .B2(n_268), .Y(n_146) );
INVx1_ASAP7_75t_L g459 ( .A(n_147), .Y(n_459) );
INVx1_ASAP7_75t_SL g147 ( .A(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_148), .B(n_306), .Y(n_375) );
AND2x2_ASAP7_75t_L g406 ( .A(n_148), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_180), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g319 ( .A(n_149), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g330 ( .A(n_149), .Y(n_330) );
AND2x2_ASAP7_75t_L g505 ( .A(n_149), .B(n_373), .Y(n_505) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx2_ASAP7_75t_L g270 ( .A(n_150), .Y(n_270) );
AND2x2_ASAP7_75t_L g358 ( .A(n_150), .B(n_320), .Y(n_358) );
AND2x2_ASAP7_75t_L g402 ( .A(n_150), .B(n_307), .Y(n_402) );
OR2x2_ASAP7_75t_L g420 ( .A(n_150), .B(n_421), .Y(n_420) );
INVx4_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g324 ( .A(n_151), .B(n_307), .Y(n_324) );
BUFx2_ASAP7_75t_L g381 ( .A(n_151), .Y(n_381) );
OR2x2_ASAP7_75t_L g389 ( .A(n_151), .B(n_347), .Y(n_389) );
INVx1_ASAP7_75t_L g444 ( .A(n_151), .Y(n_444) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_157), .Y(n_151) );
INVx2_ASAP7_75t_L g592 ( .A(n_153), .Y(n_592) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x4_ASAP7_75t_SL g176 ( .A(n_154), .B(n_177), .Y(n_176) );
INVx1_ASAP7_75t_SL g183 ( .A(n_154), .Y(n_183) );
INVx2_ASAP7_75t_L g219 ( .A(n_154), .Y(n_219) );
BUFx3_ASAP7_75t_L g548 ( .A(n_154), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_154), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g576 ( .A(n_154), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_154), .B(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_154), .B(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_167), .B(n_176), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_164), .Y(n_158) );
OAI22xp33_ASAP7_75t_L g283 ( .A1(n_160), .A2(n_227), .B1(n_284), .B2(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g566 ( .A(n_160), .Y(n_566) );
INVx4_ASAP7_75t_L g568 ( .A(n_160), .Y(n_568) );
INVx1_ASAP7_75t_L g620 ( .A(n_160), .Y(n_620) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_161), .Y(n_163) );
INVx1_ASAP7_75t_L g173 ( .A(n_161), .Y(n_173) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_161), .Y(n_175) );
INVx1_ASAP7_75t_L g191 ( .A(n_161), .Y(n_191) );
INVx1_ASAP7_75t_L g206 ( .A(n_161), .Y(n_206) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_161), .Y(n_227) );
INVx1_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
INVx1_ASAP7_75t_L g239 ( .A(n_161), .Y(n_239) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_161), .Y(n_252) );
INVx2_ASAP7_75t_L g281 ( .A(n_161), .Y(n_281) );
INVx2_ASAP7_75t_L g212 ( .A(n_163), .Y(n_212) );
INVx1_ASAP7_75t_L g583 ( .A(n_163), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_164), .A2(n_190), .B(n_192), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_164), .A2(n_311), .B(n_312), .Y(n_310) );
BUFx4f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g171 ( .A(n_166), .Y(n_171) );
INVx1_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
BUFx8_ASAP7_75t_L g208 ( .A(n_166), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B1(n_172), .B2(n_174), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_169), .A2(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
BUFx3_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_175), .A2(n_186), .B(n_188), .Y(n_185) );
INVx1_ASAP7_75t_L g256 ( .A(n_175), .Y(n_256) );
INVx3_ASAP7_75t_L g565 ( .A(n_175), .Y(n_565) );
OAI21x1_ASAP7_75t_L g184 ( .A1(n_177), .A2(n_185), .B(n_189), .Y(n_184) );
OAI21x1_ASAP7_75t_L g202 ( .A1(n_177), .A2(n_203), .B(n_209), .Y(n_202) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_177), .A2(n_221), .B(n_224), .Y(n_220) );
OAI21x1_ASAP7_75t_L g248 ( .A1(n_177), .A2(n_249), .B(n_253), .Y(n_248) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_177), .A2(n_310), .B(n_313), .Y(n_309) );
BUFx10_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx10_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
INVx1_ASAP7_75t_L g555 ( .A(n_178), .Y(n_555) );
AND2x2_ASAP7_75t_L g271 ( .A(n_180), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g383 ( .A(n_180), .B(n_360), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_180), .B(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g421 ( .A(n_181), .Y(n_421) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_181), .Y(n_426) );
AND2x2_ASAP7_75t_L g443 ( .A(n_181), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g333 ( .A(n_182), .B(n_273), .Y(n_333) );
INVx1_ASAP7_75t_L g347 ( .A(n_182), .Y(n_347) );
OAI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_193), .Y(n_182) );
INVx1_ASAP7_75t_L g257 ( .A(n_187), .Y(n_257) );
INVx1_ASAP7_75t_L g553 ( .A(n_187), .Y(n_553) );
INVx1_ASAP7_75t_SL g569 ( .A(n_187), .Y(n_569) );
INVx1_ASAP7_75t_L g611 ( .A(n_191), .Y(n_611) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g201 ( .A(n_195), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_195), .B(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_195), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g242 ( .A(n_196), .Y(n_242) );
INVx2_ASAP7_75t_L g246 ( .A(n_196), .Y(n_246) );
NAND2x1_ASAP7_75t_L g197 ( .A(n_198), .B(n_214), .Y(n_197) );
AND2x4_ASAP7_75t_L g508 ( .A(n_198), .B(n_436), .Y(n_508) );
INVxp67_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
INVxp67_ASAP7_75t_SL g267 ( .A(n_199), .Y(n_267) );
BUFx3_ASAP7_75t_L g302 ( .A(n_199), .Y(n_302) );
INVx1_ASAP7_75t_L g368 ( .A(n_199), .Y(n_368) );
AND2x2_ASAP7_75t_L g371 ( .A(n_199), .B(n_217), .Y(n_371) );
AND2x2_ASAP7_75t_L g396 ( .A(n_199), .B(n_247), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_199), .Y(n_399) );
AND2x2_ASAP7_75t_L g431 ( .A(n_199), .B(n_296), .Y(n_431) );
INVx3_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OAI21x1_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_202), .B(n_213), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g297 ( .A1(n_201), .A2(n_202), .B(n_213), .Y(n_297) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_201), .A2(n_309), .B(n_318), .Y(n_308) );
OAI21xp33_ASAP7_75t_SL g336 ( .A1(n_201), .A2(n_309), .B(n_318), .Y(n_336) );
O2A1O1Ixp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .C(n_208), .Y(n_203) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_208), .A2(n_225), .B(n_226), .Y(n_224) );
INVx6_ASAP7_75t_L g237 ( .A(n_208), .Y(n_237) );
O2A1O1Ixp5_ASAP7_75t_L g578 ( .A1(n_208), .A2(n_568), .B(n_579), .C(n_580), .Y(n_578) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_229), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g340 ( .A(n_216), .B(n_326), .Y(n_340) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g366 ( .A(n_218), .B(n_353), .Y(n_366) );
AND2x2_ASAP7_75t_L g395 ( .A(n_218), .B(n_231), .Y(n_395) );
OR2x2_ASAP7_75t_L g491 ( .A(n_218), .B(n_231), .Y(n_491) );
OAI21x1_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_218) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_219), .A2(n_248), .B(n_258), .Y(n_247) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_219), .A2(n_220), .B(n_228), .Y(n_265) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_219), .A2(n_248), .B(n_258), .Y(n_296) );
INVx2_ASAP7_75t_L g234 ( .A(n_227), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_227), .A2(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g370 ( .A(n_229), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g519 ( .A(n_229), .Y(n_519) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_230), .Y(n_261) );
OR2x2_ASAP7_75t_L g453 ( .A(n_230), .B(n_263), .Y(n_453) );
INVx1_ASAP7_75t_L g475 ( .A(n_230), .Y(n_475) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_247), .Y(n_230) );
AND2x2_ASAP7_75t_L g291 ( .A(n_231), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g326 ( .A(n_231), .B(n_296), .Y(n_326) );
INVx1_ASAP7_75t_L g353 ( .A(n_231), .Y(n_353) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_231), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_231), .B(n_247), .Y(n_440) );
AO31x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_242), .A3(n_243), .B(n_244), .Y(n_231) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_237), .B1(n_238), .B2(n_240), .Y(n_232) );
INVx1_ASAP7_75t_L g602 ( .A(n_235), .Y(n_602) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g549 ( .A1(n_237), .A2(n_550), .B1(n_552), .B2(n_553), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_237), .A2(n_564), .B1(n_567), .B2(n_569), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_237), .A2(n_582), .B(n_584), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_237), .A2(n_240), .B1(n_590), .B2(n_591), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_237), .A2(n_569), .B1(n_601), .B2(n_603), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_237), .A2(n_240), .B1(n_610), .B2(n_612), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_237), .A2(n_240), .B1(n_619), .B2(n_621), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_237), .A2(n_240), .B1(n_635), .B2(n_636), .Y(n_634) );
INVx1_ASAP7_75t_L g613 ( .A(n_239), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_240), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g317 ( .A(n_241), .Y(n_317) );
INVx2_ASAP7_75t_L g275 ( .A(n_242), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_242), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_SL g604 ( .A(n_242), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g276 ( .A(n_243), .Y(n_276) );
AO31x2_ASAP7_75t_L g588 ( .A1(n_243), .A2(n_589), .A3(n_592), .B(n_593), .Y(n_588) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_243), .A2(n_562), .A3(n_600), .B(n_604), .Y(n_599) );
AO31x2_ASAP7_75t_L g608 ( .A1(n_243), .A2(n_548), .A3(n_609), .B(n_614), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
BUFx2_ASAP7_75t_L g562 ( .A(n_246), .Y(n_562) );
AND2x2_ASAP7_75t_L g377 ( .A(n_247), .B(n_297), .Y(n_377) );
INVx2_ASAP7_75t_L g316 ( .A(n_252), .Y(n_316) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_257), .Y(n_253) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR3x1_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .C(n_266), .Y(n_260) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_263), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g325 ( .A(n_263), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g376 ( .A(n_263), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g416 ( .A(n_263), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_263), .B(n_439), .Y(n_471) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_264), .B(n_352), .Y(n_412) );
AND2x2_ASAP7_75t_L g436 ( .A(n_264), .B(n_296), .Y(n_436) );
BUFx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g292 ( .A(n_265), .Y(n_292) );
BUFx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g447 ( .A(n_267), .B(n_326), .Y(n_447) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_270), .B(n_333), .Y(n_512) );
AND2x4_ASAP7_75t_L g504 ( .A(n_271), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_271), .B(n_324), .Y(n_518) );
INVx2_ASAP7_75t_L g320 ( .A(n_272), .Y(n_320) );
INVx1_ASAP7_75t_L g323 ( .A(n_272), .Y(n_323) );
INVx2_ASAP7_75t_L g408 ( .A(n_272), .Y(n_408) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g392 ( .A(n_273), .Y(n_392) );
AOI21x1_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_286), .Y(n_273) );
NOR2xp67_ASAP7_75t_SL g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g617 ( .A(n_275), .Y(n_617) );
INVx1_ASAP7_75t_L g570 ( .A(n_276), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_282), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx2_ASAP7_75t_SL g551 ( .A(n_281), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_327), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_303), .B1(n_321), .B2(n_325), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B(n_298), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g355 ( .A(n_291), .B(n_302), .Y(n_355) );
AND2x2_ASAP7_75t_L g515 ( .A(n_291), .B(n_396), .Y(n_515) );
BUFx2_ASAP7_75t_L g386 ( .A(n_292), .Y(n_386) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g385 ( .A(n_295), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g300 ( .A(n_296), .Y(n_300) );
INVx1_ASAP7_75t_L g352 ( .A(n_296), .Y(n_352) );
INVx1_ASAP7_75t_L g477 ( .A(n_297), .Y(n_477) );
AOI31xp33_ASAP7_75t_L g495 ( .A1(n_298), .A2(n_496), .A3(n_497), .B(n_498), .Y(n_495) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_299), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_300), .B(n_395), .Y(n_494) );
INVx2_ASAP7_75t_L g522 ( .A(n_300), .Y(n_522) );
INVxp67_ASAP7_75t_SL g337 ( .A(n_301), .Y(n_337) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g350 ( .A(n_302), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_302), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g480 ( .A(n_302), .B(n_440), .Y(n_480) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_319), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g391 ( .A(n_307), .B(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g360 ( .A(n_308), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_317), .Y(n_313) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_323), .Y(n_344) );
INVx1_ASAP7_75t_L g384 ( .A(n_323), .Y(n_384) );
INVx1_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
AND2x2_ASAP7_75t_L g425 ( .A(n_324), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g481 ( .A(n_324), .B(n_408), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_325), .A2(n_398), .B(n_400), .Y(n_397) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_337), .Y(n_327) );
NAND3x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .C(n_334), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g499 ( .A(n_330), .B(n_419), .Y(n_499) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2x1_ASAP7_75t_SL g452 ( .A(n_332), .B(n_364), .Y(n_452) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_373), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_334), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_334), .B(n_443), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_334), .B(n_443), .Y(n_516) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g419 ( .A(n_336), .B(n_392), .Y(n_419) );
AND2x2_ASAP7_75t_L g339 ( .A(n_337), .B(n_340), .Y(n_339) );
AOI221x1_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_341), .B1(n_348), .B2(n_357), .C(n_361), .Y(n_338) );
AOI32xp33_ASAP7_75t_L g520 ( .A1(n_340), .A2(n_521), .A3(n_526), .B1(n_527), .B2(n_529), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_345), .B(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g359 ( .A(n_347), .B(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_347), .Y(n_363) );
OR2x2_ASAP7_75t_L g476 ( .A(n_347), .B(n_477), .Y(n_476) );
NAND3xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_354), .C(n_356), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g398 ( .A(n_351), .B(n_399), .Y(n_398) );
AND2x4_ASAP7_75t_L g415 ( .A(n_351), .B(n_416), .Y(n_415) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_354), .A2(n_451), .B1(n_453), .B2(n_454), .Y(n_450) );
INVx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g528 ( .A(n_358), .Y(n_528) );
INVx2_ASAP7_75t_L g373 ( .A(n_360), .Y(n_373) );
OAI21xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B(n_369), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g497 ( .A(n_366), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_367), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B1(n_374), .B2(n_376), .Y(n_369) );
AND2x4_ASAP7_75t_L g466 ( .A(n_372), .B(n_381), .Y(n_466) );
INVx1_ASAP7_75t_L g525 ( .A(n_373), .Y(n_525) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g404 ( .A(n_377), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_377), .B(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_377), .B(n_405), .Y(n_496) );
AOI211x1_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_385), .B(n_387), .C(n_413), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR3x2_ASAP7_75t_L g488 ( .A(n_381), .B(n_383), .C(n_384), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_382), .A2(n_404), .B1(n_406), .B2(n_409), .Y(n_403) );
NOR2x1p5_ASAP7_75t_SL g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_383), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_521) );
INVx2_ASAP7_75t_L g405 ( .A(n_386), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_393), .B(n_397), .C(n_403), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_395), .B(n_399), .Y(n_410) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_395), .B(n_502), .Y(n_510) );
OAI32xp33_ASAP7_75t_L g485 ( .A1(n_396), .A2(n_441), .A3(n_486), .B1(n_488), .B2(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g502 ( .A(n_396), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_396), .B(n_416), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_399), .B(n_433), .Y(n_468) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g446 ( .A(n_405), .B(n_431), .Y(n_446) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g455 ( .A(n_408), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g423 ( .A(n_411), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B1(n_422), .B2(n_424), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g461 ( .A(n_418), .Y(n_461) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g442 ( .A(n_419), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_419), .B(n_426), .Y(n_530) );
INVx1_ASAP7_75t_SL g456 ( .A(n_420), .Y(n_456) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_450), .C(n_457), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_441), .B(n_445), .Y(n_428) );
NOR2xp33_ASAP7_75t_SL g429 ( .A(n_430), .B(n_434), .Y(n_429) );
INVxp67_ASAP7_75t_L g462 ( .A(n_430), .Y(n_462) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx1_ASAP7_75t_L g487 ( .A(n_432), .Y(n_487) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_437), .C(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g449 ( .A(n_443), .Y(n_449) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_447), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g458 ( .A(n_446), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_451), .A2(n_502), .B1(n_503), .B2(n_506), .C(n_507), .Y(n_501) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OAI32xp33_ASAP7_75t_L g457 ( .A1(n_454), .A2(n_458), .A3(n_459), .B1(n_460), .B2(n_462), .Y(n_457) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI221xp5_ASAP7_75t_L g469 ( .A1(n_460), .A2(n_470), .B1(n_471), .B2(n_472), .C(n_478), .Y(n_469) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_482), .C(n_500), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B(n_469), .Y(n_464) );
AOI211x1_ASAP7_75t_L g482 ( .A1(n_465), .A2(n_483), .B(n_485), .C(n_492), .Y(n_482) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVxp67_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2x1_ASAP7_75t_SL g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g484 ( .A(n_475), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AO21x1_ASAP7_75t_L g492 ( .A1(n_481), .A2(n_493), .B(n_495), .Y(n_492) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g526 ( .A(n_497), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_513), .Y(n_500) );
INVx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OAI21xp33_ASAP7_75t_SL g507 ( .A1(n_508), .A2(n_509), .B(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
NOR2xp67_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g523 ( .A(n_522), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_531), .A2(n_538), .B(n_850), .C(n_861), .Y(n_537) );
OAI21xp5_ASAP7_75t_L g850 ( .A1(n_531), .A2(n_851), .B(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g851 ( .A(n_540), .Y(n_851) );
NAND4xp75_ASAP7_75t_L g540 ( .A(n_541), .B(n_690), .C(n_766), .D(n_818), .Y(n_540) );
AND3x1_ASAP7_75t_L g541 ( .A(n_542), .B(n_663), .C(n_676), .Y(n_541) );
AOI221x1_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_595), .B1(n_624), .B2(n_628), .C(n_640), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_543), .A2(n_664), .B(n_666), .C(n_667), .Y(n_663) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_558), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g627 ( .A(n_547), .Y(n_627) );
BUFx2_ASAP7_75t_L g645 ( .A(n_547), .Y(n_645) );
OR2x2_ASAP7_75t_L g687 ( .A(n_547), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g694 ( .A(n_547), .B(n_561), .Y(n_694) );
AND2x4_ASAP7_75t_L g729 ( .A(n_547), .B(n_560), .Y(n_729) );
OR2x2_ASAP7_75t_L g772 ( .A(n_547), .B(n_588), .Y(n_772) );
AO31x2_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .A3(n_554), .B(n_556), .Y(n_547) );
AO31x2_ASAP7_75t_L g616 ( .A1(n_554), .A2(n_617), .A3(n_618), .B(n_622), .Y(n_616) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g585 ( .A(n_555), .Y(n_585) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_573), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_560), .B(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_560), .Y(n_659) );
INVx2_ASAP7_75t_L g686 ( .A(n_560), .Y(n_686) );
INVx3_ASAP7_75t_L g699 ( .A(n_560), .Y(n_699) );
AND2x2_ASAP7_75t_L g817 ( .A(n_560), .B(n_646), .Y(n_817) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g626 ( .A(n_561), .B(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g682 ( .A(n_561), .Y(n_682) );
AO31x2_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .A3(n_570), .B(n_571), .Y(n_561) );
AO31x2_ASAP7_75t_L g633 ( .A1(n_570), .A2(n_617), .A3(n_634), .B(n_637), .Y(n_633) );
INVxp67_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g702 ( .A(n_574), .Y(n_702) );
INVx1_ASAP7_75t_L g829 ( .A(n_574), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_587), .Y(n_574) );
AND2x2_ASAP7_75t_L g625 ( .A(n_575), .B(n_588), .Y(n_625) );
INVx1_ASAP7_75t_L g688 ( .A(n_575), .Y(n_688) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_586), .Y(n_575) );
OAI21x1_ASAP7_75t_L g647 ( .A1(n_576), .A2(n_577), .B(n_586), .Y(n_647) );
OAI21x1_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_585), .Y(n_577) );
INVx2_ASAP7_75t_L g643 ( .A(n_587), .Y(n_643) );
AND2x2_ASAP7_75t_L g695 ( .A(n_587), .B(n_646), .Y(n_695) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_588), .Y(n_717) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_597), .A2(n_689), .B1(n_693), .B2(n_696), .Y(n_692) );
AND2x4_ASAP7_75t_L g597 ( .A(n_598), .B(n_606), .Y(n_597) );
INVx1_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g630 ( .A(n_599), .B(n_608), .Y(n_630) );
AND2x2_ASAP7_75t_L g661 ( .A(n_599), .B(n_616), .Y(n_661) );
INVx4_ASAP7_75t_SL g672 ( .A(n_599), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_599), .B(n_706), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_599), .B(n_845), .Y(n_844) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g743 ( .A(n_607), .B(n_721), .Y(n_743) );
OR2x2_ASAP7_75t_L g776 ( .A(n_607), .B(n_758), .Y(n_776) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_616), .Y(n_607) );
INVx2_ASAP7_75t_L g650 ( .A(n_608), .Y(n_650) );
INVx1_ASAP7_75t_L g655 ( .A(n_608), .Y(n_655) );
AND2x2_ASAP7_75t_L g662 ( .A(n_608), .B(n_632), .Y(n_662) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_608), .Y(n_678) );
INVx1_ASAP7_75t_L g706 ( .A(n_608), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_608), .B(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g639 ( .A(n_616), .Y(n_639) );
AND2x4_ASAP7_75t_L g649 ( .A(n_616), .B(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g675 ( .A(n_616), .Y(n_675) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_616), .Y(n_752) );
INVx1_ASAP7_75t_L g845 ( .A(n_616), .Y(n_845) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_625), .B(n_698), .Y(n_765) );
AND2x2_ASAP7_75t_L g778 ( .A(n_625), .B(n_694), .Y(n_778) );
AND2x2_ASAP7_75t_L g848 ( .A(n_625), .B(n_699), .Y(n_848) );
AND2x4_ASAP7_75t_L g683 ( .A(n_627), .B(n_646), .Y(n_683) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
AND2x2_ASAP7_75t_L g750 ( .A(n_630), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g764 ( .A(n_630), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_630), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g666 ( .A(n_631), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_631), .B(n_704), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g760 ( .A1(n_631), .A2(n_761), .B(n_764), .C(n_765), .Y(n_760) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_639), .Y(n_631) );
AND2x2_ASAP7_75t_L g731 ( .A(n_632), .B(n_672), .Y(n_731) );
INVx3_ASAP7_75t_L g758 ( .A(n_632), .Y(n_758) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g653 ( .A(n_633), .Y(n_653) );
AND2x4_ASAP7_75t_L g679 ( .A(n_633), .B(n_639), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_639), .B(n_672), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_648), .B1(n_656), .B2(n_660), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g797 ( .A(n_642), .Y(n_797) );
AND2x4_ASAP7_75t_L g708 ( .A(n_643), .B(n_688), .Y(n_708) );
INVx1_ASAP7_75t_L g728 ( .A(n_643), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_645), .A2(n_701), .B1(n_711), .B2(n_713), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_645), .B(n_702), .Y(n_759) );
NAND2x1_ASAP7_75t_L g816 ( .A(n_645), .B(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g831 ( .A(n_645), .Y(n_831) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g770 ( .A(n_647), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g689 ( .A(n_649), .B(n_671), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_649), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g730 ( .A(n_649), .B(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_649), .Y(n_804) );
NAND2x1p5_ASAP7_75t_L g811 ( .A(n_649), .B(n_712), .Y(n_811) );
AND2x4_ASAP7_75t_L g834 ( .A(n_649), .B(n_762), .Y(n_834) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx3_ASAP7_75t_L g712 ( .A(n_652), .Y(n_712) );
AND2x2_ASAP7_75t_L g724 ( .A(n_652), .B(n_717), .Y(n_724) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g674 ( .A(n_653), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g722 ( .A(n_653), .Y(n_722) );
INVx1_ASAP7_75t_L g665 ( .A(n_654), .Y(n_665) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g822 ( .A(n_655), .B(n_672), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g748 ( .A(n_657), .B(n_729), .Y(n_748) );
INVx2_ASAP7_75t_L g789 ( .A(n_657), .Y(n_789) );
AND2x4_ASAP7_75t_L g790 ( .A(n_657), .B(n_683), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_658), .B(n_708), .Y(n_838) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_661), .B(n_721), .Y(n_720) );
AND2x4_ASAP7_75t_L g733 ( .A(n_661), .B(n_678), .Y(n_733) );
INVx1_ASAP7_75t_L g825 ( .A(n_661), .Y(n_825) );
AND2x2_ASAP7_75t_L g824 ( .A(n_662), .B(n_751), .Y(n_824) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g795 ( .A1(n_666), .A2(n_796), .B1(n_798), .B2(n_800), .Y(n_795) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_670), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g704 ( .A(n_672), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g740 ( .A(n_672), .Y(n_740) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_672), .Y(n_746) );
INVx2_ASAP7_75t_L g763 ( .A(n_672), .Y(n_763) );
OR2x2_ASAP7_75t_L g784 ( .A(n_672), .B(n_747), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_672), .B(n_742), .Y(n_794) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OR2x2_ASAP7_75t_L g761 ( .A(n_674), .B(n_762), .Y(n_761) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_674), .Y(n_815) );
INVx1_ASAP7_75t_L g742 ( .A(n_675), .Y(n_742) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_680), .B(n_684), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_678), .B(n_679), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_679), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g747 ( .A(n_679), .Y(n_747) );
AND2x2_ASAP7_75t_L g821 ( .A(n_679), .B(n_822), .Y(n_821) );
AOI211x1_ASAP7_75t_SL g749 ( .A1(n_680), .A2(n_750), .B(n_753), .C(n_760), .Y(n_749) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x4_ASAP7_75t_L g806 ( .A(n_682), .B(n_683), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_683), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g799 ( .A(n_683), .Y(n_799) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_689), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g714 ( .A(n_686), .Y(n_714) );
NOR2x1p5_ASAP7_75t_L g771 ( .A(n_686), .B(n_772), .Y(n_771) );
NOR2x1_ASAP7_75t_L g715 ( .A(n_687), .B(n_716), .Y(n_715) );
NOR2xp67_ASAP7_75t_SL g788 ( .A(n_687), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g849 ( .A(n_689), .B(n_757), .Y(n_849) );
NOR2x1_ASAP7_75t_L g690 ( .A(n_691), .B(n_734), .Y(n_690) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_700), .C(n_718), .Y(n_691) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_694), .Y(n_725) );
AND2x2_ASAP7_75t_L g732 ( .A(n_694), .B(n_728), .Y(n_732) );
AND2x4_ASAP7_75t_SL g846 ( .A(n_694), .B(n_708), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_695), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_697), .A2(n_739), .B1(n_811), .B2(n_812), .Y(n_810) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AND2x4_ASAP7_75t_L g828 ( .A(n_699), .B(n_829), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B1(n_707), .B2(n_709), .Y(n_701) );
NAND2x1_ASAP7_75t_L g777 ( .A(n_704), .B(n_757), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g787 ( .A(n_704), .B(n_751), .Y(n_787) );
INVx1_ASAP7_75t_L g814 ( .A(n_704), .Y(n_814) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_707), .A2(n_833), .B(n_836), .Y(n_832) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_708), .A2(n_720), .B(n_723), .Y(n_719) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g793 ( .A(n_712), .Y(n_793) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g737 ( .A(n_715), .Y(n_737) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AOI222xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_725), .B1(n_726), .B2(n_730), .C1(n_732), .C2(n_733), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g753 ( .A1(n_720), .A2(n_754), .B(n_759), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_721), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g835 ( .A(n_721), .Y(n_835) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g841 ( .A(n_722), .Y(n_841) );
AND2x2_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
AND2x2_ASAP7_75t_L g805 ( .A(n_727), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OR2x2_ASAP7_75t_L g798 ( .A(n_728), .B(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_749), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_738), .B1(n_744), .B2(n_748), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_743), .Y(n_738) );
OR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
INVx1_ASAP7_75t_L g755 ( .A(n_741), .Y(n_755) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx4_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g783 ( .A(n_758), .B(n_775), .Y(n_783) );
OR2x2_ASAP7_75t_L g843 ( .A(n_758), .B(n_844), .Y(n_843) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND5xp2_ASAP7_75t_L g819 ( .A(n_764), .B(n_811), .C(n_820), .D(n_823), .E(n_825), .Y(n_819) );
NOR2x1_ASAP7_75t_L g766 ( .A(n_767), .B(n_802), .Y(n_766) );
NAND2xp67_ASAP7_75t_SL g767 ( .A(n_768), .B(n_785), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_773), .B1(n_778), .B2(n_779), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
NAND3xp33_ASAP7_75t_SL g773 ( .A(n_774), .B(n_776), .C(n_777), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_L g808 ( .A(n_777), .Y(n_808) );
NAND3xp33_ASAP7_75t_SL g779 ( .A(n_780), .B(n_783), .C(n_784), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g801 ( .A(n_782), .Y(n_801) );
O2A1O1Ixp33_ASAP7_75t_SL g813 ( .A1(n_783), .A2(n_814), .B(n_815), .C(n_816), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .B1(n_790), .B2(n_791), .C(n_795), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_792), .B(n_840), .Y(n_839) );
OR2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx1_ASAP7_75t_L g809 ( .A(n_796), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_807), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g812 ( .A(n_806), .Y(n_812) );
AOI211xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_809), .B(n_810), .C(n_813), .Y(n_807) );
AOI211x1_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_826), .B(n_832), .C(n_847), .Y(n_818) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2x1p5_ASAP7_75t_L g827 ( .A(n_828), .B(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
NAND2x1_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_837), .A2(n_839), .B1(n_842), .B2(n_846), .Y(n_836) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AND2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g861 ( .A(n_852), .B(n_862), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
INVx5_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
BUFx10_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_869), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx8_ASAP7_75t_SL g867 ( .A(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_870), .B(n_892), .Y(n_869) );
AOI31xp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_882), .A3(n_883), .B(n_886), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_871), .B(n_894), .Y(n_893) );
AO22x1_ASAP7_75t_L g871 ( .A1(n_872), .A2(n_874), .B1(n_880), .B2(n_881), .Y(n_871) );
CKINVDCx5p33_ASAP7_75t_R g880 ( .A(n_872), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_874), .Y(n_881) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g895 ( .A(n_882), .Y(n_895) );
INVx1_ASAP7_75t_L g894 ( .A(n_883), .Y(n_894) );
BUFx2_ASAP7_75t_SL g883 ( .A(n_884), .Y(n_883) );
INVx4_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NOR2xp33_ASAP7_75t_SL g886 ( .A(n_887), .B(n_891), .Y(n_886) );
INVx5_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_895), .Y(n_892) );
NOR2xp33_ASAP7_75t_R g896 ( .A(n_897), .B(n_898), .Y(n_896) );
endmodule