module fake_jpeg_16875_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_40),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_15),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_23),
.B(n_26),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_21),
.B(n_23),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_41),
.A2(n_28),
.B(n_18),
.C(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_22),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_31),
.A2(n_16),
.B1(n_27),
.B2(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_57),
.B1(n_39),
.B2(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_30),
.B1(n_20),
.B2(n_27),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_35),
.B(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_54),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_20),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_27),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_31),
.A2(n_16),
.B1(n_30),
.B2(n_21),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_33),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_48),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_34),
.B(n_32),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_69),
.B(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_28),
.Y(n_93)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_50),
.Y(n_84)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_57),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_35),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_97),
.B(n_101),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_89),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_39),
.B1(n_51),
.B2(n_41),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_39),
.B1(n_56),
.B2(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_92),
.B1(n_80),
.B2(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_66),
.A2(n_56),
.B1(n_38),
.B2(n_59),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_95),
.B(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_18),
.B(n_38),
.C(n_29),
.D(n_25),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_78),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_65),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_25),
.B1(n_29),
.B2(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_102),
.B1(n_92),
.B2(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_111),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_95),
.C(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_71),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_114),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_24),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_64),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_97),
.Y(n_135)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_118),
.A2(n_100),
.B1(n_102),
.B2(n_84),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_122),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_59),
.C(n_55),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_49),
.C(n_2),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_115),
.B(n_118),
.C(n_85),
.D(n_114),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_123),
.B(n_141),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_105),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_135),
.Y(n_143)
);

OAI322xp33_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_103),
.A3(n_105),
.B1(n_111),
.B2(n_120),
.C1(n_122),
.C2(n_117),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_89),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_136),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_85),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

A2O1A1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_118),
.A2(n_85),
.B(n_91),
.C(n_97),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_72),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_35),
.C(n_38),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_106),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_68),
.B1(n_29),
.B2(n_25),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_49),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_168)
);

OAI322xp33_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_127),
.A3(n_132),
.B1(n_126),
.B2(n_4),
.C1(n_5),
.C2(n_8),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_134),
.B(n_110),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_148),
.B(n_152),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_141),
.C(n_126),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_10),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_162),
.C(n_163),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_147),
.A2(n_123),
.B1(n_132),
.B2(n_131),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_14),
.C(n_13),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_132),
.C(n_10),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_1),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_145),
.A2(n_1),
.B(n_2),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

BUFx12f_ASAP7_75t_SL g165 ( 
.A(n_156),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_165),
.A2(n_142),
.B(n_4),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_180),
.Y(n_182)
);

NAND4xp25_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_157),
.C(n_147),
.D(n_149),
.Y(n_175)
);

NOR2xp67_ASAP7_75t_SL g187 ( 
.A(n_175),
.B(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_176),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_157),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_179),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_170),
.B(n_142),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_166),
.B1(n_164),
.B2(n_162),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_168),
.B1(n_160),
.B2(n_164),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_184),
.B(n_177),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_171),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_11),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_188),
.B(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_195),
.B(n_197),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_173),
.B(n_181),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_3),
.B(n_8),
.C(n_191),
.D(n_196),
.Y(n_202)
);

OAI21x1_ASAP7_75t_SL g199 ( 
.A1(n_190),
.A2(n_11),
.B(n_12),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_199),
.B(n_3),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_8),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_200),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_203),
.Y(n_206)
);


endmodule