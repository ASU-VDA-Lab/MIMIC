module real_aes_6979_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_733;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g579 ( .A1(n_0), .A2(n_157), .B(n_580), .C(n_583), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_1), .B(n_524), .Y(n_584) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_2), .B(n_91), .C(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g444 ( .A(n_2), .Y(n_444) );
INVx1_ASAP7_75t_L g191 ( .A(n_3), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_4), .B(n_149), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_5), .A2(n_493), .B(n_518), .Y(n_517) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_6), .A2(n_134), .B(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_7), .A2(n_35), .B1(n_143), .B2(n_221), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_8), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_9), .B(n_134), .Y(n_160) );
AND2x6_ASAP7_75t_L g158 ( .A(n_10), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_11), .A2(n_158), .B(n_483), .C(n_485), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_108), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_12), .B(n_36), .Y(n_445) );
INVx1_ASAP7_75t_L g139 ( .A(n_13), .Y(n_139) );
INVx1_ASAP7_75t_L g184 ( .A(n_14), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_15), .B(n_147), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_16), .B(n_149), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_17), .B(n_135), .Y(n_196) );
AO32x2_ASAP7_75t_L g218 ( .A1(n_18), .A2(n_134), .A3(n_164), .B1(n_175), .B2(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_19), .B(n_143), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_20), .B(n_135), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_21), .A2(n_54), .B1(n_143), .B2(n_221), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g243 ( .A1(n_22), .A2(n_82), .B1(n_143), .B2(n_147), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_23), .B(n_143), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_24), .A2(n_175), .B(n_483), .C(n_544), .Y(n_543) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_25), .A2(n_175), .B(n_483), .C(n_512), .Y(n_511) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_26), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_27), .B(n_177), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_28), .A2(n_493), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_29), .B(n_177), .Y(n_215) );
INVx2_ASAP7_75t_L g145 ( .A(n_30), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_31), .A2(n_495), .B(n_503), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_32), .B(n_143), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_33), .B(n_177), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_34), .B(n_229), .Y(n_513) );
INVx1_ASAP7_75t_L g108 ( .A(n_36), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_37), .B(n_542), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_38), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_39), .A2(n_78), .B1(n_460), .B2(n_461), .Y(n_459) );
CKINVDCx16_ASAP7_75t_R g461 ( .A(n_39), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_40), .B(n_149), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_41), .B(n_493), .Y(n_510) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_42), .A2(n_79), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_42), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_43), .A2(n_495), .B(n_497), .C(n_503), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_44), .A2(n_459), .B1(n_462), .B2(n_463), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_44), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_45), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g581 ( .A(n_46), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_47), .A2(n_92), .B1(n_221), .B2(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g498 ( .A(n_48), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_49), .B(n_143), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_50), .B(n_143), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_51), .B(n_121), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_51), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_52), .B(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_53), .B(n_155), .Y(n_154) );
AOI22xp33_ASAP7_75t_SL g200 ( .A1(n_55), .A2(n_59), .B1(n_143), .B2(n_147), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_56), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_57), .B(n_143), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_58), .B(n_143), .Y(n_226) );
INVx1_ASAP7_75t_L g159 ( .A(n_60), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_61), .B(n_493), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_62), .B(n_524), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_63), .A2(n_155), .B(n_187), .C(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_64), .B(n_143), .Y(n_192) );
INVx1_ASAP7_75t_L g138 ( .A(n_65), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_66), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_67), .B(n_149), .Y(n_534) );
AO32x2_ASAP7_75t_L g239 ( .A1(n_68), .A2(n_134), .A3(n_175), .B1(n_240), .B2(n_244), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_69), .B(n_150), .Y(n_486) );
INVx1_ASAP7_75t_L g170 ( .A(n_70), .Y(n_170) );
INVx1_ASAP7_75t_L g210 ( .A(n_71), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g578 ( .A(n_72), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_73), .B(n_500), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g555 ( .A1(n_74), .A2(n_483), .B(n_503), .C(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_75), .B(n_147), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_76), .Y(n_519) );
INVx1_ASAP7_75t_L g112 ( .A(n_77), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_78), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_79), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_79), .A2(n_125), .B1(n_126), .B2(n_436), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_80), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_81), .B(n_499), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_83), .B(n_221), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_84), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_85), .B(n_147), .Y(n_214) );
INVx2_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_87), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_88), .A2(n_105), .B1(n_113), .B2(n_766), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_89), .B(n_174), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_90), .B(n_147), .Y(n_146) );
OR2x2_ASAP7_75t_L g441 ( .A(n_91), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g469 ( .A(n_91), .B(n_443), .Y(n_469) );
INVx2_ASAP7_75t_L g757 ( .A(n_91), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_93), .A2(n_103), .B1(n_147), .B2(n_148), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_94), .B(n_493), .Y(n_530) );
INVx1_ASAP7_75t_L g533 ( .A(n_95), .Y(n_533) );
INVxp67_ASAP7_75t_L g522 ( .A(n_96), .Y(n_522) );
AOI222xp33_ASAP7_75t_SL g457 ( .A1(n_97), .A2(n_458), .B1(n_464), .B2(n_758), .C1(n_759), .C2(n_763), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_98), .B(n_147), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_99), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g479 ( .A(n_100), .Y(n_479) );
INVx1_ASAP7_75t_L g557 ( .A(n_101), .Y(n_557) );
AND2x2_ASAP7_75t_L g505 ( .A(n_102), .B(n_177), .Y(n_505) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g767 ( .A(n_106), .Y(n_767) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AOI22x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_118), .B1(n_454), .B2(n_457), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g456 ( .A(n_117), .Y(n_456) );
AOI211xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_446), .B(n_447), .C(n_451), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_437), .C(n_440), .Y(n_119) );
INVxp67_ASAP7_75t_L g448 ( .A(n_120), .Y(n_448) );
INVx1_ASAP7_75t_L g439 ( .A(n_121), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_436), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g436 ( .A(n_126), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g126 ( .A(n_127), .B(n_360), .Y(n_126) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_128), .B(n_318), .Y(n_127) );
NOR4xp25_ASAP7_75t_L g128 ( .A(n_129), .B(n_258), .C(n_294), .D(n_308), .Y(n_128) );
OAI221xp5_ASAP7_75t_SL g129 ( .A1(n_130), .A2(n_202), .B1(n_234), .B2(n_245), .C(n_249), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_130), .B(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_178), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_161), .Y(n_132) );
AND2x2_ASAP7_75t_L g255 ( .A(n_133), .B(n_162), .Y(n_255) );
INVx3_ASAP7_75t_L g263 ( .A(n_133), .Y(n_263) );
AND2x2_ASAP7_75t_L g317 ( .A(n_133), .B(n_181), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_133), .B(n_180), .Y(n_353) );
AND2x2_ASAP7_75t_L g411 ( .A(n_133), .B(n_273), .Y(n_411) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_140), .B(n_160), .Y(n_133) );
INVx4_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_134), .A2(n_510), .B(n_511), .Y(n_509) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_134), .Y(n_516) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g164 ( .A(n_135), .Y(n_164) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g177 ( .A(n_136), .B(n_137), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_152), .B(n_158), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_149), .Y(n_141) );
INVx3_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_143), .Y(n_559) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g221 ( .A(n_144), .Y(n_221) );
BUFx3_ASAP7_75t_L g242 ( .A(n_144), .Y(n_242) );
AND2x6_ASAP7_75t_L g483 ( .A(n_144), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx2_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_149), .A2(n_167), .B(n_168), .Y(n_166) );
O2A1O1Ixp5_ASAP7_75t_SL g208 ( .A1(n_149), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g521 ( .A(n_149), .B(n_522), .Y(n_521) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g240 ( .A1(n_150), .A2(n_174), .B1(n_241), .B2(n_243), .Y(n_240) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_151), .Y(n_189) );
INVx1_ASAP7_75t_L g229 ( .A(n_151), .Y(n_229) );
AND2x2_ASAP7_75t_L g481 ( .A(n_151), .B(n_156), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_151), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .Y(n_152) );
INVx2_ASAP7_75t_L g171 ( .A(n_155), .Y(n_171) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_157), .A2(n_171), .B(n_191), .C(n_192), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_157), .A2(n_174), .B1(n_199), .B2(n_200), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_157), .A2(n_174), .B1(n_220), .B2(n_222), .Y(n_219) );
BUFx3_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g182 ( .A1(n_158), .A2(n_183), .B(n_190), .Y(n_182) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_158), .A2(n_208), .B(n_212), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_158), .A2(n_225), .B(n_230), .Y(n_224) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_158), .B(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g493 ( .A(n_158), .B(n_481), .Y(n_493) );
INVx4_ASAP7_75t_SL g504 ( .A(n_158), .Y(n_504) );
AND2x2_ASAP7_75t_L g246 ( .A(n_161), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g260 ( .A(n_161), .B(n_181), .Y(n_260) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_162), .B(n_181), .Y(n_275) );
AND2x2_ASAP7_75t_L g287 ( .A(n_162), .B(n_263), .Y(n_287) );
OR2x2_ASAP7_75t_L g289 ( .A(n_162), .B(n_247), .Y(n_289) );
AND2x2_ASAP7_75t_L g324 ( .A(n_162), .B(n_247), .Y(n_324) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_162), .Y(n_369) );
INVx1_ASAP7_75t_L g377 ( .A(n_162), .Y(n_377) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_176), .Y(n_162) );
OA21x2_ASAP7_75t_L g181 ( .A1(n_163), .A2(n_182), .B(n_193), .Y(n_181) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_164), .B(n_489), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_175), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .C(n_173), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_171), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_173), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx4_ASAP7_75t_L g582 ( .A(n_174), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g197 ( .A(n_175), .B(n_198), .C(n_201), .Y(n_197) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_177), .A2(n_207), .B(n_215), .Y(n_206) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_177), .A2(n_224), .B(n_233), .Y(n_223) );
INVx2_ASAP7_75t_L g244 ( .A(n_177), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_177), .A2(n_492), .B(n_494), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_177), .A2(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g550 ( .A(n_177), .Y(n_550) );
OAI221xp5_ASAP7_75t_L g294 ( .A1(n_178), .A2(n_295), .B1(n_299), .B2(n_303), .C(n_304), .Y(n_294) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g254 ( .A(n_179), .B(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_194), .Y(n_179) );
INVx2_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
AND2x2_ASAP7_75t_L g306 ( .A(n_180), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g325 ( .A(n_180), .B(n_263), .Y(n_325) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g388 ( .A(n_181), .B(n_263), .Y(n_388) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .C(n_187), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_185), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_185), .A2(n_513), .B(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_187), .A2(n_557), .B(n_558), .C(n_559), .Y(n_556) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_188), .A2(n_213), .B(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g500 ( .A(n_189), .Y(n_500) );
AND2x2_ASAP7_75t_L g310 ( .A(n_194), .B(n_255), .Y(n_310) );
OAI322xp33_ASAP7_75t_L g378 ( .A1(n_194), .A2(n_334), .A3(n_379), .B1(n_381), .B2(n_384), .C1(n_386), .C2(n_390), .Y(n_378) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_195), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g274 ( .A(n_195), .Y(n_274) );
AND2x2_ASAP7_75t_L g383 ( .A(n_195), .B(n_263), .Y(n_383) );
AND2x2_ASAP7_75t_L g415 ( .A(n_195), .B(n_287), .Y(n_415) );
OR2x2_ASAP7_75t_L g418 ( .A(n_195), .B(n_419), .Y(n_418) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_197), .Y(n_195) );
INVx1_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
AO21x1_ASAP7_75t_L g247 ( .A1(n_198), .A2(n_201), .B(n_248), .Y(n_247) );
AO21x2_ASAP7_75t_L g477 ( .A1(n_201), .A2(n_478), .B(n_488), .Y(n_477) );
INVx3_ASAP7_75t_L g524 ( .A(n_201), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_201), .B(n_536), .Y(n_535) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_201), .A2(n_554), .B(n_561), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_201), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_216), .Y(n_203) );
INVx1_ASAP7_75t_L g431 ( .A(n_204), .Y(n_431) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g236 ( .A(n_205), .B(n_223), .Y(n_236) );
INVx2_ASAP7_75t_L g271 ( .A(n_205), .Y(n_271) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g293 ( .A(n_206), .Y(n_293) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_206), .Y(n_301) );
OR2x2_ASAP7_75t_L g425 ( .A(n_206), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g250 ( .A(n_216), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g290 ( .A(n_216), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g342 ( .A(n_216), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
AND2x2_ASAP7_75t_L g237 ( .A(n_217), .B(n_238), .Y(n_237) );
NOR2xp67_ASAP7_75t_L g297 ( .A(n_217), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g351 ( .A(n_217), .B(n_239), .Y(n_351) );
OR2x2_ASAP7_75t_L g359 ( .A(n_217), .B(n_293), .Y(n_359) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx2_ASAP7_75t_L g268 ( .A(n_218), .Y(n_268) );
AND2x2_ASAP7_75t_L g278 ( .A(n_218), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g302 ( .A(n_218), .B(n_223), .Y(n_302) );
AND2x2_ASAP7_75t_L g366 ( .A(n_218), .B(n_239), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_223), .B(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_223), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g279 ( .A(n_223), .Y(n_279) );
INVx1_ASAP7_75t_L g284 ( .A(n_223), .Y(n_284) );
AND2x2_ASAP7_75t_L g296 ( .A(n_223), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_223), .Y(n_374) );
INVx1_ASAP7_75t_L g426 ( .A(n_223), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g403 ( .A(n_235), .B(n_312), .Y(n_403) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g330 ( .A(n_237), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g429 ( .A(n_237), .B(n_364), .Y(n_429) );
INVx1_ASAP7_75t_L g251 ( .A(n_238), .Y(n_251) );
AND2x2_ASAP7_75t_L g277 ( .A(n_238), .B(n_271), .Y(n_277) );
BUFx2_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_239), .Y(n_257) );
INVx1_ASAP7_75t_L g267 ( .A(n_239), .Y(n_267) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_242), .Y(n_502) );
INVx2_ASAP7_75t_L g583 ( .A(n_242), .Y(n_583) );
INVx1_ASAP7_75t_L g547 ( .A(n_244), .Y(n_547) );
NOR2xp67_ASAP7_75t_L g405 ( .A(n_245), .B(n_252), .Y(n_405) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI32xp33_ASAP7_75t_L g249 ( .A1(n_246), .A2(n_250), .A3(n_252), .B1(n_254), .B2(n_256), .Y(n_249) );
AND2x2_ASAP7_75t_L g389 ( .A(n_246), .B(n_262), .Y(n_389) );
AND2x2_ASAP7_75t_L g427 ( .A(n_246), .B(n_325), .Y(n_427) );
INVx1_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_251), .B(n_313), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_252), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_252), .B(n_255), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_252), .B(n_324), .Y(n_406) );
OR2x2_ASAP7_75t_L g420 ( .A(n_252), .B(n_289), .Y(n_420) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g347 ( .A(n_253), .B(n_255), .Y(n_347) );
OR2x2_ASAP7_75t_L g356 ( .A(n_253), .B(n_343), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_255), .B(n_306), .Y(n_328) );
INVx2_ASAP7_75t_L g343 ( .A(n_257), .Y(n_343) );
OR2x2_ASAP7_75t_L g358 ( .A(n_257), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_257), .B(n_374), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_257), .A2(n_350), .B(n_431), .C(n_432), .Y(n_430) );
OAI321xp33_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .A3(n_269), .B1(n_272), .B2(n_276), .C(n_280), .Y(n_258) );
INVx1_ASAP7_75t_L g371 ( .A(n_259), .Y(n_371) );
NAND2x1p5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g382 ( .A(n_260), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g334 ( .A(n_262), .Y(n_334) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_263), .B(n_377), .Y(n_394) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_264), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_407), .Y(n_401) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_268), .Y(n_265) );
AND2x2_ASAP7_75t_L g339 ( .A(n_266), .B(n_313), .Y(n_339) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_267), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g312 ( .A(n_268), .Y(n_312) );
A2O1A1Ixp33_ASAP7_75t_L g354 ( .A1(n_269), .A2(n_310), .B(n_355), .C(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g321 ( .A(n_271), .B(n_278), .Y(n_321) );
BUFx2_ASAP7_75t_L g331 ( .A(n_271), .Y(n_331) );
INVx1_ASAP7_75t_L g346 ( .A(n_271), .Y(n_346) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OR2x2_ASAP7_75t_L g352 ( .A(n_274), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g435 ( .A(n_274), .Y(n_435) );
INVx1_ASAP7_75t_L g428 ( .A(n_275), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_L g281 ( .A(n_277), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g385 ( .A(n_277), .B(n_302), .Y(n_385) );
INVx1_ASAP7_75t_L g314 ( .A(n_278), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_285), .B1(n_288), .B2(n_290), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_282), .B(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g350 ( .A(n_283), .B(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_SL g313 ( .A(n_284), .B(n_293), .Y(n_313) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g305 ( .A(n_287), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_292), .A2(n_410), .B1(n_412), .B2(n_413), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g298 ( .A(n_293), .Y(n_298) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_293), .Y(n_364) );
INVx1_ASAP7_75t_SL g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_296), .B(n_415), .Y(n_414) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_297), .A2(n_302), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_300), .B(n_310), .Y(n_407) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g376 ( .A(n_301), .Y(n_376) );
AND2x2_ASAP7_75t_L g335 ( .A(n_302), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g424 ( .A(n_302), .Y(n_424) );
INVx1_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
INVx1_ASAP7_75t_L g395 ( .A(n_306), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B1(n_314), .B2(n_315), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_312), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g380 ( .A(n_313), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_313), .B(n_351), .Y(n_417) );
OR2x2_ASAP7_75t_L g390 ( .A(n_314), .B(n_343), .Y(n_390) );
INVx1_ASAP7_75t_L g329 ( .A(n_315), .Y(n_329) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_317), .B(n_368), .Y(n_367) );
NOR3xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_337), .C(n_348), .Y(n_318) );
OAI211xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_322), .B(n_326), .C(n_332), .Y(n_319) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_321), .A2(n_392), .B1(n_396), .B2(n_399), .C(n_401), .Y(n_391) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g333 ( .A(n_324), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g387 ( .A(n_324), .B(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g372 ( .A1(n_325), .A2(n_373), .B(n_375), .C(n_377), .Y(n_372) );
INVx2_ASAP7_75t_L g419 ( .A(n_325), .Y(n_419) );
OAI21xp5_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_329), .B(n_330), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g398 ( .A(n_331), .B(n_351), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_335), .Y(n_332) );
OAI21xp5_ASAP7_75t_SL g337 ( .A1(n_338), .A2(n_340), .B(n_341), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI21xp5_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_344), .B(n_347), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_342), .B(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_347), .B(n_434), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B(n_354), .Y(n_348) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g375 ( .A(n_351), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND4x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_391), .C(n_408), .D(n_430), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_378), .Y(n_361) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_367), .B(n_370), .C(n_372), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_366), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_377), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g412 ( .A(n_387), .Y(n_412) );
INVx2_ASAP7_75t_SL g400 ( .A(n_388), .Y(n_400) );
OR2x2_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g413 ( .A(n_398), .Y(n_413) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_416), .Y(n_408) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
OAI221xp5_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_418), .B1(n_420), .B2(n_421), .C(n_422), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_427), .B1(n_428), .B2(n_429), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g449 ( .A(n_437), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_SL g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g450 ( .A(n_441), .Y(n_450) );
BUFx2_ASAP7_75t_L g452 ( .A(n_441), .Y(n_452) );
NOR2x2_ASAP7_75t_L g765 ( .A(n_442), .B(n_757), .Y(n_765) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g756 ( .A(n_443), .B(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
AOI211xp5_ASAP7_75t_L g447 ( .A1(n_446), .A2(n_448), .B(n_449), .C(n_450), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_451), .B(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g758 ( .A(n_458), .Y(n_758) );
INVx1_ASAP7_75t_L g462 ( .A(n_459), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g464 ( .A1(n_465), .A2(n_467), .B1(n_470), .B2(n_754), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g759 ( .A1(n_466), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_759) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g760 ( .A(n_468), .Y(n_760) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g761 ( .A(n_470), .Y(n_761) );
OR3x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_652), .C(n_717), .Y(n_470) );
NAND4xp25_ASAP7_75t_SL g471 ( .A(n_472), .B(n_593), .C(n_619), .D(n_642), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_525), .B1(n_563), .B2(n_570), .C(n_585), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_474), .A2(n_586), .B1(n_610), .B2(n_741), .Y(n_740) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_506), .Y(n_474) );
INVx1_ASAP7_75t_SL g646 ( .A(n_475), .Y(n_646) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
OR2x2_ASAP7_75t_L g568 ( .A(n_476), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g588 ( .A(n_476), .B(n_507), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_476), .B(n_515), .Y(n_601) );
AND2x2_ASAP7_75t_L g618 ( .A(n_476), .B(n_490), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_476), .B(n_566), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_476), .B(n_617), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_476), .B(n_506), .Y(n_739) );
AOI211xp5_ASAP7_75t_SL g750 ( .A1(n_476), .A2(n_656), .B(n_751), .C(n_752), .Y(n_750) );
INVx5_ASAP7_75t_SL g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_477), .B(n_507), .Y(n_622) );
AND2x2_ASAP7_75t_L g625 ( .A(n_477), .B(n_508), .Y(n_625) );
OR2x2_ASAP7_75t_L g670 ( .A(n_477), .B(n_507), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_477), .B(n_515), .Y(n_679) );
OAI21xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_482), .Y(n_478) );
INVx5_ASAP7_75t_L g496 ( .A(n_483), .Y(n_496) );
INVx5_ASAP7_75t_SL g569 ( .A(n_490), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_490), .B(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_490), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g673 ( .A(n_490), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g705 ( .A(n_490), .B(n_515), .Y(n_705) );
OR2x2_ASAP7_75t_L g711 ( .A(n_490), .B(n_601), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_490), .B(n_661), .Y(n_720) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_505), .Y(n_490) );
BUFx2_ASAP7_75t_L g542 ( .A(n_493), .Y(n_542) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_496), .A2(n_504), .B(n_519), .C(n_520), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_SL g577 ( .A1(n_496), .A2(n_504), .B(n_578), .C(n_579), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B(n_501), .C(n_502), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_499), .A2(n_502), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
AND2x2_ASAP7_75t_L g602 ( .A(n_507), .B(n_569), .Y(n_602) );
INVx1_ASAP7_75t_SL g615 ( .A(n_507), .Y(n_615) );
OR2x2_ASAP7_75t_L g650 ( .A(n_507), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g656 ( .A(n_507), .B(n_515), .Y(n_656) );
AND2x2_ASAP7_75t_L g714 ( .A(n_507), .B(n_566), .Y(n_714) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_508), .B(n_569), .Y(n_641) );
INVx3_ASAP7_75t_L g566 ( .A(n_515), .Y(n_566) );
OR2x2_ASAP7_75t_L g607 ( .A(n_515), .B(n_569), .Y(n_607) );
AND2x2_ASAP7_75t_L g617 ( .A(n_515), .B(n_615), .Y(n_617) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_515), .Y(n_665) );
AND2x2_ASAP7_75t_L g674 ( .A(n_515), .B(n_588), .Y(n_674) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_515) );
OA21x2_ASAP7_75t_L g575 ( .A1(n_524), .A2(n_576), .B(n_584), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_525), .A2(n_691), .B1(n_693), .B2(n_695), .C(n_698), .Y(n_690) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_537), .Y(n_526) );
AND2x2_ASAP7_75t_L g664 ( .A(n_527), .B(n_645), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_527), .B(n_723), .Y(n_727) );
OR2x2_ASAP7_75t_L g748 ( .A(n_527), .B(n_749), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_527), .B(n_753), .Y(n_752) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx5_ASAP7_75t_L g595 ( .A(n_528), .Y(n_595) );
AND2x2_ASAP7_75t_L g672 ( .A(n_528), .B(n_539), .Y(n_672) );
AND2x2_ASAP7_75t_L g733 ( .A(n_528), .B(n_612), .Y(n_733) );
AND2x2_ASAP7_75t_L g746 ( .A(n_528), .B(n_566), .Y(n_746) );
OR2x6_ASAP7_75t_L g528 ( .A(n_529), .B(n_535), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_551), .Y(n_537) );
AND2x4_ASAP7_75t_L g573 ( .A(n_538), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g591 ( .A(n_538), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g598 ( .A(n_538), .Y(n_598) );
AND2x2_ASAP7_75t_L g667 ( .A(n_538), .B(n_645), .Y(n_667) );
AND2x2_ASAP7_75t_L g677 ( .A(n_538), .B(n_595), .Y(n_677) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_538), .Y(n_685) );
AND2x2_ASAP7_75t_L g697 ( .A(n_538), .B(n_575), .Y(n_697) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_538), .B(n_629), .Y(n_701) );
AND2x2_ASAP7_75t_L g738 ( .A(n_538), .B(n_733), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_538), .B(n_612), .Y(n_749) );
OR2x2_ASAP7_75t_L g751 ( .A(n_538), .B(n_687), .Y(n_751) );
INVx5_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g637 ( .A(n_539), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g647 ( .A(n_539), .B(n_592), .Y(n_647) );
AND2x2_ASAP7_75t_L g659 ( .A(n_539), .B(n_575), .Y(n_659) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_539), .Y(n_689) );
AND2x4_ASAP7_75t_L g723 ( .A(n_539), .B(n_574), .Y(n_723) );
OR2x6_ASAP7_75t_L g539 ( .A(n_540), .B(n_548), .Y(n_539) );
AOI21xp5_ASAP7_75t_SL g540 ( .A1(n_541), .A2(n_543), .B(n_547), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
BUFx2_ASAP7_75t_L g572 ( .A(n_551), .Y(n_572) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g612 ( .A(n_552), .Y(n_612) );
AND2x2_ASAP7_75t_L g645 ( .A(n_552), .B(n_575), .Y(n_645) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g592 ( .A(n_553), .B(n_575), .Y(n_592) );
BUFx2_ASAP7_75t_L g638 ( .A(n_553), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_565), .B(n_646), .Y(n_725) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_566), .B(n_588), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_566), .B(n_569), .Y(n_627) );
AND2x2_ASAP7_75t_L g682 ( .A(n_566), .B(n_618), .Y(n_682) );
AOI221xp5_ASAP7_75t_SL g619 ( .A1(n_567), .A2(n_620), .B1(n_628), .B2(n_630), .C(n_634), .Y(n_619) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g614 ( .A(n_568), .B(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g655 ( .A(n_568), .B(n_656), .Y(n_655) );
OAI321xp33_ASAP7_75t_L g662 ( .A1(n_568), .A2(n_621), .A3(n_663), .B1(n_665), .B2(n_666), .C(n_668), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_569), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_572), .B(n_723), .Y(n_741) );
AND2x2_ASAP7_75t_L g628 ( .A(n_573), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_573), .B(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_574), .Y(n_604) );
AND2x2_ASAP7_75t_L g611 ( .A(n_574), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_574), .B(n_686), .Y(n_716) );
INVx1_ASAP7_75t_L g753 ( .A(n_574), .Y(n_753) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B(n_590), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
A2O1A1Ixp33_ASAP7_75t_L g745 ( .A1(n_587), .A2(n_697), .B(n_746), .C(n_747), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_588), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_588), .B(n_626), .Y(n_692) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g635 ( .A(n_592), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_592), .B(n_595), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_592), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_592), .B(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_596), .B1(n_608), .B2(n_613), .Y(n_593) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g609 ( .A(n_595), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g632 ( .A(n_595), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g644 ( .A(n_595), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_595), .B(n_638), .Y(n_680) );
OR2x2_ASAP7_75t_L g687 ( .A(n_595), .B(n_612), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_595), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g737 ( .A(n_595), .B(n_723), .Y(n_737) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .B1(n_603), .B2(n_605), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g643 ( .A(n_598), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_601), .A2(n_616), .B1(n_684), .B2(n_688), .Y(n_683) );
INVx1_ASAP7_75t_L g731 ( .A(n_602), .Y(n_731) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_606), .A2(n_643), .B1(n_646), .B2(n_647), .C(n_648), .Y(n_642) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g621 ( .A(n_607), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_611), .B(n_677), .Y(n_709) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_612), .Y(n_629) );
INVx1_ASAP7_75t_L g633 ( .A(n_612), .Y(n_633) );
NAND2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
INVx1_ASAP7_75t_L g651 ( .A(n_618), .Y(n_651) );
AND2x2_ASAP7_75t_L g660 ( .A(n_618), .B(n_661), .Y(n_660) );
NAND2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g704 ( .A(n_625), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_628), .A2(n_654), .B1(n_657), .B2(n_660), .C(n_662), .Y(n_653) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_632), .B(n_689), .Y(n_688) );
AOI21xp33_ASAP7_75t_SL g634 ( .A1(n_635), .A2(n_636), .B(n_639), .Y(n_634) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_639), .Y(n_736) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OR2x2_ASAP7_75t_L g678 ( .A(n_641), .B(n_679), .Y(n_678) );
INVx1_ASAP7_75t_SL g699 ( .A(n_644), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_644), .B(n_704), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_647), .B(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_671), .C(n_690), .D(n_703), .Y(n_652) );
INVx1_ASAP7_75t_SL g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g661 ( .A(n_656), .Y(n_661) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g694 ( .A(n_665), .B(n_670), .Y(n_694) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B(n_675), .C(n_683), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g742 ( .A1(n_673), .A2(n_715), .B(n_743), .C(n_750), .Y(n_742) );
INVx1_ASAP7_75t_SL g702 ( .A(n_674), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B1(n_680), .B2(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g706 ( .A(n_680), .Y(n_706) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_686), .B(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_686), .B(n_697), .Y(n_730) );
INVx2_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g707 ( .A(n_697), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_700), .B(n_702), .Y(n_698) );
INVxp33_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI322xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_706), .A3(n_707), .B1(n_708), .B2(n_710), .C1(n_712), .C2(n_715), .Y(n_703) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g717 ( .A(n_718), .B(n_735), .C(n_742), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_724), .B2(n_726), .C(n_728), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g734 ( .A(n_723), .Y(n_734) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_735) );
NAND2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVxp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g762 ( .A(n_755), .Y(n_762) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
endmodule