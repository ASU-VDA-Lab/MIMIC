module fake_jpeg_19305_n_144 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_144);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx4f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_1),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_36),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

HAxp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_1),
.CON(n_72),
.SN(n_72)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_77),
.B1(n_51),
.B2(n_57),
.Y(n_89)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_75),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_77),
.A2(n_58),
.B1(n_55),
.B2(n_68),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_69),
.B1(n_66),
.B2(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_72),
.B(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_90),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_74),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_88),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_56),
.B1(n_47),
.B2(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_3),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_62),
.B1(n_53),
.B2(n_63),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_66),
.B1(n_65),
.B2(n_64),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_87),
.B1(n_67),
.B2(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_49),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_26),
.B1(n_43),
.B2(n_40),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_118)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_3),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_111),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_4),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_117),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_99),
.B1(n_7),
.B2(n_13),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_12),
.B(n_14),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_27),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_15),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_128),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_114),
.A2(n_16),
.B1(n_18),
.B2(n_22),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_111),
.Y(n_133)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_131),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_124),
.B(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_124),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_133),
.B(n_123),
.C(n_132),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_108),
.B1(n_125),
.B2(n_115),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_138),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_139),
.A2(n_28),
.B(n_29),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_107),
.B1(n_110),
.B2(n_34),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_142),
.A2(n_30),
.B(n_32),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_37),
.Y(n_144)
);


endmodule