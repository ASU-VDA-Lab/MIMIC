module real_aes_4145_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_503;
wire n_635;
wire n_357;
wire n_287;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_892;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_397;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_928;
wire n_637;
wire n_653;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_946;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_949;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_0), .A2(n_222), .B1(n_390), .B2(n_391), .Y(n_441) );
AO22x2_ASAP7_75t_L g419 ( .A1(n_1), .A2(n_420), .B1(n_443), .B2(n_444), .Y(n_419) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_1), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_1), .A2(n_50), .B1(n_706), .B2(n_709), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_2), .A2(n_57), .B1(n_257), .B2(n_599), .Y(n_903) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_3), .Y(n_664) );
AND2x4_ASAP7_75t_L g679 ( .A(n_3), .B(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g689 ( .A(n_3), .B(n_237), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_4), .A2(n_187), .B1(n_257), .B2(n_282), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_5), .A2(n_89), .B1(n_390), .B2(n_391), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_6), .A2(n_212), .B1(n_292), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_7), .A2(n_10), .B1(n_384), .B2(n_385), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_8), .A2(n_13), .B1(n_506), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_9), .A2(n_200), .B1(n_474), .B2(n_506), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_11), .A2(n_108), .B1(n_643), .B2(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_12), .B(n_432), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_14), .A2(n_75), .B1(n_503), .B2(n_600), .Y(n_905) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_15), .A2(n_74), .B1(n_699), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_16), .A2(n_119), .B1(n_382), .B2(n_391), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_17), .A2(n_110), .B1(n_334), .B2(n_337), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_18), .A2(n_177), .B1(n_450), .B2(n_451), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_19), .Y(n_536) );
INVx1_ASAP7_75t_L g686 ( .A(n_20), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_21), .A2(n_192), .B1(n_466), .B2(n_468), .Y(n_465) );
INVx1_ASAP7_75t_L g493 ( .A(n_22), .Y(n_493) );
INVx1_ASAP7_75t_L g541 ( .A(n_23), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_24), .A2(n_100), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g578 ( .A(n_25), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_26), .A2(n_149), .B1(n_387), .B2(n_388), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_27), .A2(n_72), .B1(n_692), .B2(n_722), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_28), .A2(n_130), .B1(n_368), .B2(n_372), .Y(n_532) );
INVx1_ASAP7_75t_SL g755 ( .A(n_29), .Y(n_755) );
XNOR2x1_ASAP7_75t_L g485 ( .A(n_30), .B(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_31), .A2(n_157), .B1(n_646), .B2(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g898 ( .A(n_32), .Y(n_898) );
INVx1_ASAP7_75t_L g279 ( .A(n_33), .Y(n_279) );
INVxp67_ASAP7_75t_L g332 ( .A(n_33), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_33), .B(n_182), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_34), .A2(n_114), .B1(n_368), .B2(n_384), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_35), .A2(n_84), .B1(n_676), .B2(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_36), .B(n_453), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_37), .A2(n_95), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_38), .A2(n_116), .B1(n_473), .B2(n_649), .Y(n_648) );
XNOR2x1_ASAP7_75t_L g620 ( .A(n_39), .B(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_40), .A2(n_66), .B1(n_381), .B2(n_382), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g941 ( .A1(n_41), .A2(n_97), .B1(n_257), .B2(n_942), .Y(n_941) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_42), .B(n_263), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_43), .A2(n_215), .B1(n_314), .B2(n_506), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_44), .A2(n_80), .B1(n_301), .B2(n_304), .Y(n_300) );
AOI21xp33_ASAP7_75t_SL g422 ( .A1(n_45), .A2(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g525 ( .A(n_46), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_47), .A2(n_96), .B1(n_320), .B2(n_928), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_48), .A2(n_229), .B1(n_371), .B2(n_372), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_49), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_51), .A2(n_150), .B1(n_342), .B2(n_346), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_52), .A2(n_205), .B1(n_369), .B2(n_371), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_53), .A2(n_248), .B1(n_688), .B2(n_723), .Y(n_743) );
BUFx2_ASAP7_75t_L g430 ( .A(n_54), .Y(n_430) );
INVxp67_ASAP7_75t_R g690 ( .A(n_55), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_56), .A2(n_94), .B1(n_384), .B2(n_385), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_58), .A2(n_183), .B1(n_384), .B2(n_385), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_59), .A2(n_236), .B1(n_302), .B2(n_471), .Y(n_564) );
INVx2_ASAP7_75t_L g662 ( .A(n_60), .Y(n_662) );
INVx1_ASAP7_75t_L g678 ( .A(n_61), .Y(n_678) );
AND2x4_ASAP7_75t_L g683 ( .A(n_61), .B(n_662), .Y(n_683) );
INVx1_ASAP7_75t_SL g700 ( .A(n_61), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_62), .A2(n_186), .B1(n_387), .B2(n_388), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_63), .A2(n_139), .B1(n_334), .B2(n_346), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_64), .A2(n_165), .B1(n_468), .B2(n_529), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_65), .A2(n_147), .B1(n_320), .B2(n_323), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_67), .B(n_613), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_68), .A2(n_153), .B1(n_323), .B2(n_930), .Y(n_929) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_69), .A2(n_173), .B1(n_699), .B2(n_713), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g603 ( .A1(n_70), .A2(n_226), .B1(n_257), .B2(n_282), .Y(n_603) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_71), .Y(n_263) );
XNOR2x2_ASAP7_75t_SL g561 ( .A(n_73), .B(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_76), .A2(n_184), .B1(n_387), .B2(n_388), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_77), .A2(n_162), .B1(n_308), .B2(n_314), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_78), .A2(n_243), .B1(n_385), .B2(n_390), .Y(n_410) );
INVx1_ASAP7_75t_L g514 ( .A(n_79), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g895 ( .A1(n_81), .A2(n_896), .B(n_897), .Y(n_895) );
INVx1_ASAP7_75t_L g926 ( .A(n_82), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_83), .A2(n_85), .B1(n_372), .B2(n_381), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g684 ( .A(n_86), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_87), .A2(n_142), .B1(n_676), .B2(n_774), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_88), .A2(n_199), .B1(n_552), .B2(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_90), .A2(n_136), .B1(n_450), .B2(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g264 ( .A(n_91), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_91), .B(n_181), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_92), .A2(n_888), .B1(n_906), .B2(n_907), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_92), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_93), .A2(n_230), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_98), .A2(n_195), .B1(n_368), .B2(n_369), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_99), .A2(n_137), .B1(n_346), .B2(n_456), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_101), .A2(n_217), .B1(n_523), .B2(n_582), .C(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g701 ( .A(n_102), .Y(n_701) );
XNOR2x1_ASAP7_75t_L g400 ( .A(n_103), .B(n_401), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_103), .A2(n_143), .B1(n_722), .B2(n_723), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_104), .A2(n_161), .B1(n_615), .B2(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g591 ( .A(n_105), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_106), .A2(n_190), .B1(n_282), .B2(n_602), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g439 ( .A1(n_107), .A2(n_241), .B1(n_381), .B2(n_382), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_109), .A2(n_123), .B1(n_624), .B2(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g585 ( .A(n_111), .Y(n_585) );
INVx1_ASAP7_75t_L g637 ( .A(n_112), .Y(n_637) );
INVx1_ASAP7_75t_L g425 ( .A(n_113), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_115), .A2(n_148), .B1(n_688), .B2(n_692), .Y(n_757) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_117), .A2(n_374), .B(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_118), .A2(n_140), .B1(n_297), .B2(n_503), .Y(n_936) );
INVx1_ASAP7_75t_L g408 ( .A(n_120), .Y(n_408) );
INVx1_ASAP7_75t_L g495 ( .A(n_121), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_122), .A2(n_167), .B1(n_508), .B2(n_545), .Y(n_544) );
XOR2x2_ASAP7_75t_L g519 ( .A(n_124), .B(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_125), .A2(n_210), .B1(n_372), .B2(n_437), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_126), .A2(n_128), .B1(n_450), .B2(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_127), .A2(n_320), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g573 ( .A(n_129), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_131), .A2(n_132), .B1(n_471), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g446 ( .A(n_133), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_133), .A2(n_219), .B1(n_706), .B2(n_709), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_134), .B(n_339), .Y(n_403) );
INVx1_ASAP7_75t_L g704 ( .A(n_135), .Y(n_704) );
INVx1_ASAP7_75t_L g702 ( .A(n_138), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_141), .A2(n_172), .B1(n_651), .B2(n_652), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_144), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g361 ( .A(n_145), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_146), .A2(n_194), .B1(n_302), .B2(n_501), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_151), .A2(n_218), .B1(n_257), .B2(n_470), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_152), .A2(n_171), .B1(n_627), .B2(n_629), .Y(n_626) );
OA22x2_ASAP7_75t_L g269 ( .A1(n_154), .A2(n_182), .B1(n_263), .B2(n_267), .Y(n_269) );
INVx1_ASAP7_75t_L g288 ( .A(n_154), .Y(n_288) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_155), .A2(n_632), .B(n_635), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_156), .A2(n_245), .B1(n_282), .B2(n_508), .Y(n_507) );
XOR2x2_ASAP7_75t_L g253 ( .A(n_158), .B(n_254), .Y(n_253) );
AOI221x1_ASAP7_75t_L g922 ( .A1(n_159), .A2(n_207), .B1(n_634), .B2(n_923), .C(n_925), .Y(n_922) );
INVx1_ASAP7_75t_L g640 ( .A(n_160), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_163), .A2(n_166), .B1(n_387), .B2(n_388), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_164), .A2(n_175), .B1(n_599), .B2(n_600), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_168), .A2(n_232), .B1(n_503), .B2(n_556), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_169), .A2(n_228), .B1(n_390), .B2(n_391), .Y(n_527) );
INVx1_ASAP7_75t_L g580 ( .A(n_170), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_174), .A2(n_204), .B1(n_369), .B2(n_371), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_176), .B(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_178), .B(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g434 ( .A(n_179), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_180), .A2(n_209), .B1(n_387), .B2(n_388), .Y(n_442) );
INVx1_ASAP7_75t_L g281 ( .A(n_181), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_181), .B(n_286), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g289 ( .A1(n_182), .A2(n_202), .B(n_290), .Y(n_289) );
CKINVDCx6p67_ASAP7_75t_R g681 ( .A(n_185), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_188), .A2(n_246), .B1(n_676), .B2(n_725), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_189), .A2(n_211), .B1(n_566), .B2(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g491 ( .A(n_191), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_193), .A2(n_227), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI221x1_ASAP7_75t_SL g538 ( .A1(n_196), .A2(n_197), .B1(n_320), .B2(n_539), .C(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g609 ( .A(n_198), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_201), .A2(n_242), .B1(n_522), .B2(n_523), .C(n_524), .Y(n_521) );
INVx1_ASAP7_75t_L g266 ( .A(n_202), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_202), .B(n_231), .Y(n_355) );
AOI21xp33_ASAP7_75t_L g607 ( .A1(n_203), .A2(n_320), .B(n_608), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g509 ( .A1(n_206), .A2(n_234), .B1(n_510), .B2(n_511), .C(n_513), .Y(n_509) );
INVx1_ASAP7_75t_L g756 ( .A(n_208), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_208), .A2(n_913), .B1(n_916), .B2(n_949), .Y(n_912) );
OAI21x1_ASAP7_75t_L g919 ( .A1(n_208), .A2(n_920), .B(n_943), .Y(n_919) );
INVx1_ASAP7_75t_L g459 ( .A(n_213), .Y(n_459) );
INVx1_ASAP7_75t_L g376 ( .A(n_214), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_216), .A2(n_233), .B1(n_473), .B2(n_474), .Y(n_554) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_220), .A2(n_374), .B(n_375), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_221), .A2(n_225), .B1(n_292), .B2(n_297), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_223), .A2(n_238), .B1(n_257), .B2(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_224), .A2(n_339), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_231), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_235), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g680 ( .A(n_237), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_239), .A2(n_240), .B1(n_473), .B2(n_474), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_244), .A2(n_247), .B1(n_474), .B2(n_506), .Y(n_505) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_479), .B(n_656), .C(n_665), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_250), .A2(n_479), .B(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g250 ( .A1(n_251), .A2(n_394), .B1(n_477), .B2(n_478), .Y(n_250) );
INVx1_ASAP7_75t_L g477 ( .A(n_251), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_253), .B1(n_358), .B2(n_392), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2x1_ASAP7_75t_L g254 ( .A(n_255), .B(n_318), .Y(n_254) );
NAND4xp25_ASAP7_75t_SL g255 ( .A(n_256), .B(n_291), .C(n_300), .D(n_307), .Y(n_255) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_258), .Y(n_501) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_258), .Y(n_566) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_270), .Y(n_258) );
AND2x4_ASAP7_75t_L g303 ( .A(n_259), .B(n_295), .Y(n_303) );
AND2x4_ASAP7_75t_L g311 ( .A(n_259), .B(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g315 ( .A(n_259), .B(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g381 ( .A(n_259), .B(n_299), .Y(n_381) );
AND2x4_ASAP7_75t_L g387 ( .A(n_259), .B(n_312), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_259), .B(n_316), .Y(n_388) );
AND2x4_ASAP7_75t_L g390 ( .A(n_259), .B(n_295), .Y(n_390) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_268), .Y(n_259) );
AND2x2_ASAP7_75t_L g322 ( .A(n_260), .B(n_269), .Y(n_322) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g294 ( .A(n_261), .B(n_269), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
NAND2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g267 ( .A(n_263), .Y(n_267) );
INVx3_ASAP7_75t_L g274 ( .A(n_263), .Y(n_274) );
NAND2xp33_ASAP7_75t_L g280 ( .A(n_263), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_263), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_264), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_266), .A2(n_290), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g330 ( .A(n_269), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g283 ( .A(n_270), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g382 ( .A(n_270), .B(n_284), .Y(n_382) );
AND2x4_ASAP7_75t_L g385 ( .A(n_270), .B(n_294), .Y(n_385) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g299 ( .A(n_271), .Y(n_299) );
OR2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
AND2x4_ASAP7_75t_L g295 ( .A(n_272), .B(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g312 ( .A(n_272), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
AND2x2_ASAP7_75t_L g326 ( .A(n_272), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_274), .B(n_279), .Y(n_278) );
INVxp67_ASAP7_75t_L g286 ( .A(n_274), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g356 ( .A(n_275), .B(n_285), .C(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g296 ( .A(n_276), .Y(n_296) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
BUFx3_ASAP7_75t_L g644 ( .A(n_282), .Y(n_644) );
BUFx12f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx6_ASAP7_75t_L g464 ( .A(n_283), .Y(n_464) );
AND2x4_ASAP7_75t_L g306 ( .A(n_284), .B(n_295), .Y(n_306) );
AND2x4_ASAP7_75t_L g347 ( .A(n_284), .B(n_316), .Y(n_347) );
AND2x4_ASAP7_75t_L g372 ( .A(n_284), .B(n_316), .Y(n_372) );
AND2x4_ASAP7_75t_L g391 ( .A(n_284), .B(n_295), .Y(n_391) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_289), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
BUFx8_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_293), .Y(n_503) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x4_ASAP7_75t_L g298 ( .A(n_294), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_316), .Y(n_340) );
AND2x2_ASAP7_75t_L g345 ( .A(n_294), .B(n_312), .Y(n_345) );
AND2x4_ASAP7_75t_L g369 ( .A(n_294), .B(n_312), .Y(n_369) );
AND2x4_ASAP7_75t_L g384 ( .A(n_294), .B(n_295), .Y(n_384) );
AND2x2_ASAP7_75t_L g467 ( .A(n_294), .B(n_295), .Y(n_467) );
AND2x2_ASAP7_75t_L g583 ( .A(n_294), .B(n_316), .Y(n_583) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_297), .Y(n_643) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_298), .Y(n_468) );
BUFx12f_ASAP7_75t_L g508 ( .A(n_298), .Y(n_508) );
BUFx3_ASAP7_75t_L g602 ( .A(n_298), .Y(n_602) );
BUFx12f_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx12f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_303), .Y(n_470) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_303), .Y(n_599) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g471 ( .A(n_305), .Y(n_471) );
INVx2_ASAP7_75t_L g556 ( .A(n_305), .Y(n_556) );
INVx4_ASAP7_75t_L g600 ( .A(n_305), .Y(n_600) );
INVx1_ASAP7_75t_L g653 ( .A(n_305), .Y(n_653) );
INVx8_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx4f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx12f_ASAP7_75t_L g473 ( .A(n_311), .Y(n_473) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_311), .Y(n_506) );
AND2x4_ASAP7_75t_L g321 ( .A(n_312), .B(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g368 ( .A(n_312), .B(n_322), .Y(n_368) );
AND2x4_ASAP7_75t_L g316 ( .A(n_313), .B(n_317), .Y(n_316) );
BUFx3_ASAP7_75t_L g649 ( .A(n_314), .Y(n_649) );
BUFx5_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_315), .Y(n_474) );
INVx1_ASAP7_75t_L g597 ( .A(n_315), .Y(n_597) );
AND2x4_ASAP7_75t_L g336 ( .A(n_316), .B(n_322), .Y(n_336) );
AND2x2_ASAP7_75t_L g374 ( .A(n_316), .B(n_322), .Y(n_374) );
NAND4xp25_ASAP7_75t_L g318 ( .A(n_319), .B(n_333), .C(n_341), .D(n_348), .Y(n_318) );
INVx4_ASAP7_75t_L g496 ( .A(n_320), .Y(n_496) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx3_ASAP7_75t_L g423 ( .A(n_321), .Y(n_423) );
BUFx3_ASAP7_75t_L g628 ( .A(n_321), .Y(n_628) );
INVx1_ASAP7_75t_L g893 ( .A(n_321), .Y(n_893) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g451 ( .A(n_324), .Y(n_451) );
INVx2_ASAP7_75t_L g549 ( .A(n_324), .Y(n_549) );
INVx2_ASAP7_75t_L g615 ( .A(n_324), .Y(n_615) );
INVx5_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx4f_ASAP7_75t_L g498 ( .A(n_325), .Y(n_498) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_330), .Y(n_325) );
AND2x2_ASAP7_75t_L g371 ( .A(n_326), .B(n_330), .Y(n_371) );
AND2x4_ASAP7_75t_L g432 ( .A(n_326), .B(n_330), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_L g352 ( .A(n_328), .Y(n_352) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx3_ASAP7_75t_L g611 ( .A(n_335), .Y(n_611) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_336), .Y(n_437) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_336), .Y(n_456) );
BUFx3_ASAP7_75t_L g510 ( .A(n_336), .Y(n_510) );
BUFx8_ASAP7_75t_SL g551 ( .A(n_336), .Y(n_551) );
INVx2_ASAP7_75t_L g924 ( .A(n_336), .Y(n_924) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g366 ( .A(n_340), .Y(n_366) );
INVx3_ASAP7_75t_L g454 ( .A(n_340), .Y(n_454) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g616 ( .A(n_343), .Y(n_616) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g932 ( .A(n_344), .Y(n_932) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g450 ( .A(n_345), .Y(n_450) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_345), .Y(n_490) );
INVx3_ASAP7_75t_L g492 ( .A(n_346), .Y(n_492) );
BUFx3_ASAP7_75t_L g928 ( .A(n_346), .Y(n_928) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_347), .Y(n_552) );
INVx2_ASAP7_75t_SL g542 ( .A(n_349), .Y(n_542) );
INVx2_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_350), .Y(n_460) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_350), .Y(n_586) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx3_ASAP7_75t_L g378 ( .A(n_351), .Y(n_378) );
AO21x2_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_353), .B(n_356), .Y(n_351) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_353), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx3_ASAP7_75t_L g393 ( .A(n_360), .Y(n_393) );
XNOR2x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_379), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .C(n_370), .D(n_373), .Y(n_363) );
BUFx3_ASAP7_75t_L g896 ( .A(n_365), .Y(n_896) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_366), .Y(n_512) );
INVx2_ASAP7_75t_L g574 ( .A(n_368), .Y(n_574) );
INVx2_ASAP7_75t_L g435 ( .A(n_369), .Y(n_435) );
INVx1_ASAP7_75t_L g577 ( .A(n_369), .Y(n_577) );
INVx2_ASAP7_75t_L g579 ( .A(n_372), .Y(n_579) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_374), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_377), .B(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g516 ( .A(n_377), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_377), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_377), .B(n_926), .Y(n_925) );
INVx4_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g426 ( .A(n_378), .Y(n_426) );
NAND4xp25_ASAP7_75t_L g379 ( .A(n_380), .B(n_383), .C(n_386), .D(n_389), .Y(n_379) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g478 ( .A(n_394), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_414), .B1(n_415), .B2(n_475), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_397), .Y(n_476) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_409), .Y(n_401) );
NAND4xp25_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .C(n_405), .D(n_406), .Y(n_402) );
NAND4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .C(n_412), .D(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
XOR2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_445), .Y(n_418) );
INVx1_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
NOR2x1_ASAP7_75t_L g420 ( .A(n_421), .B(n_438), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_427), .C(n_436), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_426), .B(n_609), .Y(n_608) );
INVx4_ASAP7_75t_L g639 ( .A(n_426), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_433), .B2(n_435), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
OAI21xp5_ASAP7_75t_L g897 ( .A1(n_431), .A2(n_898), .B(n_899), .Y(n_897) );
INVx4_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
CKINVDCx9p33_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
NAND4xp25_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .C(n_441), .D(n_442), .Y(n_438) );
XNOR2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NOR2xp67_ASAP7_75t_L g447 ( .A(n_448), .B(n_461), .Y(n_447) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .C(n_455), .D(n_457), .Y(n_448) );
INVx2_ASAP7_75t_L g630 ( .A(n_450), .Y(n_630) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g522 ( .A(n_454), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_L g900 ( .A(n_460), .Y(n_900) );
NAND4xp25_ASAP7_75t_SL g461 ( .A(n_462), .B(n_465), .C(n_469), .D(n_472), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx5_ASAP7_75t_L g545 ( .A(n_464), .Y(n_545) );
INVx3_ASAP7_75t_L g567 ( .A(n_464), .Y(n_567) );
INVx1_ASAP7_75t_L g942 ( .A(n_464), .Y(n_942) );
BUFx4f_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_467), .Y(n_529) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_470), .Y(n_646) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
XNOR2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_558), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OA22x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_517), .B1(n_518), .B2(n_557), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g557 ( .A(n_484), .Y(n_557) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND4xp75_ASAP7_75t_L g486 ( .A(n_487), .B(n_499), .C(n_504), .D(n_509), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_488) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_497), .Y(n_494) );
INVx2_ASAP7_75t_SL g636 ( .A(n_498), .Y(n_636) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
BUFx3_ASAP7_75t_L g647 ( .A(n_501), .Y(n_647) );
BUFx3_ASAP7_75t_L g651 ( .A(n_503), .Y(n_651) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_507), .Y(n_504) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g539 ( .A(n_512), .Y(n_539) );
INVx2_ASAP7_75t_L g634 ( .A(n_512), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
XNOR2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_535), .Y(n_518) );
NAND3x1_ASAP7_75t_L g520 ( .A(n_521), .B(n_526), .C(n_530), .Y(n_520) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND4x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .C(n_533), .D(n_534), .Y(n_530) );
XOR2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
NAND4xp75_ASAP7_75t_L g537 ( .A(n_538), .B(n_543), .C(n_547), .D(n_553), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .Y(n_543) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_551), .Y(n_624) );
BUFx3_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_619), .B1(n_620), .B2(n_654), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g655 ( .A(n_560), .Y(n_655) );
AO22x2_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_587), .B1(n_617), .B2(n_618), .Y(n_560) );
INVx2_ASAP7_75t_L g617 ( .A(n_561), .Y(n_617) );
NAND4xp75_ASAP7_75t_L g562 ( .A(n_563), .B(n_568), .C(n_571), .D(n_581), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B(n_575), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_576) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g618 ( .A(n_589), .Y(n_618) );
INVx2_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
XNOR2x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_604), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_598), .C(n_601), .D(n_603), .Y(n_593) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_612), .C(n_614), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_641), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .C(n_631), .Y(n_622) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_640), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND4xp25_ASAP7_75t_SL g641 ( .A(n_642), .B(n_645), .C(n_648), .D(n_650), .Y(n_641) );
BUFx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx10_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_663), .C(n_664), .Y(n_659) );
AND2x2_ASAP7_75t_L g910 ( .A(n_660), .B(n_911), .Y(n_910) );
AND2x2_ASAP7_75t_L g914 ( .A(n_660), .B(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OA21x2_ASAP7_75t_L g950 ( .A1(n_661), .A2(n_700), .B(n_951), .Y(n_950) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g677 ( .A(n_662), .B(n_678), .Y(n_677) );
AND3x4_ASAP7_75t_L g699 ( .A(n_662), .B(n_679), .C(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g915 ( .A(n_663), .B(n_911), .Y(n_915) );
INVx1_ASAP7_75t_L g911 ( .A(n_664), .Y(n_911) );
OAI221xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_886), .B1(n_887), .B2(n_908), .C(n_912), .Y(n_665) );
AND5x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_830), .C(n_847), .D(n_856), .E(n_876), .Y(n_666) );
AOI222xp33_ASAP7_75t_SL g667 ( .A1(n_668), .A2(n_753), .B1(n_767), .B2(n_776), .C1(n_809), .C2(n_829), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_747), .B1(n_753), .B2(n_758), .C(n_763), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_726), .C(n_739), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_693), .Y(n_670) );
AND2x2_ASAP7_75t_L g881 ( .A(n_671), .B(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_672), .A2(n_727), .B1(n_732), .B2(n_736), .C(n_738), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_672), .B(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_L g826 ( .A(n_672), .Y(n_826) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx3_ASAP7_75t_L g734 ( .A(n_673), .Y(n_734) );
AND2x2_ASAP7_75t_L g750 ( .A(n_673), .B(n_748), .Y(n_750) );
OR2x2_ASAP7_75t_L g784 ( .A(n_673), .B(n_742), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_673), .B(n_696), .Y(n_786) );
AND2x2_ASAP7_75t_L g798 ( .A(n_673), .B(n_742), .Y(n_798) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_685), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_681), .B1(n_682), .B2(n_684), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g754 ( .A1(n_675), .A2(n_682), .B1(n_755), .B2(n_756), .C(n_757), .Y(n_754) );
INVx3_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
AND2x4_ASAP7_75t_L g688 ( .A(n_677), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g709 ( .A(n_677), .B(n_689), .Y(n_709) );
AND2x2_ASAP7_75t_L g722 ( .A(n_677), .B(n_689), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_679), .B(n_683), .Y(n_682) );
AND2x4_ASAP7_75t_L g713 ( .A(n_679), .B(n_683), .Y(n_713) );
AND2x4_ASAP7_75t_L g725 ( .A(n_679), .B(n_683), .Y(n_725) );
CKINVDCx5p33_ASAP7_75t_R g951 ( .A(n_679), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_682), .A2(n_698), .B1(n_701), .B2(n_702), .Y(n_697) );
BUFx2_ASAP7_75t_L g886 ( .A(n_682), .Y(n_886) );
AND2x4_ASAP7_75t_L g692 ( .A(n_683), .B(n_689), .Y(n_692) );
AND2x2_ASAP7_75t_L g706 ( .A(n_683), .B(n_689), .Y(n_706) );
AND2x2_ASAP7_75t_L g723 ( .A(n_683), .B(n_689), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_690), .B2(n_691), .Y(n_685) );
INVx3_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_693), .B(n_792), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_710), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_694), .B(n_729), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_694), .B(n_792), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_694), .B(n_771), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_694), .B(n_728), .Y(n_885) );
INVx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
CKINVDCx6p67_ASAP7_75t_R g735 ( .A(n_696), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_696), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g779 ( .A(n_696), .B(n_752), .Y(n_779) );
AND2x2_ASAP7_75t_L g789 ( .A(n_696), .B(n_734), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_696), .B(n_734), .Y(n_817) );
AND2x2_ASAP7_75t_L g836 ( .A(n_696), .B(n_802), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_696), .B(n_731), .Y(n_872) );
OR2x6_ASAP7_75t_SL g696 ( .A(n_697), .B(n_703), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B1(n_707), .B2(n_708), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g791 ( .A(n_710), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_710), .B(n_728), .Y(n_851) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_715), .Y(n_710) );
CKINVDCx6p67_ASAP7_75t_R g731 ( .A(n_711), .Y(n_731) );
INVx1_ASAP7_75t_L g762 ( .A(n_711), .Y(n_762) );
OR2x2_ASAP7_75t_L g766 ( .A(n_711), .B(n_716), .Y(n_766) );
OAI32xp33_ASAP7_75t_L g782 ( .A1(n_711), .A2(n_766), .A3(n_783), .B1(n_784), .B2(n_785), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_711), .B(n_716), .Y(n_800) );
AND2x2_ASAP7_75t_L g802 ( .A(n_711), .B(n_729), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g866 ( .A(n_711), .B(n_730), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_711), .B(n_752), .Y(n_880) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
INVx2_ASAP7_75t_SL g775 ( .A(n_713), .Y(n_775) );
OR2x2_ASAP7_75t_L g783 ( .A(n_715), .B(n_729), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_715), .B(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g833 ( .A(n_715), .B(n_731), .Y(n_833) );
INVx1_ASAP7_75t_L g871 ( .A(n_715), .Y(n_871) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_716), .Y(n_730) );
AND2x2_ASAP7_75t_L g822 ( .A(n_716), .B(n_720), .Y(n_822) );
AND2x4_ASAP7_75t_SL g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g737 ( .A(n_719), .Y(n_737) );
AND2x2_ASAP7_75t_L g746 ( .A(n_719), .B(n_731), .Y(n_746) );
AND2x2_ASAP7_75t_L g752 ( .A(n_719), .B(n_730), .Y(n_752) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g729 ( .A(n_720), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .Y(n_720) );
OAI211xp5_ASAP7_75t_SL g834 ( .A1(n_727), .A2(n_785), .B(n_835), .C(n_837), .Y(n_834) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_SL g728 ( .A(n_729), .B(n_731), .Y(n_728) );
AND2x2_ASAP7_75t_L g794 ( .A(n_729), .B(n_795), .Y(n_794) );
OAI21xp33_ASAP7_75t_L g824 ( .A1(n_729), .A2(n_733), .B(n_746), .Y(n_824) );
AND2x2_ASAP7_75t_L g863 ( .A(n_729), .B(n_839), .Y(n_863) );
OAI222xp33_ASAP7_75t_L g739 ( .A1(n_730), .A2(n_740), .B1(n_745), .B2(n_747), .C1(n_749), .C2(n_751), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_730), .B(n_761), .Y(n_760) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_730), .A2(n_798), .B1(n_811), .B2(n_812), .Y(n_810) );
AND2x2_ASAP7_75t_L g795 ( .A(n_731), .B(n_735), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_731), .B(n_752), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_731), .B(n_822), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_731), .B(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_731), .B(n_779), .Y(n_858) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_733), .B(n_768), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AND2x2_ASAP7_75t_L g741 ( .A(n_734), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g764 ( .A(n_734), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_734), .B(n_790), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_734), .B(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_734), .B(n_863), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_735), .B(n_741), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_735), .B(n_760), .Y(n_759) );
NOR2x1p5_ASAP7_75t_L g765 ( .A(n_735), .B(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_735), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g814 ( .A(n_735), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_735), .B(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g839 ( .A(n_735), .B(n_761), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_735), .B(n_750), .Y(n_849) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_735), .B(n_784), .Y(n_855) );
INVx1_ASAP7_75t_L g816 ( .A(n_736), .Y(n_816) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g877 ( .A(n_740), .Y(n_877) );
INVx1_ASAP7_75t_L g823 ( .A(n_741), .Y(n_823) );
INVx2_ASAP7_75t_L g748 ( .A(n_742), .Y(n_748) );
AND2x2_ASAP7_75t_L g861 ( .A(n_742), .B(n_771), .Y(n_861) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g801 ( .A1(n_746), .A2(n_802), .B1(n_803), .B2(n_805), .C(n_806), .Y(n_801) );
AOI211xp5_ASAP7_75t_L g818 ( .A1(n_746), .A2(n_819), .B(n_820), .C(n_827), .Y(n_818) );
OAI211xp5_ASAP7_75t_SL g776 ( .A1(n_747), .A2(n_777), .B(n_780), .C(n_801), .Y(n_776) );
INVx3_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g790 ( .A(n_748), .B(n_771), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_748), .B(n_770), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_748), .B(n_771), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_749), .A2(n_865), .B1(n_867), .B2(n_869), .C(n_873), .Y(n_864) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
BUFx3_ASAP7_75t_L g829 ( .A(n_754), .Y(n_829) );
NOR3xp33_ASAP7_75t_L g944 ( .A(n_756), .B(n_935), .C(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AND2x2_ASAP7_75t_L g778 ( .A(n_761), .B(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx3_ASAP7_75t_L g781 ( .A(n_767), .Y(n_781) );
OAI311xp33_ASAP7_75t_L g820 ( .A1(n_767), .A2(n_821), .A3(n_823), .B1(n_824), .C1(n_825), .Y(n_820) );
INVx3_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx3_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_769), .B(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_770), .B(n_794), .Y(n_793) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g804 ( .A(n_771), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_771), .B(n_798), .Y(n_808) );
AND2x2_ASAP7_75t_L g845 ( .A(n_771), .B(n_846), .Y(n_845) );
AND2x4_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AOI211xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B(n_787), .C(n_796), .Y(n_780) );
INVx1_ASAP7_75t_L g846 ( .A(n_784), .Y(n_846) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_790), .B1(n_791), .B2(n_792), .C(n_793), .Y(n_787) );
INVx1_ASAP7_75t_L g812 ( .A(n_790), .Y(n_812) );
OAI221xp5_ASAP7_75t_SL g809 ( .A1(n_792), .A2(n_810), .B1(n_813), .B2(n_815), .C(n_818), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_795), .B(n_822), .Y(n_875) );
AOI21xp33_ASAP7_75t_SL g796 ( .A1(n_797), .A2(n_799), .B(n_800), .Y(n_796) );
AOI211xp5_ASAP7_75t_SL g856 ( .A1(n_798), .A2(n_857), .B(n_859), .C(n_864), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_800), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g878 ( .A(n_800), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_802), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g828 ( .A(n_802), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g865 ( .A(n_802), .B(n_866), .Y(n_865) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_808), .Y(n_806) );
INVx1_ASAP7_75t_L g811 ( .A(n_807), .Y(n_811) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_812), .A2(n_819), .B1(n_831), .B2(n_834), .C(n_840), .Y(n_830) );
CKINVDCx14_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
AND2x2_ASAP7_75t_L g838 ( .A(n_822), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g843 ( .A(n_822), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_826), .B(n_836), .Y(n_835) );
AOI322xp5_ASAP7_75t_L g876 ( .A1(n_829), .A2(n_861), .A3(n_877), .B1(n_878), .B2(n_879), .C1(n_881), .C2(n_884), .Y(n_876) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_844), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_846), .B(n_868), .Y(n_867) );
OAI21xp33_ASAP7_75t_L g873 ( .A1(n_846), .A2(n_861), .B(n_874), .Y(n_873) );
AOI211xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_850), .B(n_852), .C(n_853), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVxp67_ASAP7_75t_SL g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_862), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
INVx1_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_SL g907 ( .A(n_888), .Y(n_907) );
HB1xp67_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
NOR2x1_ASAP7_75t_SL g889 ( .A(n_890), .B(n_901), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g890 ( .A(n_891), .B(n_894), .C(n_895), .Y(n_890) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND4xp25_ASAP7_75t_SL g901 ( .A(n_902), .B(n_903), .C(n_904), .D(n_905), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_909), .Y(n_908) );
BUFx3_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
BUFx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NOR2x1_ASAP7_75t_L g920 ( .A(n_921), .B(n_933), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_927), .C(n_929), .Y(n_921) );
INVx1_ASAP7_75t_L g947 ( .A(n_922), .Y(n_947) );
INVx2_ASAP7_75t_SL g923 ( .A(n_924), .Y(n_923) );
INVxp67_ASAP7_75t_SL g948 ( .A(n_927), .Y(n_948) );
INVx1_ASAP7_75t_L g945 ( .A(n_929), .Y(n_945) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g933 ( .A(n_934), .B(n_938), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
NOR3xp33_ASAP7_75t_L g946 ( .A(n_939), .B(n_947), .C(n_948), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_940), .B(n_941), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_946), .Y(n_943) );
BUFx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
endmodule