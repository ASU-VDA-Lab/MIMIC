module fake_jpeg_17131_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_34),
.B(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_42),
.Y(n_47)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_25),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_66),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_69),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_32),
.Y(n_63)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_28),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_8),
.B(n_9),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_28),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_10),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_37),
.B(n_33),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_29),
.B1(n_24),
.B2(n_66),
.Y(n_74)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_20),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_91),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_72),
.B(n_74),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_40),
.B1(n_26),
.B2(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_81),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_3),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_77),
.C(n_89),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_26),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_67),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_3),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_83),
.Y(n_103)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_19),
.B1(n_7),
.B2(n_6),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_8),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_70),
.Y(n_104)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

CKINVDCx11_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_88),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_52),
.A2(n_19),
.B1(n_9),
.B2(n_10),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_63),
.B(n_50),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_64),
.Y(n_107)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_62),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_79),
.B(n_73),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_95),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_102),
.B(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_56),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_105),
.B(n_106),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_56),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_109),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_59),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_77),
.C(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_12),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_58),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_14),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_115),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_133),
.B(n_124),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_80),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.C(n_123),
.Y(n_137)
);

NOR4xp25_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_72),
.C(n_92),
.D(n_91),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_126),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_73),
.C(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_125),
.A2(n_129),
.B(n_100),
.Y(n_140)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_76),
.C(n_90),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_75),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_74),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_R g133 ( 
.A(n_101),
.B(n_78),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_108),
.B(n_110),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_139),
.B(n_148),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_108),
.C(n_97),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_120),
.C(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_128),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_99),
.B1(n_111),
.B2(n_114),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_149),
.B1(n_121),
.B2(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_146),
.A2(n_147),
.B1(n_87),
.B2(n_96),
.Y(n_151)
);

AOI21x1_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_99),
.B(n_114),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_102),
.B(n_116),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_152),
.Y(n_164)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_156),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_117),
.C(n_53),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_93),
.Y(n_169)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_159),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_147),
.A2(n_142),
.B1(n_141),
.B2(n_136),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_141),
.B1(n_138),
.B2(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_162),
.B(n_164),
.Y(n_172)
);

FAx1_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_139),
.CI(n_148),
.CON(n_165),
.SN(n_165)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_165),
.B(n_93),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_156),
.A2(n_140),
.B1(n_135),
.B2(n_149),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_151),
.B1(n_150),
.B2(n_155),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_157),
.C(n_158),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_173),
.C(n_161),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_14),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_175),
.B(n_167),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_53),
.B(n_61),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_178),
.B(n_163),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_179),
.C(n_165),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_162),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_166),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_182),
.C(n_61),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_165),
.B(n_53),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_61),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_185),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);


endmodule