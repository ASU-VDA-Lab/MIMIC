module fake_netlist_1_6200_n_720 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_720);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_720;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_141;
wire n_119;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g79 ( .A(n_65), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_28), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_64), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_7), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_26), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_27), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_36), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_60), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_44), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_52), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_25), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_37), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_72), .Y(n_94) );
INVxp67_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_54), .Y(n_96) );
NOR2xp67_ASAP7_75t_L g97 ( .A(n_21), .B(n_77), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_29), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_5), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_43), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_40), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_15), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_16), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_78), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_5), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_69), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_74), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_30), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_62), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_12), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_56), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_38), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_45), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_10), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_34), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_35), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_67), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_23), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_19), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_32), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_33), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_116), .B(n_0), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_81), .B(n_0), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_79), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_79), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_100), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_83), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_98), .B(n_1), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_83), .B(n_1), .Y(n_140) );
BUFx8_ASAP7_75t_L g141 ( .A(n_127), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_124), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_83), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_87), .Y(n_145) );
AOI22x1_ASAP7_75t_SL g146 ( .A1(n_118), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_127), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_124), .B(n_2), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_106), .B(n_6), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_127), .Y(n_150) );
NOR2x1_ASAP7_75t_L g151 ( .A(n_89), .B(n_6), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_127), .Y(n_153) );
BUFx8_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_118), .B(n_7), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_93), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_126), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_80), .B(n_84), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_99), .B(n_8), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_107), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_96), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_110), .B(n_8), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_113), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_102), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_121), .B(n_9), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_104), .Y(n_168) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_125), .B(n_49), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_105), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_108), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_171), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_134), .B(n_109), .Y(n_173) );
NAND2xp33_ASAP7_75t_L g174 ( .A(n_171), .B(n_111), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_162), .B(n_109), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_149), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_154), .B(n_111), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_130), .Y(n_180) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_171), .B(n_122), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_171), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_154), .B(n_129), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
NOR2x1p5_ASAP7_75t_L g185 ( .A(n_137), .B(n_122), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_171), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_171), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_130), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_134), .B(n_95), .Y(n_190) );
BUFx10_ASAP7_75t_L g191 ( .A(n_129), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_132), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_145), .B(n_90), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_132), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_145), .B(n_123), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_139), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_141), .Y(n_199) );
INVx5_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_135), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_148), .Y(n_202) );
INVxp33_ASAP7_75t_SL g203 ( .A(n_149), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_154), .B(n_90), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_148), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_154), .B(n_115), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_165), .B(n_88), .Y(n_207) );
AND2x6_ASAP7_75t_L g208 ( .A(n_129), .B(n_112), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
OR2x2_ASAP7_75t_L g211 ( .A(n_156), .B(n_120), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_135), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_152), .B(n_88), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_159), .B(n_115), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_152), .B(n_101), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_158), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_159), .B(n_119), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_155), .B(n_85), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_155), .B(n_117), .Y(n_223) );
BUFx6f_ASAP7_75t_SL g224 ( .A(n_169), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_161), .A2(n_114), .B1(n_103), .B2(n_82), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_169), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_157), .B(n_103), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_128), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_128), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_135), .Y(n_230) );
BUFx8_ASAP7_75t_SL g231 ( .A(n_164), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g232 ( .A1(n_167), .A2(n_82), .B1(n_97), .B2(n_13), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_157), .B(n_10), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_160), .B(n_50), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_143), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_160), .B(n_47), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_213), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_179), .B(n_191), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_213), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_175), .B(n_170), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_218), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_218), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_179), .B(n_169), .Y(n_244) );
AND2x4_ASAP7_75t_L g245 ( .A(n_215), .B(n_151), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_224), .A2(n_170), .B1(n_166), .B2(n_151), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
NAND3xp33_ASAP7_75t_SL g248 ( .A(n_177), .B(n_140), .C(n_163), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_175), .B(n_170), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_228), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_224), .A2(n_168), .B1(n_163), .B2(n_166), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_173), .B(n_166), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_228), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_224), .A2(n_166), .B1(n_168), .B2(n_163), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_194), .B(n_168), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_215), .B(n_221), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_179), .B(n_141), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_221), .B(n_128), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_220), .B(n_142), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_207), .B(n_128), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_229), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_205), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_205), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_220), .B(n_142), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_207), .B(n_142), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_220), .B(n_131), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_217), .B(n_142), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_190), .B(n_222), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_211), .B(n_131), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_216), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_199), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_191), .B(n_141), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_226), .A2(n_146), .B1(n_131), .B2(n_147), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_234), .B(n_131), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_208), .B(n_138), .Y(n_277) );
INVx3_ASAP7_75t_L g278 ( .A(n_191), .Y(n_278) );
NAND2xp33_ASAP7_75t_L g279 ( .A(n_208), .B(n_153), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_176), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_183), .B(n_146), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_211), .B(n_11), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_176), .Y(n_283) );
OAI22xp5_ASAP7_75t_SL g284 ( .A1(n_225), .A2(n_13), .B1(n_14), .B2(n_144), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_176), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_199), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_180), .A2(n_143), .B1(n_144), .B2(n_147), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_208), .B(n_138), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_227), .B(n_14), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_200), .B(n_138), .Y(n_290) );
NOR2x1p5_ASAP7_75t_L g291 ( .A(n_231), .B(n_185), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_208), .B(n_138), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_172), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_184), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_203), .A2(n_143), .B1(n_147), .B2(n_144), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_189), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_200), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_193), .A2(n_153), .B1(n_150), .B2(n_136), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_197), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_209), .B(n_138), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_198), .B(n_138), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_172), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_209), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_210), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_182), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_SL g306 ( .A1(n_235), .A2(n_153), .B(n_150), .C(n_136), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_214), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_238), .B(n_203), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_239), .A2(n_206), .B(n_178), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_239), .A2(n_204), .B(n_200), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
OAI21xp5_ASAP7_75t_L g312 ( .A1(n_253), .A2(n_208), .B(n_196), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_240), .B(n_245), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_244), .A2(n_208), .B1(n_202), .B2(n_200), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_244), .A2(n_202), .B1(n_200), .B2(n_223), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_267), .Y(n_316) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_252), .A2(n_202), .B(n_174), .Y(n_317) );
BUFx4f_ASAP7_75t_L g318 ( .A(n_282), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_270), .B(n_202), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_245), .B(n_202), .Y(n_320) );
OR2x4_ASAP7_75t_L g321 ( .A(n_281), .B(n_231), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_291), .B(n_233), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_256), .B(n_232), .Y(n_323) );
NOR2xp33_ASAP7_75t_SL g324 ( .A(n_286), .B(n_187), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_272), .B(n_237), .Y(n_325) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_284), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_241), .B(n_174), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_267), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_251), .A2(n_186), .B1(n_187), .B2(n_182), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_251), .A2(n_186), .B1(n_230), .B2(n_212), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_263), .A2(n_181), .B(n_236), .C(n_212), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_259), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_250), .Y(n_333) );
AOI33xp33_ASAP7_75t_L g334 ( .A1(n_274), .A2(n_236), .A3(n_230), .B1(n_201), .B2(n_195), .B3(n_192), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
AOI221x1_ASAP7_75t_L g336 ( .A1(n_248), .A2(n_133), .B1(n_136), .B2(n_150), .C(n_153), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_264), .A2(n_181), .B(n_195), .C(n_192), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_272), .B(n_201), .Y(n_338) );
CKINVDCx8_ASAP7_75t_R g339 ( .A(n_281), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_289), .B(n_17), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_269), .A2(n_188), .B(n_22), .C(n_24), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_255), .A2(n_188), .B(n_153), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_278), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_261), .B(n_18), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_280), .A2(n_153), .B(n_150), .Y(n_345) );
INVx5_ASAP7_75t_L g346 ( .A(n_278), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_303), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_249), .B(n_150), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_294), .A2(n_150), .B(n_136), .C(n_133), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_266), .B(n_133), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_260), .B(n_133), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_254), .B(n_136), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_260), .B(n_136), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_283), .Y(n_355) );
O2A1O1Ixp5_ASAP7_75t_L g356 ( .A1(n_257), .A2(n_31), .B(n_39), .C(n_41), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_257), .A2(n_133), .B(n_46), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_296), .A2(n_42), .B(n_51), .C(n_53), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_285), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_273), .A2(n_133), .B(n_57), .Y(n_360) );
OAI21x1_ASAP7_75t_L g361 ( .A1(n_277), .A2(n_55), .B(n_58), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_333), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_354), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_308), .B(n_265), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_323), .A2(n_265), .B1(n_304), .B2(n_299), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g366 ( .A1(n_312), .A2(n_273), .B(n_307), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_313), .B(n_275), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_332), .B(n_349), .Y(n_368) );
BUFx10_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
BUFx2_ASAP7_75t_R g370 ( .A(n_339), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_326), .A2(n_246), .B1(n_268), .B2(n_295), .Y(n_371) );
OAI22x1_ASAP7_75t_L g372 ( .A1(n_340), .A2(n_275), .B1(n_300), .B2(n_297), .Y(n_372) );
O2A1O1Ixp5_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_306), .B(n_271), .C(n_276), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_347), .B(n_258), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_348), .A2(n_262), .B(n_279), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_318), .A2(n_301), .B1(n_287), .B2(n_243), .C(n_247), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_318), .A2(n_242), .B1(n_301), .B2(n_297), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_320), .B(n_287), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_328), .B(n_320), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_327), .A2(n_288), .B(n_292), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_319), .A2(n_290), .B1(n_298), .B2(n_302), .Y(n_382) );
INVx3_ASAP7_75t_SL g383 ( .A(n_322), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_355), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_334), .A2(n_290), .B(n_298), .C(n_306), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_340), .A2(n_305), .B1(n_293), .B2(n_63), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_309), .A2(n_59), .B(n_61), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
CKINVDCx11_ASAP7_75t_R g390 ( .A(n_322), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_315), .A2(n_66), .B1(n_68), .B2(n_75), .Y(n_391) );
AO31x2_ASAP7_75t_L g392 ( .A1(n_336), .A2(n_76), .A3(n_337), .B(n_331), .Y(n_392) );
OAI21xp5_ASAP7_75t_L g393 ( .A1(n_317), .A2(n_342), .B(n_314), .Y(n_393) );
AO32x2_ASAP7_75t_L g394 ( .A1(n_329), .A2(n_330), .A3(n_361), .B1(n_341), .B2(n_356), .Y(n_394) );
A2O1A1Ixp33_ASAP7_75t_L g395 ( .A1(n_344), .A2(n_358), .B(n_310), .C(n_357), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_364), .B(n_322), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_365), .A2(n_346), .B1(n_335), .B2(n_343), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g399 ( .A1(n_395), .A2(n_324), .B(n_351), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_384), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_366), .A2(n_324), .B(n_325), .Y(n_401) );
BUFx8_ASAP7_75t_L g402 ( .A(n_380), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_360), .B(n_345), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_365), .A2(n_338), .B1(n_343), .B2(n_311), .C(n_350), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_368), .B(n_346), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_387), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_389), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
AOI21xp5_ASAP7_75t_L g409 ( .A1(n_393), .A2(n_345), .B(n_311), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_367), .B(n_346), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_371), .A2(n_321), .B1(n_335), .B2(n_377), .C(n_374), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_392), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_372), .B(n_335), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_378), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_375), .B(n_381), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_383), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_383), .B(n_390), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_371), .A2(n_391), .B1(n_376), .B2(n_382), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_391), .A2(n_382), .B1(n_370), .B2(n_385), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_392), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_373), .A2(n_388), .B(n_394), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_369), .B(n_392), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_394), .Y(n_424) );
AO21x2_ASAP7_75t_L g425 ( .A1(n_422), .A2(n_392), .B(n_394), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_407), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_407), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_411), .B(n_369), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_400), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g430 ( .A1(n_423), .A2(n_394), .B(n_420), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_406), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_400), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_412), .B(n_406), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
OR2x6_ASAP7_75t_L g436 ( .A(n_414), .B(n_417), .Y(n_436) );
BUFx2_ASAP7_75t_L g437 ( .A(n_414), .Y(n_437) );
AOI21xp5_ASAP7_75t_SL g438 ( .A1(n_419), .A2(n_397), .B(n_421), .Y(n_438) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_421), .A2(n_413), .B(n_416), .Y(n_439) );
OR2x2_ASAP7_75t_L g440 ( .A(n_408), .B(n_405), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_408), .Y(n_441) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_413), .A2(n_424), .B(n_399), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_410), .Y(n_445) );
OAI211xp5_ASAP7_75t_L g446 ( .A1(n_396), .A2(n_418), .B(n_415), .C(n_404), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_403), .A2(n_409), .B(n_401), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
OA21x2_ASAP7_75t_L g449 ( .A1(n_415), .A2(n_418), .B(n_402), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_402), .B(n_412), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_402), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_412), .B(n_407), .Y(n_452) );
AOI21x1_ASAP7_75t_L g453 ( .A1(n_423), .A2(n_421), .B(n_399), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_400), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_407), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
OAI211xp5_ASAP7_75t_L g461 ( .A1(n_411), .A2(n_274), .B(n_225), .C(n_339), .Y(n_461) );
NOR2x1_ASAP7_75t_L g462 ( .A(n_449), .B(n_443), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_432), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_443), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_431), .B(n_432), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_450), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_431), .B(n_458), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_434), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_445), .B(n_441), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_441), .B(n_457), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_427), .B(n_454), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_456), .B(n_437), .Y(n_473) );
INVx2_ASAP7_75t_SL g474 ( .A(n_459), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_435), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_454), .B(n_460), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_456), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_458), .Y(n_480) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_430), .A2(n_448), .B(n_453), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_460), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_429), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_426), .B(n_455), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_440), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_426), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_437), .B(n_440), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_456), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_455), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_459), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_459), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_436), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_456), .B(n_436), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_456), .B(n_452), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_452), .B(n_444), .Y(n_497) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_453), .A2(n_425), .B(n_439), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_436), .B(n_433), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_439), .Y(n_500) );
BUFx3_ASAP7_75t_L g501 ( .A(n_449), .Y(n_501) );
INVx3_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_439), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_425), .B(n_451), .Y(n_505) );
INVxp67_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_442), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_449), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_442), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_449), .A2(n_428), .B1(n_425), .B2(n_447), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_447), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_463), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_505), .B(n_447), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_505), .B(n_438), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_463), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_501), .B(n_438), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_505), .B(n_446), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_501), .B(n_461), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_505), .B(n_496), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_468), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_501), .B(n_508), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_496), .B(n_497), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_497), .B(n_465), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_508), .B(n_462), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_462), .B(n_473), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_468), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_465), .B(n_491), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_467), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_491), .B(n_478), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_486), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_472), .B(n_478), .Y(n_535) );
AND2x4_ASAP7_75t_L g536 ( .A(n_473), .B(n_479), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_475), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_466), .B(n_506), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_476), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_469), .B(n_483), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_464), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_483), .B(n_488), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_467), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_472), .B(n_485), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_485), .B(n_511), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_464), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_488), .B(n_495), .Y(n_547) );
NOR2xp67_ASAP7_75t_L g548 ( .A(n_464), .B(n_502), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_500), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_473), .B(n_482), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_476), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_473), .B(n_482), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_477), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_499), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_477), .B(n_480), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_500), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_495), .B(n_499), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_489), .B(n_494), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_487), .B(n_490), .Y(n_560) );
INVx4_ASAP7_75t_L g561 ( .A(n_484), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_502), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_487), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_490), .B(n_504), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_484), .B(n_494), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_504), .B(n_512), .C(n_510), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_492), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_513), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_524), .B(n_470), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_523), .B(n_474), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_523), .B(n_474), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_567), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_534), .B(n_493), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_555), .B(n_512), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_567), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_524), .B(n_493), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_513), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_544), .B(n_502), .Y(n_578) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_561), .B(n_502), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_516), .Y(n_580) );
NAND2x1_ASAP7_75t_L g581 ( .A(n_525), .B(n_503), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_516), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_555), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_521), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_544), .B(n_503), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_533), .B(n_507), .Y(n_586) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_519), .A2(n_507), .B(n_510), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_535), .B(n_503), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_521), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_533), .B(n_510), .Y(n_591) );
NAND2x1p5_ASAP7_75t_L g592 ( .A(n_561), .B(n_503), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_535), .B(n_481), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_527), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_530), .B(n_509), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_560), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_554), .B(n_481), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_547), .B(n_509), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_528), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_547), .B(n_509), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_558), .B(n_498), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_560), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_546), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_558), .B(n_498), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_529), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_530), .B(n_498), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_564), .B(n_498), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_532), .B(n_481), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_564), .B(n_529), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_541), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_522), .B(n_548), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_531), .B(n_551), .Y(n_613) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_561), .B(n_525), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_531), .B(n_551), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_520), .B(n_550), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_520), .B(n_550), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_532), .B(n_543), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_537), .B(n_539), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_537), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_543), .B(n_542), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_610), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_593), .B(n_540), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_608), .B(n_545), .Y(n_624) );
BUFx2_ASAP7_75t_SL g625 ( .A(n_611), .Y(n_625) );
AND2x4_ASAP7_75t_L g626 ( .A(n_614), .B(n_522), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_610), .Y(n_627) );
INVx2_ASAP7_75t_SL g628 ( .A(n_576), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_583), .B(n_545), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_621), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_612), .B(n_522), .Y(n_631) );
INVx2_ASAP7_75t_SL g632 ( .A(n_570), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_569), .B(n_565), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_572), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_579), .A2(n_538), .B(n_525), .C(n_541), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_613), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_608), .B(n_574), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_572), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_574), .B(n_556), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_595), .B(n_565), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_595), .B(n_552), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_613), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_578), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_615), .Y(n_644) );
OAI21xp33_ASAP7_75t_L g645 ( .A1(n_588), .A2(n_515), .B(n_518), .Y(n_645) );
AOI21xp33_ASAP7_75t_SL g646 ( .A1(n_579), .A2(n_517), .B(n_526), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_586), .B(n_539), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_586), .B(n_556), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_604), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_591), .B(n_552), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_615), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_619), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_616), .B(n_515), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_617), .B(n_536), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_619), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g656 ( .A1(n_592), .A2(n_517), .B(n_526), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_607), .B(n_601), .Y(n_657) );
OR2x2_ASAP7_75t_L g658 ( .A(n_591), .B(n_518), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_585), .B(n_536), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g660 ( .A(n_635), .B(n_604), .C(n_581), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_636), .Y(n_661) );
OAI32xp33_ASAP7_75t_L g662 ( .A1(n_649), .A2(n_592), .A3(n_573), .B1(n_605), .B2(n_618), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_645), .A2(n_573), .B1(n_519), .B2(n_517), .Y(n_663) );
OAI322xp33_ASAP7_75t_L g664 ( .A1(n_624), .A2(n_600), .A3(n_598), .B1(n_602), .B2(n_596), .C1(n_609), .C2(n_575), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_642), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_644), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_625), .B(n_571), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_651), .Y(n_668) );
NOR2x1_ASAP7_75t_L g669 ( .A(n_649), .B(n_626), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_630), .A2(n_519), .B1(n_517), .B2(n_612), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_637), .B(n_620), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_652), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_622), .B(n_597), .Y(n_673) );
INVxp67_ASAP7_75t_L g674 ( .A(n_655), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_627), .A2(n_587), .B1(n_603), .B2(n_599), .C(n_594), .Y(n_675) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_646), .A2(n_587), .B(n_526), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_626), .B(n_562), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_628), .B(n_582), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_631), .B(n_514), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_639), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_639), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_659), .B(n_536), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_671), .Y(n_683) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_669), .B(n_631), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_671), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_667), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_674), .B(n_632), .Y(n_687) );
OAI221xp5_ASAP7_75t_L g688 ( .A1(n_660), .A2(n_657), .B1(n_624), .B2(n_637), .C(n_648), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_662), .A2(n_657), .B(n_638), .C(n_634), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_661), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_665), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_676), .A2(n_653), .B1(n_623), .B2(n_629), .Y(n_692) );
OAI31xp33_ASAP7_75t_SL g693 ( .A1(n_679), .A2(n_654), .A3(n_643), .B(n_656), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_679), .Y(n_694) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_677), .Y(n_695) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_664), .A2(n_623), .B(n_648), .C(n_647), .Y(n_696) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_684), .B(n_663), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_692), .A2(n_678), .B1(n_670), .B2(n_680), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_688), .A2(n_672), .B(n_668), .Y(n_699) );
O2A1O1Ixp5_ASAP7_75t_L g700 ( .A1(n_683), .A2(n_666), .B(n_681), .C(n_673), .Y(n_700) );
BUFx6f_ASAP7_75t_L g701 ( .A(n_687), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_696), .A2(n_675), .B1(n_647), .B2(n_658), .C(n_633), .Y(n_702) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_693), .A2(n_640), .B(n_641), .C(n_650), .Y(n_703) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_689), .A2(n_584), .B1(n_606), .B2(n_590), .C(n_589), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_697), .B(n_686), .C(n_685), .Y(n_705) );
NOR4xp25_ASAP7_75t_L g706 ( .A(n_703), .B(n_691), .C(n_690), .D(n_694), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_699), .A2(n_695), .B1(n_687), .B2(n_580), .C(n_577), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g708 ( .A(n_701), .B(n_695), .Y(n_708) );
OAI211xp5_ASAP7_75t_L g709 ( .A1(n_701), .A2(n_695), .B(n_682), .C(n_514), .Y(n_709) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_708), .B(n_704), .C(n_702), .D(n_700), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_705), .B(n_698), .C(n_562), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_706), .B(n_568), .Y(n_712) );
OR4x2_ASAP7_75t_L g713 ( .A(n_710), .B(n_709), .C(n_707), .D(n_559), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_714), .B(n_711), .Y(n_715) );
OR2x6_ASAP7_75t_L g716 ( .A(n_715), .B(n_713), .Y(n_716) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_716), .A2(n_713), .B1(n_562), .B2(n_566), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_553), .B(n_559), .Y(n_718) );
AO221x2_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_553), .B1(n_563), .B2(n_549), .C(n_557), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_563), .B(n_549), .Y(n_720) );
endmodule