module fake_jpeg_27713_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_43),
.B(n_22),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_44),
.B(n_51),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_18),
.B1(n_32),
.B2(n_28),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_27),
.B1(n_23),
.B2(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_52),
.Y(n_61)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_42),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_21),
.B1(n_29),
.B2(n_30),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_65),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_35),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_69),
.B1(n_85),
.B2(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_24),
.B1(n_14),
.B2(n_11),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_49),
.A2(n_39),
.B1(n_27),
.B2(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_77),
.B1(n_60),
.B2(n_47),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_59),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_86),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_32),
.B1(n_23),
.B2(n_25),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_16),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_25),
.C(n_22),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_29),
.C(n_21),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_22),
.B1(n_30),
.B2(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_31),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_88),
.B(n_89),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_48),
.B(n_57),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_26),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_96),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_72),
.A2(n_57),
.B1(n_47),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_98),
.B1(n_68),
.B2(n_83),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_24),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_61),
.A2(n_75),
.B1(n_63),
.B2(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_89),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_64),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_110),
.B(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_16),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_103),
.B(n_107),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_64),
.B(n_0),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_84),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_110),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_69),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_121),
.B(n_54),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_122),
.A2(n_117),
.B1(n_113),
.B2(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_11),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_125),
.B(n_126),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_98),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_62),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_1),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_130),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_62),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_133),
.A2(n_90),
.B(n_70),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_102),
.C(n_99),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_146),
.C(n_124),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_112),
.A2(n_105),
.B(n_90),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_139),
.B(n_150),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_138),
.B(n_156),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_153),
.B(n_113),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_109),
.B1(n_97),
.B2(n_81),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_145),
.A2(n_120),
.B1(n_127),
.B2(n_126),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_88),
.C(n_109),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_111),
.B(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_97),
.B(n_2),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_151),
.A2(n_118),
.B(n_130),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_1),
.C(n_2),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_3),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_159),
.C(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_131),
.C(n_121),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_165),
.B1(n_149),
.B2(n_137),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_161),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_143),
.B(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_118),
.B1(n_114),
.B2(n_116),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_144),
.B1(n_149),
.B2(n_148),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_116),
.C(n_4),
.Y(n_166)
);

OAI322xp33_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_143),
.A3(n_152),
.B1(n_9),
.B2(n_10),
.C1(n_6),
.C2(n_7),
.Y(n_186)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_135),
.B(n_5),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_172),
.Y(n_183)
);

OAI321xp33_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_84),
.C(n_6),
.Y(n_173)
);

XNOR2x1_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_5),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_151),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_170),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_185),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_136),
.C(n_147),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_182),
.C(n_169),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_141),
.C(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_179),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_170),
.B(n_164),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_163),
.B1(n_174),
.B2(n_141),
.Y(n_193)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_193),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_180),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_198),
.C(n_185),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_176),
.C(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_176),
.C(n_183),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_165),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_197),
.Y(n_208)
);

AO21x2_ASAP7_75t_L g207 ( 
.A1(n_199),
.A2(n_193),
.B(n_140),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_145),
.B1(n_161),
.B2(n_205),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_203),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_204),
.A2(n_177),
.B(n_178),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_209),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_184),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_207),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_207),
.B(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_215),
.B(n_152),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_215),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_214),
.C(n_173),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_220),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_9),
.Y(n_224)
);


endmodule