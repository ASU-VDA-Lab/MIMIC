module fake_netlist_1_9254_n_41 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx2_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
INVx3_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_4), .B(n_1), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_1), .B(n_3), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_0), .B(n_11), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_14), .B(n_12), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_14), .B(n_8), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_13), .B1(n_15), .B2(n_17), .C(n_18), .Y(n_23) );
OAI21xp5_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_12), .B(n_18), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_12), .B(n_15), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_22), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
OAI321xp33_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_26), .A3(n_17), .B1(n_16), .B2(n_27), .C(n_19), .Y(n_31) );
OAI221xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_26), .B1(n_16), .B2(n_25), .C(n_5), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_16), .B1(n_2), .B2(n_3), .Y(n_33) );
OAI211xp5_ASAP7_75t_SL g34 ( .A1(n_31), .A2(n_0), .B(n_2), .C(n_5), .Y(n_34) );
INVxp67_ASAP7_75t_SL g35 ( .A(n_33), .Y(n_35) );
AND4x2_ASAP7_75t_L g36 ( .A(n_34), .B(n_6), .C(n_7), .D(n_16), .Y(n_36) );
NOR2x1_ASAP7_75t_L g37 ( .A(n_32), .B(n_16), .Y(n_37) );
XOR2xp5_ASAP7_75t_L g38 ( .A(n_36), .B(n_6), .Y(n_38) );
OR3x1_ASAP7_75t_L g39 ( .A(n_37), .B(n_7), .C(n_16), .Y(n_39) );
OAI22x1_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_35), .B1(n_39), .B2(n_37), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_40), .Y(n_41) );
endmodule