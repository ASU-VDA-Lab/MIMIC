module real_aes_462_n_255 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_255);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_255;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_693;
wire n_281;
wire n_496;
wire n_468;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_598;
wire n_404;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_668;
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_0), .A2(n_103), .B1(n_411), .B2(n_504), .Y(n_610) );
XNOR2x1_ASAP7_75t_L g544 ( .A(n_1), .B(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_2), .A2(n_237), .B1(n_381), .B2(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_3), .A2(n_189), .B1(n_373), .B2(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_4), .B(n_343), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_5), .A2(n_191), .B1(n_406), .B2(n_484), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_6), .A2(n_135), .B1(n_399), .B2(n_548), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_7), .A2(n_26), .B1(n_348), .B2(n_655), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_8), .A2(n_111), .B1(n_733), .B2(n_734), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_9), .A2(n_203), .B1(n_536), .B2(n_626), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_10), .A2(n_163), .B1(n_415), .B2(n_640), .Y(n_639) );
AO22x2_ASAP7_75t_L g282 ( .A1(n_11), .A2(n_172), .B1(n_279), .B2(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g709 ( .A(n_11), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_12), .A2(n_106), .B1(n_319), .B2(n_433), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g372 ( .A1(n_13), .A2(n_228), .B1(n_373), .B2(n_374), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_14), .A2(n_174), .B1(n_428), .B2(n_575), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_15), .A2(n_43), .B1(n_323), .B2(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g511 ( .A(n_16), .Y(n_511) );
INVx1_ASAP7_75t_L g531 ( .A(n_17), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_18), .A2(n_193), .B1(n_539), .B2(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g506 ( .A(n_19), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_20), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_21), .A2(n_68), .B1(n_516), .B2(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_22), .A2(n_164), .B1(n_292), .B2(n_433), .Y(n_559) );
AO22x2_ASAP7_75t_L g278 ( .A1(n_23), .A2(n_54), .B1(n_279), .B2(n_280), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g707 ( .A(n_23), .B(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_24), .A2(n_207), .B1(n_409), .B2(n_619), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g369 ( .A1(n_25), .A2(n_81), .B1(n_370), .B2(n_371), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_27), .A2(n_115), .B1(n_318), .B2(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_28), .A2(n_204), .B1(n_386), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_29), .A2(n_171), .B1(n_323), .B2(n_326), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_30), .A2(n_144), .B1(n_275), .B2(n_413), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_31), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_32), .A2(n_79), .B1(n_382), .B2(n_433), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_33), .A2(n_39), .B1(n_685), .B2(n_727), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_34), .A2(n_148), .B1(n_339), .B2(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_35), .A2(n_139), .B1(n_381), .B2(n_382), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_36), .A2(n_126), .B1(n_318), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_37), .A2(n_124), .B1(n_378), .B2(n_379), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_38), .A2(n_76), .B1(n_397), .B2(n_724), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_40), .A2(n_69), .B1(n_379), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_41), .A2(n_153), .B1(n_468), .B2(n_470), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_42), .A2(n_58), .B1(n_298), .B2(n_304), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_44), .A2(n_104), .B1(n_428), .B2(n_575), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_45), .A2(n_128), .B1(n_484), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_46), .A2(n_232), .B1(n_642), .B2(n_644), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_47), .A2(n_236), .B1(n_293), .B2(n_433), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_48), .A2(n_109), .B1(n_468), .B2(n_470), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_49), .A2(n_119), .B1(n_370), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_50), .A2(n_150), .B1(n_385), .B2(n_386), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_51), .A2(n_64), .B1(n_558), .B2(n_646), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_52), .A2(n_133), .B1(n_366), .B2(n_367), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_53), .A2(n_86), .B1(n_293), .B2(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_55), .A2(n_186), .B1(n_366), .B2(n_367), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_56), .A2(n_60), .B1(n_413), .B2(n_489), .Y(n_611) );
AOI22xp33_ASAP7_75t_SL g450 ( .A1(n_57), .A2(n_99), .B1(n_373), .B2(n_374), .Y(n_450) );
AO222x2_ASAP7_75t_SL g448 ( .A1(n_59), .A2(n_168), .B1(n_185), .B2(n_363), .C1(n_366), .C2(n_367), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_61), .A2(n_131), .B1(n_308), .B2(n_311), .Y(n_307) );
OA22x2_ASAP7_75t_L g560 ( .A1(n_62), .A2(n_561), .B1(n_562), .B2(n_586), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_62), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_63), .A2(n_142), .B1(n_415), .B2(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g279 ( .A(n_65), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_66), .A2(n_93), .B1(n_481), .B2(n_482), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_67), .A2(n_240), .B1(n_406), .B2(n_407), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_70), .A2(n_178), .B1(n_382), .B2(n_388), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_71), .A2(n_215), .B1(n_366), .B2(n_367), .Y(n_667) );
AOI22x1_ASAP7_75t_L g463 ( .A1(n_72), .A2(n_464), .B1(n_465), .B2(n_490), .Y(n_463) );
INVx1_ASAP7_75t_L g490 ( .A(n_72), .Y(n_490) );
INVx1_ASAP7_75t_L g523 ( .A(n_73), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_74), .A2(n_169), .B1(n_650), .B2(n_651), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_75), .A2(n_137), .B1(n_472), .B2(n_473), .Y(n_471) );
AOI222xp33_ASAP7_75t_L g627 ( .A1(n_77), .A2(n_92), .B1(n_175), .B2(n_424), .C1(n_567), .C2(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_78), .A2(n_84), .B1(n_402), .B2(n_403), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_80), .A2(n_107), .B1(n_482), .B2(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_82), .A2(n_222), .B1(n_378), .B2(n_379), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_83), .A2(n_146), .B1(n_335), .B2(n_719), .Y(n_718) );
INVx1_ASAP7_75t_SL g287 ( .A(n_85), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_85), .B(n_121), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_87), .A2(n_123), .B1(n_402), .B2(n_403), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_88), .A2(n_252), .B1(n_299), .B2(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_89), .A2(n_158), .B1(n_473), .B2(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g262 ( .A(n_90), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_91), .A2(n_206), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_94), .A2(n_199), .B1(n_370), .B2(n_371), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_95), .A2(n_125), .B1(n_366), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g435 ( .A1(n_96), .A2(n_132), .B1(n_385), .B2(n_386), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_97), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_98), .A2(n_173), .B1(n_273), .B2(n_292), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_100), .A2(n_213), .B1(n_481), .B2(n_487), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_101), .A2(n_166), .B1(n_378), .B2(n_379), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_102), .A2(n_165), .B1(n_642), .B2(n_644), .Y(n_641) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_105), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_108), .B(n_343), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_110), .A2(n_225), .B1(n_403), .B2(n_626), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g255 ( .A1(n_112), .A2(n_256), .B(n_265), .C(n_711), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_113), .A2(n_210), .B1(n_348), .B2(n_350), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_114), .A2(n_167), .B1(n_333), .B2(n_338), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_116), .A2(n_151), .B1(n_608), .B2(n_609), .Y(n_607) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_117), .A2(n_161), .B1(n_378), .B2(n_379), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_118), .A2(n_230), .B1(n_396), .B2(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g697 ( .A(n_120), .Y(n_697) );
AO22x2_ASAP7_75t_L g290 ( .A1(n_121), .A2(n_188), .B1(n_279), .B2(n_291), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_122), .A2(n_143), .B1(n_651), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_127), .A2(n_235), .B1(n_335), .B2(n_475), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_129), .A2(n_243), .B1(n_315), .B2(n_317), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_130), .A2(n_248), .B1(n_409), .B2(n_411), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_134), .A2(n_254), .B1(n_520), .B2(n_556), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_136), .A2(n_198), .B1(n_324), .B2(n_655), .Y(n_722) );
INVx1_ASAP7_75t_L g288 ( .A(n_138), .Y(n_288) );
INVx1_ASAP7_75t_L g533 ( .A(n_140), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_141), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_145), .B(n_478), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_147), .A2(n_205), .B1(n_487), .B2(n_489), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_149), .A2(n_233), .B1(n_311), .B2(n_409), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_152), .B(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_154), .A2(n_157), .B1(n_385), .B2(n_386), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_155), .A2(n_238), .B1(n_323), .B2(n_350), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_156), .B(n_344), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_159), .B(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_160), .A2(n_239), .B1(n_539), .B2(n_540), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_162), .A2(n_217), .B1(n_508), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_170), .A2(n_221), .B1(n_388), .B2(n_389), .Y(n_387) );
XNOR2x1_ASAP7_75t_L g499 ( .A(n_176), .B(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_177), .A2(n_184), .B1(n_381), .B2(n_389), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_179), .B(n_343), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_180), .A2(n_713), .B1(n_714), .B2(n_737), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_180), .Y(n_737) );
INVx1_ASAP7_75t_L g657 ( .A(n_181), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_182), .A2(n_190), .B1(n_370), .B2(n_371), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_183), .A2(n_216), .B1(n_381), .B2(n_382), .Y(n_380) );
AOI221x1_ASAP7_75t_L g515 ( .A1(n_187), .A2(n_208), .B1(n_308), .B2(n_516), .C(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g505 ( .A(n_192), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_194), .B(n_478), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_195), .A2(n_234), .B1(n_472), .B2(n_473), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_196), .A2(n_197), .B1(n_311), .B2(n_504), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_200), .A2(n_251), .B1(n_382), .B2(n_433), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_201), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g705 ( .A(n_201), .Y(n_705) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_202), .Y(n_364) );
INVx1_ASAP7_75t_L g259 ( .A(n_209), .Y(n_259) );
AND2x2_ASAP7_75t_R g739 ( .A(n_209), .B(n_705), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_211), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_212), .B(n_394), .Y(n_393) );
XNOR2xp5_ASAP7_75t_L g740 ( .A(n_214), .B(n_715), .Y(n_740) );
INVxp67_ASAP7_75t_L g745 ( .A(n_214), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_218), .A2(n_249), .B1(n_381), .B2(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_219), .A2(n_246), .B1(n_475), .B2(n_476), .Y(n_474) );
INVxp67_ASAP7_75t_L g264 ( .A(n_220), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_223), .Y(n_576) );
AOI22x1_ASAP7_75t_SL g597 ( .A1(n_224), .A2(n_598), .B1(n_599), .B2(n_612), .Y(n_597) );
INVx1_ASAP7_75t_L g612 ( .A(n_224), .Y(n_612) );
XNOR2xp5_ASAP7_75t_L g269 ( .A(n_226), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g522 ( .A(n_227), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_229), .A2(n_250), .B1(n_385), .B2(n_386), .Y(n_458) );
INVx1_ASAP7_75t_L g510 ( .A(n_231), .Y(n_510) );
INVx1_ASAP7_75t_L g527 ( .A(n_241), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_242), .B(n_344), .Y(n_422) );
OA22x2_ASAP7_75t_L g613 ( .A1(n_244), .A2(n_614), .B1(n_615), .B2(n_630), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_244), .Y(n_614) );
AO21x2_ASAP7_75t_L g632 ( .A1(n_244), .A2(n_615), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g416 ( .A(n_245), .Y(n_416) );
XNOR2xp5_ASAP7_75t_L g358 ( .A(n_247), .B(n_359), .Y(n_358) );
AOI22x1_ASAP7_75t_L g445 ( .A1(n_253), .A2(n_446), .B1(n_459), .B2(n_460), .Y(n_445) );
INVx1_ASAP7_75t_L g460 ( .A(n_253), .Y(n_460) );
BUFx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR2x1_ASAP7_75t_R g257 ( .A(n_258), .B(n_260), .Y(n_257) );
OR2x2_ASAP7_75t_L g744 ( .A(n_258), .B(n_261), .Y(n_744) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_259), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_495), .B(n_701), .C(n_702), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_266), .B(n_495), .Y(n_701) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_354), .B1(n_355), .B2(n_494), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_269), .Y(n_494) );
NOR2xp67_ASAP7_75t_L g270 ( .A(n_271), .B(n_321), .Y(n_270) );
NAND4xp25_ASAP7_75t_L g271 ( .A(n_272), .B(n_297), .C(n_307), .D(n_314), .Y(n_271) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_274), .A2(n_510), .B1(n_511), .B2(n_512), .Y(n_509) );
INVx3_ASAP7_75t_L g558 ( .A(n_274), .Y(n_558) );
INVx1_ASAP7_75t_SL g687 ( .A(n_274), .Y(n_687) );
INVx2_ASAP7_75t_L g727 ( .A(n_274), .Y(n_727) );
INVx6_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
BUFx3_ASAP7_75t_L g489 ( .A(n_275), .Y(n_489) );
AND2x4_ASAP7_75t_L g275 ( .A(n_276), .B(n_284), .Y(n_275) );
AND2x4_ASAP7_75t_L g310 ( .A(n_276), .B(n_294), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_276), .B(n_303), .Y(n_316) );
AND2x2_ASAP7_75t_L g346 ( .A(n_276), .B(n_329), .Y(n_346) );
AND2x4_ASAP7_75t_L g363 ( .A(n_276), .B(n_329), .Y(n_363) );
AND2x6_ASAP7_75t_L g381 ( .A(n_276), .B(n_303), .Y(n_381) );
AND2x2_ASAP7_75t_L g385 ( .A(n_276), .B(n_284), .Y(n_385) );
AND2x2_ASAP7_75t_L g388 ( .A(n_276), .B(n_294), .Y(n_388) );
AND2x2_ASAP7_75t_L g584 ( .A(n_276), .B(n_284), .Y(n_584) );
AND2x4_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g296 ( .A(n_278), .B(n_282), .Y(n_296) );
INVx1_ASAP7_75t_L g302 ( .A(n_278), .Y(n_302) );
AND2x4_ASAP7_75t_L g320 ( .A(n_278), .B(n_281), .Y(n_320) );
INVx2_ASAP7_75t_L g280 ( .A(n_279), .Y(n_280) );
INVx1_ASAP7_75t_L g283 ( .A(n_279), .Y(n_283) );
OAI22x1_ASAP7_75t_L g285 ( .A1(n_279), .A2(n_286), .B1(n_287), .B2(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_279), .Y(n_286) );
INVx1_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
INVxp67_ASAP7_75t_L g353 ( .A(n_281), .Y(n_353) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g301 ( .A(n_282), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g325 ( .A(n_284), .B(n_301), .Y(n_325) );
AND2x2_ASAP7_75t_L g341 ( .A(n_284), .B(n_320), .Y(n_341) );
AND2x4_ASAP7_75t_L g366 ( .A(n_284), .B(n_320), .Y(n_366) );
AND2x4_ASAP7_75t_L g370 ( .A(n_284), .B(n_301), .Y(n_370) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_289), .Y(n_284) );
INVx2_ASAP7_75t_L g295 ( .A(n_285), .Y(n_295) );
AND2x2_ASAP7_75t_L g329 ( .A(n_285), .B(n_290), .Y(n_329) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_285), .Y(n_337) );
AND2x4_ASAP7_75t_L g294 ( .A(n_289), .B(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_290), .B(n_295), .Y(n_303) );
BUFx2_ASAP7_75t_L g306 ( .A(n_290), .Y(n_306) );
BUFx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
BUFx3_ASAP7_75t_L g413 ( .A(n_293), .Y(n_413) );
BUFx2_ASAP7_75t_SL g516 ( .A(n_293), .Y(n_516) );
BUFx2_ASAP7_75t_SL g733 ( .A(n_293), .Y(n_733) );
AND2x4_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
AND2x4_ASAP7_75t_L g313 ( .A(n_294), .B(n_301), .Y(n_313) );
AND2x4_ASAP7_75t_L g319 ( .A(n_294), .B(n_320), .Y(n_319) );
AND2x6_ASAP7_75t_L g382 ( .A(n_294), .B(n_301), .Y(n_382) );
AND2x4_ASAP7_75t_L g386 ( .A(n_294), .B(n_296), .Y(n_386) );
AND2x2_ASAP7_75t_L g389 ( .A(n_294), .B(n_320), .Y(n_389) );
AND2x4_ASAP7_75t_L g305 ( .A(n_296), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g336 ( .A(n_296), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_296), .B(n_337), .Y(n_367) );
AND2x4_ASAP7_75t_L g379 ( .A(n_296), .B(n_306), .Y(n_379) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_296), .B(n_337), .Y(n_424) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx3_ASAP7_75t_L g406 ( .A(n_300), .Y(n_406) );
INVx2_ASAP7_75t_L g521 ( .A(n_300), .Y(n_521) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_301), .B(n_303), .Y(n_378) );
AND2x2_ASAP7_75t_L g672 ( .A(n_301), .B(n_303), .Y(n_672) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_302), .Y(n_331) );
AND2x4_ASAP7_75t_L g349 ( .A(n_303), .B(n_320), .Y(n_349) );
AND2x2_ASAP7_75t_L g373 ( .A(n_303), .B(n_320), .Y(n_373) );
AND2x2_ASAP7_75t_L g575 ( .A(n_303), .B(n_320), .Y(n_575) );
BUFx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx3_ASAP7_75t_L g407 ( .A(n_305), .Y(n_407) );
BUFx2_ASAP7_75t_L g484 ( .A(n_305), .Y(n_484) );
INVx5_ASAP7_75t_SL g524 ( .A(n_305), .Y(n_524) );
INVx3_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g415 ( .A(n_309), .Y(n_415) );
INVx3_ASAP7_75t_L g433 ( .A(n_309), .Y(n_433) );
INVx2_ASAP7_75t_SL g481 ( .A(n_309), .Y(n_481) );
INVx4_ASAP7_75t_L g736 ( .A(n_309), .Y(n_736) );
INVx8_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_SL g411 ( .A(n_312), .Y(n_411) );
INVx2_ASAP7_75t_L g482 ( .A(n_312), .Y(n_482) );
INVx2_ASAP7_75t_L g508 ( .A(n_312), .Y(n_508) );
INVx2_ASAP7_75t_L g619 ( .A(n_312), .Y(n_619) );
INVx8_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx3_ASAP7_75t_L g410 ( .A(n_316), .Y(n_410) );
BUFx2_ASAP7_75t_L g504 ( .A(n_316), .Y(n_504) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g438 ( .A(n_319), .Y(n_438) );
BUFx3_ASAP7_75t_L g514 ( .A(n_319), .Y(n_514) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_319), .Y(n_675) );
NAND4xp25_ASAP7_75t_L g321 ( .A(n_322), .B(n_332), .C(n_342), .D(n_347), .Y(n_321) );
BUFx6f_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g570 ( .A(n_324), .Y(n_570) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_325), .Y(n_402) );
INVx3_ASAP7_75t_L g469 ( .A(n_325), .Y(n_469) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx2_ASAP7_75t_L g656 ( .A(n_327), .Y(n_656) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx3_ASAP7_75t_L g403 ( .A(n_328), .Y(n_403) );
BUFx4f_ASAP7_75t_L g470 ( .A(n_328), .Y(n_470) );
INVx1_ASAP7_75t_L g537 ( .A(n_328), .Y(n_537) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AND2x4_ASAP7_75t_L g352 ( .A(n_329), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_330), .Y(n_371) );
AND2x2_ASAP7_75t_L g374 ( .A(n_329), .B(n_353), .Y(n_374) );
AND2x2_ASAP7_75t_L g428 ( .A(n_329), .B(n_353), .Y(n_428) );
AND2x2_ASAP7_75t_L g666 ( .A(n_329), .B(n_330), .Y(n_666) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OAI222xp33_ASAP7_75t_L g526 ( .A1(n_334), .A2(n_527), .B1(n_528), .B2(n_531), .C1(n_532), .C2(n_533), .Y(n_526) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
BUFx12f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx3_ASAP7_75t_L g400 ( .A(n_336), .Y(n_400) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g532 ( .A(n_339), .Y(n_532) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g548 ( .A(n_340), .Y(n_548) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx5_ASAP7_75t_L g475 ( .A(n_341), .Y(n_475) );
BUFx3_ASAP7_75t_L g652 ( .A(n_341), .Y(n_652) );
BUFx3_ASAP7_75t_L g721 ( .A(n_341), .Y(n_721) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx4_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
INVx4_ASAP7_75t_SL g478 ( .A(n_345), .Y(n_478) );
INVx3_ASAP7_75t_SL g530 ( .A(n_345), .Y(n_530) );
BUFx2_ASAP7_75t_L g691 ( .A(n_345), .Y(n_691) );
INVx6_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx2_ASAP7_75t_L g539 ( .A(n_348), .Y(n_539) );
BUFx2_ASAP7_75t_L g724 ( .A(n_348), .Y(n_724) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
BUFx2_ASAP7_75t_L g472 ( .A(n_349), .Y(n_472) );
BUFx3_ASAP7_75t_L g550 ( .A(n_349), .Y(n_550) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
INVx2_ASAP7_75t_L g473 ( .A(n_351), .Y(n_473) );
INVx2_ASAP7_75t_L g540 ( .A(n_351), .Y(n_540) );
INVx6_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AOI22xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_441), .B1(n_442), .B2(n_492), .Y(n_355) );
AO22x1_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_417), .B1(n_418), .B2(n_440), .Y(n_356) );
INVx2_ASAP7_75t_L g440 ( .A(n_357), .Y(n_440) );
AO22x2_ASAP7_75t_L g493 ( .A1(n_357), .A2(n_417), .B1(n_418), .B2(n_440), .Y(n_493) );
XOR2x1_ASAP7_75t_SL g357 ( .A(n_358), .B(n_390), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_360), .B(n_375), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_361), .B(n_368), .Y(n_360) );
OAI21xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_364), .B(n_365), .Y(n_361) );
INVx2_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g567 ( .A(n_363), .Y(n_567) );
INVx1_ASAP7_75t_SL g629 ( .A(n_366), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_372), .Y(n_368) );
INVxp67_ASAP7_75t_L g577 ( .A(n_374), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_383), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_380), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_384), .B(n_387), .Y(n_383) );
XNOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_416), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_404), .Y(n_391) );
NAND4xp25_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .C(n_398), .D(n_401), .Y(n_392) );
BUFx2_ASAP7_75t_L g650 ( .A(n_399), .Y(n_650) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g476 ( .A(n_400), .Y(n_476) );
INVx3_ASAP7_75t_L g694 ( .A(n_400), .Y(n_694) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .C(n_412), .D(n_414), .Y(n_404) );
INVx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g486 ( .A(n_410), .Y(n_486) );
INVx2_ASAP7_75t_SL g731 ( .A(n_410), .Y(n_731) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_413), .Y(n_646) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
XOR2x2_ASAP7_75t_L g418 ( .A(n_419), .B(n_439), .Y(n_418) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_420), .B(n_429), .Y(n_419) );
NOR2x1_ASAP7_75t_L g420 ( .A(n_421), .B(n_425), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_434), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_461), .B1(n_462), .B2(n_491), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g459 ( .A(n_446), .Y(n_459) );
NAND2x1_ASAP7_75t_SL g446 ( .A(n_447), .B(n_452), .Y(n_446) );
NOR2xp67_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
NOR2x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_479), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_471), .C(n_474), .D(n_477), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx4_ASAP7_75t_L g626 ( .A(n_469), .Y(n_626) );
NAND4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_483), .C(n_485), .D(n_488), .Y(n_479) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_487), .Y(n_640) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
XNOR2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_590), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_541), .B1(n_542), .B2(n_588), .Y(n_497) );
INVxp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g589 ( .A(n_499), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_515), .C(n_525), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_509), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_502) );
INVx2_ASAP7_75t_L g682 ( .A(n_503), .Y(n_682) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_517) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_520), .Y(n_729) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g608 ( .A(n_521), .Y(n_608) );
INVx1_ASAP7_75t_L g643 ( .A(n_521), .Y(n_643) );
INVx2_ASAP7_75t_L g556 ( .A(n_524), .Y(n_556) );
INVx3_ASAP7_75t_L g609 ( .A(n_524), .Y(n_609) );
INVx2_ASAP7_75t_L g644 ( .A(n_524), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_534), .Y(n_525) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_537), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_568) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AO22x2_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_560), .B2(n_587), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_553), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_549), .C(n_551), .D(n_552), .Y(n_546) );
NAND4xp25_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .C(n_557), .D(n_559), .Y(n_553) );
INVx2_ASAP7_75t_L g587 ( .A(n_560), .Y(n_587) );
INVx1_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_578), .Y(n_562) );
NOR3xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .C(n_572), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_565), .B(n_566), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_574), .B1(n_576), .B2(n_577), .Y(n_572) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OAI22xp5_ASAP7_75t_SL g590 ( .A1(n_591), .A2(n_592), .B1(n_659), .B2(n_700), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_635), .B2(n_658), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22x1_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B1(n_613), .B2(n_631), .Y(n_595) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_605), .Y(n_599) );
NAND4xp25_ASAP7_75t_SL g600 ( .A(n_601), .B(n_602), .C(n_603), .D(n_604), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .C(n_610), .D(n_611), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_614), .Y(n_634) );
INVx1_ASAP7_75t_L g630 ( .A(n_615), .Y(n_630) );
NOR2x1_ASAP7_75t_SL g633 ( .A(n_615), .B(n_634), .Y(n_633) );
NAND4xp75_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .C(n_623), .D(n_627), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
AND2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_631), .A2(n_660), .B1(n_698), .B2(n_699), .Y(n_659) );
INVx3_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_632), .Y(n_699) );
INVx2_ASAP7_75t_L g658 ( .A(n_635), .Y(n_658) );
XNOR2x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_657), .Y(n_635) );
NOR2xp67_ASAP7_75t_L g636 ( .A(n_637), .B(n_647), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .C(n_641), .D(n_645), .Y(n_637) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND4xp25_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .C(n_653), .D(n_654), .Y(n_647) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g700 ( .A(n_659), .Y(n_700) );
INVx1_ASAP7_75t_L g698 ( .A(n_660), .Y(n_698) );
XOR2x1_ASAP7_75t_L g660 ( .A(n_661), .B(n_678), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
XNOR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_677), .Y(n_662) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_664), .B(n_670), .Y(n_663) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .C(n_668), .D(n_669), .Y(n_664) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .C(n_674), .D(n_676), .Y(n_670) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_675), .Y(n_685) );
XOR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_697), .Y(n_678) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_688), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .C(n_684), .D(n_686), .Y(n_680) );
NAND4xp25_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .C(n_695), .D(n_696), .Y(n_688) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_706), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_704), .B(n_707), .Y(n_743) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
OAI222xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_738), .B1(n_740), .B2(n_741), .C1(n_744), .C2(n_745), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_725), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .C(n_722), .D(n_723), .Y(n_716) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_726), .B(n_728), .C(n_730), .D(n_732), .Y(n_725) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
CKINVDCx6p67_ASAP7_75t_R g742 ( .A(n_743), .Y(n_742) );
endmodule