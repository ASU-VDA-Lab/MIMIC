module fake_jpeg_7210_n_256 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_256);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_34),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_17),
.B(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_13),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_35),
.A2(n_26),
.B1(n_17),
.B2(n_19),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_47),
.B1(n_16),
.B2(n_25),
.Y(n_70)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_26),
.B1(n_13),
.B2(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_24),
.B1(n_15),
.B2(n_18),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_54),
.B1(n_31),
.B2(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_31),
.A2(n_29),
.B1(n_23),
.B2(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_82)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_28),
.C(n_36),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_59),
.C(n_16),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_28),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_37),
.B1(n_36),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_52),
.B1(n_41),
.B2(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_42),
.Y(n_81)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_67),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_50),
.B1(n_20),
.B2(n_25),
.Y(n_92)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_72),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_76),
.A2(n_82),
.B1(n_60),
.B2(n_65),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_43),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_84),
.C(n_20),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_57),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_44),
.A3(n_36),
.B1(n_37),
.B2(n_30),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_63),
.B(n_66),
.C(n_30),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_65),
.B1(n_69),
.B2(n_67),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_56),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_95),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_101),
.B(n_102),
.Y(n_114)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_106),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_84),
.A2(n_59),
.B(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_103),
.A2(n_109),
.B1(n_77),
.B2(n_74),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_104),
.A2(n_108),
.B1(n_111),
.B2(n_99),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_113),
.B1(n_77),
.B2(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_71),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_25),
.B(n_18),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_88),
.B(n_18),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_77),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.C(n_15),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_85),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_87),
.C(n_83),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_73),
.B1(n_63),
.B2(n_37),
.Y(n_113)
);

XOR2x2_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_86),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_116),
.B(n_119),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_78),
.B(n_75),
.C(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_121),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_111),
.A2(n_78),
.B1(n_75),
.B2(n_74),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_126),
.B1(n_130),
.B2(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_109),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_123),
.Y(n_137)
);

NOR2x1_ASAP7_75t_R g124 ( 
.A(n_98),
.B(n_20),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_107),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_133),
.B1(n_105),
.B2(n_101),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_91),
.B1(n_73),
.B2(n_30),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_131),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_15),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_132),
.C(n_102),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_89),
.B1(n_68),
.B2(n_36),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_155),
.B1(n_115),
.B2(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_142),
.A2(n_144),
.B(n_147),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_108),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_138),
.B(n_140),
.Y(n_170)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_148),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_132),
.C(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_156),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_99),
.B1(n_89),
.B2(n_97),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_27),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_32),
.B(n_27),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_128),
.B1(n_119),
.B2(n_114),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_162),
.C(n_165),
.Y(n_181)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_0),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_164),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_127),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_147),
.B1(n_137),
.B2(n_144),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_134),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_97),
.C(n_80),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_172),
.C(n_175),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_8),
.C(n_9),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_142),
.C(n_143),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_139),
.B(n_9),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_169),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_170),
.A2(n_27),
.B(n_21),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_32),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_151),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_27),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_178),
.B(n_182),
.CI(n_168),
.CON(n_194),
.SN(n_194)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_150),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_185),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_186),
.B1(n_191),
.B2(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_173),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_184),
.A2(n_192),
.B(n_161),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_142),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_172),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_177),
.Y(n_198)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_202),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_166),
.C(n_171),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_207),
.C(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_201),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_169),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_203),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_182),
.A2(n_170),
.B1(n_167),
.B2(n_175),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_204),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_32),
.C(n_21),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_178),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_208),
.Y(n_215)
);

FAx1_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_185),
.CI(n_187),
.CON(n_209),
.SN(n_209)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_209),
.A2(n_211),
.B(n_197),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_196),
.A2(n_187),
.B(n_189),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_212),
.A2(n_205),
.B1(n_204),
.B2(n_202),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_206),
.A2(n_21),
.B(n_6),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_195),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_210),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_6),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_231),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_194),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_225),
.B(n_227),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_200),
.C(n_207),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_232),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_229),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_230),
.A2(n_209),
.B1(n_211),
.B2(n_217),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_199),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_11),
.C(n_10),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_236),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_225),
.A2(n_217),
.B1(n_10),
.B2(n_7),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_1),
.C(n_2),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_7),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_0),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_240),
.B(n_1),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_243),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_237),
.A2(n_227),
.B(n_223),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_246),
.C(n_1),
.Y(n_247)
);

NOR2x1p5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_1),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_238),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_247),
.A2(n_248),
.B(n_241),
.C(n_4),
.Y(n_250)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_238),
.B(n_3),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_251),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_2),
.B(n_4),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_2),
.C(n_4),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_4),
.Y(n_256)
);


endmodule