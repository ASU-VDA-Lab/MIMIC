module fake_netlist_6_84_n_2184 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2184);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2184;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_137),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_19),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_185),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_49),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_141),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_6),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_71),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_142),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_117),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_190),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_77),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_199),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_83),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_69),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_79),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_105),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_79),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_145),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_27),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_88),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_64),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_180),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_187),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_72),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_168),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_11),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_186),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_208),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_71),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_94),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_84),
.Y(n_275)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_60),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_12),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_163),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_204),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_200),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_48),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_30),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_206),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_103),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_113),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_74),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_92),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_34),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_63),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_57),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_97),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_166),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_96),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_124),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_181),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_57),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_165),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_151),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_135),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_189),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_21),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_149),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_196),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_211),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_146),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_221),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_131),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_34),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_31),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_191),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_150),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_119),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_226),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_179),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_52),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_52),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_111),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_81),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_107),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_80),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_62),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_35),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_228),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_127),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_139),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_77),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_114),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_74),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_183),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_219),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_155),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_42),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_87),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_167),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_65),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_205),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_3),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_69),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_37),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_35),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_123),
.Y(n_344)
);

BUFx10_ASAP7_75t_L g345 ( 
.A(n_61),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_61),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_81),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_184),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_148),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_9),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_108),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_25),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_214),
.Y(n_353)
);

BUFx10_ASAP7_75t_L g354 ( 
.A(n_10),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_126),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_28),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_112),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_86),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_174),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_3),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_129),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_68),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_192),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_222),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g366 ( 
.A(n_201),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_116),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_156),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_2),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_216),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_33),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_73),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_59),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_121),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_202),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_209),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_133),
.Y(n_377)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_58),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_212),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_230),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_172),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_32),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_227),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_193),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_72),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_14),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_176),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_43),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_23),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_65),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_45),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_210),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_16),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_30),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_115),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_82),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_161),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_50),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_99),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_203),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_89),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_140),
.Y(n_402)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_160),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_218),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_25),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_55),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_18),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_32),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_53),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_58),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_85),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_17),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_169),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_47),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_31),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_164),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_173),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_24),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_78),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_26),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_122),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_18),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_80),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_170),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_39),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_91),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_134),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_11),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_59),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_157),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_93),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_217),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_56),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_60),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_22),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_0),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_224),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_2),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_175),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_215),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_46),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_110),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_144),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_13),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_29),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_104),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_62),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_147),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_49),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_43),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_28),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_197),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_1),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_188),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_319),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_280),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_281),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_326),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_292),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_336),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_292),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_365),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_292),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_379),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_404),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_436),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_329),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_358),
.B(n_0),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_292),
.Y(n_469)
);

BUFx2_ASAP7_75t_SL g470 ( 
.A(n_248),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_413),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_426),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_367),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_362),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_306),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_434),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_289),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_292),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_385),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_292),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_293),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_292),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_433),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_295),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_296),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_301),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_302),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_438),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_252),
.B(n_1),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_305),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_265),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_272),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_282),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_303),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_443),
.B(n_4),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_292),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_321),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g500 ( 
.A(n_235),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_308),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_378),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_325),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_310),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_378),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_244),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_378),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_378),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_378),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_340),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_313),
.Y(n_511)
);

INVxp33_ASAP7_75t_SL g512 ( 
.A(n_235),
.Y(n_512)
);

INVxp67_ASAP7_75t_SL g513 ( 
.A(n_265),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_341),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_346),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_378),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_369),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_378),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_248),
.B(n_4),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_257),
.B(n_5),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_244),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_315),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_371),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_R g524 ( 
.A(n_276),
.B(n_5),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_242),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_241),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_345),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_242),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_372),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_373),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_R g531 ( 
.A(n_276),
.B(n_6),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_316),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_242),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_242),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_242),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_382),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_386),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_312),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_312),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_312),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_312),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_333),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_388),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_312),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_331),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_389),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_275),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_331),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_331),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_391),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_331),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_331),
.Y(n_552)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_254),
.B(n_7),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_276),
.B(n_8),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_420),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_420),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_393),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_394),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_420),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_420),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_256),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_345),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_264),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_453),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_345),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_267),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_277),
.B(n_8),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_278),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g570 ( 
.A(n_354),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_334),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_354),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_337),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_339),
.Y(n_574)
);

INVxp33_ASAP7_75t_SL g575 ( 
.A(n_238),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_255),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_538),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_456),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_513),
.B(n_547),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_533),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_477),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_533),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_538),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_539),
.B(n_275),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_539),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_481),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_484),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_485),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_483),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_491),
.B(n_255),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_457),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_548),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_486),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_555),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_458),
.Y(n_597)
);

INVx6_ASAP7_75t_L g598 ( 
.A(n_491),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_488),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_525),
.Y(n_601)
);

AOI22x1_ASAP7_75t_SL g602 ( 
.A1(n_460),
.A2(n_338),
.B1(n_343),
.B2(n_273),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_528),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_470),
.B(n_554),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_534),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_487),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_490),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_535),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_540),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_501),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_470),
.B(n_368),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_544),
.Y(n_613)
);

BUFx8_ASAP7_75t_L g614 ( 
.A(n_466),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_545),
.B(n_368),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_549),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_488),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_459),
.B(n_232),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_504),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_551),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_552),
.B(n_397),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_462),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_556),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_560),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_521),
.B(n_397),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_561),
.B(n_249),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_511),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_482),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_522),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_461),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_532),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_463),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_455),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_506),
.B(n_283),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_467),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_482),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_497),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_542),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_506),
.B(n_249),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_571),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_469),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_478),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_497),
.B(n_268),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_562),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_480),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_573),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_496),
.B(n_268),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_502),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_505),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_507),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_507),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_474),
.B(n_266),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_508),
.Y(n_654)
);

INVx6_ASAP7_75t_L g655 ( 
.A(n_553),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_574),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_509),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_516),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_518),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_519),
.B(n_411),
.Y(n_660)
);

CKINVDCx20_ASAP7_75t_R g661 ( 
.A(n_464),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_493),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_576),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_553),
.A2(n_320),
.B(n_279),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_465),
.Y(n_666)
);

CKINVDCx20_ASAP7_75t_R g667 ( 
.A(n_471),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_564),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_472),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_493),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_568),
.Y(n_671)
);

INVx4_ASAP7_75t_SL g672 ( 
.A(n_660),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_645),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_655),
.A2(n_495),
.B1(n_489),
.B2(n_468),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_604),
.B(n_279),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_631),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_578),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_584),
.B(n_567),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_631),
.Y(n_679)
);

INVx6_ASAP7_75t_L g680 ( 
.A(n_598),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_579),
.B(n_474),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_585),
.B(n_563),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_660),
.B(n_476),
.Y(n_683)
);

INVx5_ASAP7_75t_L g684 ( 
.A(n_660),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_633),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_654),
.Y(n_686)
);

INVx5_ASAP7_75t_L g687 ( 
.A(n_660),
.Y(n_687)
);

INVxp33_ASAP7_75t_L g688 ( 
.A(n_634),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_633),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_660),
.A2(n_671),
.B1(n_568),
.B2(n_655),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_660),
.A2(n_283),
.B1(n_520),
.B2(n_359),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_577),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_577),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_653),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_642),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_671),
.B(n_500),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_585),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_642),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_660),
.B(n_476),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_643),
.B(n_494),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_654),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_598),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_671),
.B(n_500),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_643),
.Y(n_704)
);

OR2x6_ASAP7_75t_L g705 ( 
.A(n_617),
.B(n_572),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_598),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_598),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_636),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_662),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_655),
.A2(n_359),
.B1(n_364),
.B2(n_320),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_584),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_646),
.B(n_494),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_646),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_649),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_649),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_650),
.B(n_499),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_583),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_612),
.B(n_479),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_637),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_593),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_650),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_644),
.B(n_364),
.Y(n_723)
);

INVx4_ASAP7_75t_L g724 ( 
.A(n_654),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_637),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_655),
.B(n_512),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_584),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_652),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_635),
.B(n_499),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_658),
.B(n_659),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_640),
.B(n_510),
.C(n_503),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_665),
.A2(n_416),
.B1(n_421),
.B2(n_399),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_657),
.Y(n_735)
);

AND2x4_ASAP7_75t_L g736 ( 
.A(n_584),
.B(n_569),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_615),
.B(n_503),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_665),
.A2(n_416),
.B1(n_421),
.B2(n_399),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_657),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_668),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_644),
.A2(n_446),
.B1(n_291),
.B2(n_298),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_652),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_668),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_654),
.Y(n_744)
);

OAI22xp33_ASAP7_75t_L g745 ( 
.A1(n_626),
.A2(n_531),
.B1(n_524),
.B2(n_347),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_615),
.B(n_510),
.Y(n_746)
);

AND3x2_ASAP7_75t_L g747 ( 
.A(n_617),
.B(n_466),
.C(n_446),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_654),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_615),
.B(n_512),
.Y(n_749)
);

BUFx4f_ASAP7_75t_L g750 ( 
.A(n_592),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_654),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_615),
.B(n_514),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_644),
.B(n_411),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_644),
.A2(n_311),
.B1(n_318),
.B2(n_287),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_621),
.B(n_411),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_629),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_635),
.B(n_514),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_629),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_629),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_621),
.B(n_515),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_610),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_638),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_601),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_638),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_603),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_603),
.Y(n_766)
);

OR2x6_ASAP7_75t_L g767 ( 
.A(n_591),
.B(n_498),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_621),
.B(n_515),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_621),
.B(n_575),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_638),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_610),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_618),
.B(n_517),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_605),
.B(n_575),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_618),
.B(n_411),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_638),
.B(n_651),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_627),
.B(n_411),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_600),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_605),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_608),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_608),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_651),
.B(n_517),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_609),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_R g783 ( 
.A(n_581),
.B(n_523),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_651),
.B(n_523),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_592),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_609),
.Y(n_786)
);

INVx4_ASAP7_75t_SL g787 ( 
.A(n_627),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_613),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_670),
.B(n_529),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_613),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_651),
.B(n_529),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_627),
.B(n_239),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_587),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_616),
.Y(n_794)
);

INVx5_ASAP7_75t_L g795 ( 
.A(n_627),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_616),
.Y(n_796)
);

OR2x6_ASAP7_75t_L g797 ( 
.A(n_614),
.B(n_323),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_623),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_623),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_620),
.B(n_530),
.Y(n_800)
);

AND2x2_ASAP7_75t_SL g801 ( 
.A(n_648),
.B(n_442),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_614),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_580),
.B(n_530),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_614),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_625),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_620),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_624),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_625),
.Y(n_808)
);

BUFx8_ASAP7_75t_SL g809 ( 
.A(n_597),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_586),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_622),
.Y(n_811)
);

INVx8_ASAP7_75t_L g812 ( 
.A(n_588),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_624),
.B(n_536),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_580),
.Y(n_814)
);

OAI22xp33_ASAP7_75t_L g815 ( 
.A1(n_664),
.A2(n_290),
.B1(n_526),
.B2(n_527),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_586),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_614),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_661),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_582),
.B(n_536),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_582),
.B(n_537),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_664),
.A2(n_324),
.B1(n_342),
.B2(n_335),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_663),
.B(n_537),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_663),
.B(n_543),
.Y(n_823)
);

INVxp33_ASAP7_75t_L g824 ( 
.A(n_589),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_602),
.A2(n_473),
.B1(n_356),
.B2(n_441),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_589),
.B(n_442),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_594),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_594),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_596),
.B(n_543),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_801),
.B(n_546),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_690),
.B(n_442),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_785),
.B(n_546),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_801),
.B(n_550),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_711),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_690),
.B(n_550),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_694),
.B(n_557),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_720),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_681),
.B(n_475),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_684),
.B(n_442),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_727),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_676),
.B(n_558),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_684),
.B(n_442),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_679),
.B(n_558),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_727),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_720),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_708),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_685),
.B(n_565),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_684),
.B(n_448),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_696),
.B(n_565),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_702),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_725),
.Y(n_851)
);

OAI22xp33_ASAP7_75t_L g852 ( 
.A1(n_674),
.A2(n_570),
.B1(n_566),
.B2(n_300),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_696),
.A2(n_309),
.B1(n_366),
.B2(n_307),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_740),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_703),
.B(n_590),
.Y(n_855)
);

NAND2x1_ASAP7_75t_L g856 ( 
.A(n_756),
.B(n_596),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_743),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_689),
.B(n_243),
.Y(n_858)
);

NAND2xp33_ASAP7_75t_L g859 ( 
.A(n_691),
.B(n_448),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_695),
.B(n_250),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_785),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_698),
.B(n_263),
.Y(n_862)
);

INVxp33_ASAP7_75t_L g863 ( 
.A(n_773),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_703),
.A2(n_403),
.B1(n_344),
.B2(n_348),
.Y(n_864)
);

NAND2xp33_ASAP7_75t_L g865 ( 
.A(n_691),
.B(n_448),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_704),
.B(n_284),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_714),
.B(n_285),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_700),
.B(n_595),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_763),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_713),
.B(n_606),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_684),
.B(n_448),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_702),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_765),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_766),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_715),
.B(n_286),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_750),
.A2(n_297),
.B1(n_353),
.B2(n_351),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_687),
.B(n_448),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_716),
.B(n_722),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_750),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_730),
.B(n_288),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_725),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_675),
.A2(n_290),
.B1(n_431),
.B2(n_381),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_822),
.Y(n_883)
);

OR2x2_ASAP7_75t_L g884 ( 
.A(n_697),
.B(n_607),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_710),
.A2(n_349),
.B1(n_328),
.B2(n_322),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_734),
.B(n_294),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_717),
.B(n_611),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_687),
.B(n_299),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_L g889 ( 
.A(n_733),
.B(n_304),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_814),
.B(n_314),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_709),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_728),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_742),
.Y(n_893)
);

NOR2xp67_ASAP7_75t_SL g894 ( 
.A(n_687),
.B(n_317),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_729),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_731),
.B(n_363),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_742),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_778),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_823),
.B(n_383),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_757),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_823),
.B(n_427),
.Y(n_901)
);

INVx8_ASAP7_75t_L g902 ( 
.A(n_675),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_810),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_726),
.B(n_732),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_810),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_773),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_812),
.B(n_452),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_706),
.Y(n_908)
);

AO22x1_ASAP7_75t_L g909 ( 
.A1(n_726),
.A2(n_259),
.B1(n_269),
.B2(n_261),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_688),
.B(n_619),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_816),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_779),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_688),
.B(n_781),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_749),
.A2(n_414),
.B(n_422),
.C(n_425),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_687),
.B(n_454),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_675),
.A2(n_398),
.B1(n_350),
.B2(n_352),
.Y(n_916)
);

AND2x4_ASAP7_75t_SL g917 ( 
.A(n_709),
.B(n_666),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_784),
.B(n_628),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_733),
.B(n_355),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_710),
.B(n_599),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_738),
.B(n_599),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_738),
.B(n_357),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_820),
.B(n_361),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_802),
.B(n_630),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_791),
.B(n_632),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_816),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_820),
.B(n_370),
.Y(n_927)
);

NOR2xp67_ASAP7_75t_SL g928 ( 
.A(n_683),
.B(n_360),
.Y(n_928)
);

AO22x1_ASAP7_75t_L g929 ( 
.A1(n_749),
.A2(n_238),
.B1(n_246),
.B2(n_251),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_675),
.A2(n_429),
.B1(n_408),
.B2(n_447),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_678),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_737),
.B(n_639),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_780),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_756),
.B(n_829),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_756),
.B(n_374),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_746),
.B(n_641),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_789),
.B(n_647),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_678),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_829),
.B(n_375),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_782),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_752),
.B(n_656),
.Y(n_941)
);

NAND2x1_ASAP7_75t_L g942 ( 
.A(n_712),
.B(n_390),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_719),
.B(n_246),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_786),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_788),
.B(n_376),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_790),
.B(n_377),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_794),
.B(n_380),
.Y(n_947)
);

OR2x2_ASAP7_75t_L g948 ( 
.A(n_767),
.B(n_251),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_796),
.B(n_384),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_806),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_692),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_800),
.B(n_354),
.Y(n_952)
);

NAND2xp33_ASAP7_75t_L g953 ( 
.A(n_675),
.B(n_233),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_792),
.A2(n_405),
.B1(n_449),
.B2(n_451),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_807),
.B(n_387),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_813),
.B(n_392),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_769),
.A2(n_395),
.B1(n_396),
.B2(n_233),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_692),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_760),
.B(n_768),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_813),
.B(n_234),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_R g961 ( 
.A(n_783),
.B(n_667),
.Y(n_961)
);

NOR3xp33_ASAP7_75t_L g962 ( 
.A(n_815),
.B(n_259),
.C(n_261),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_678),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_L g964 ( 
.A(n_741),
.B(n_234),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_769),
.B(n_450),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_693),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_709),
.B(n_450),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_712),
.B(n_236),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_809),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_736),
.Y(n_970)
);

INVxp67_ASAP7_75t_L g971 ( 
.A(n_783),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_L g972 ( 
.A1(n_792),
.A2(n_406),
.B1(n_419),
.B2(n_444),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_736),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_758),
.B(n_236),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_792),
.A2(n_406),
.B1(n_419),
.B2(n_444),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_758),
.B(n_237),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_745),
.B(n_237),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_693),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_767),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_723),
.A2(n_269),
.B1(n_423),
.B2(n_418),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_706),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_759),
.B(n_240),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_701),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_672),
.B(n_240),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_736),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_723),
.A2(n_409),
.B(n_445),
.C(n_428),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_759),
.B(n_245),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_803),
.A2(n_402),
.B1(n_247),
.B2(n_440),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_762),
.B(n_245),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_762),
.B(n_247),
.Y(n_990)
);

O2A1O1Ixp5_ASAP7_75t_L g991 ( 
.A1(n_755),
.A2(n_258),
.B(n_440),
.C(n_439),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_819),
.B(n_669),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_741),
.A2(n_435),
.B(n_423),
.C(n_418),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_735),
.A2(n_435),
.B1(n_415),
.B2(n_412),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_934),
.A2(n_921),
.B(n_831),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_959),
.A2(n_699),
.B(n_673),
.C(n_772),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_904),
.B(n_777),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_856),
.A2(n_748),
.B(n_744),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_952),
.A2(n_863),
.B(n_849),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_850),
.Y(n_1000)
);

OAI321xp33_ASAP7_75t_L g1001 ( 
.A1(n_906),
.A2(n_821),
.A3(n_754),
.B1(n_797),
.B2(n_682),
.C(n_705),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_850),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_883),
.A2(n_707),
.B1(n_680),
.B2(n_739),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_831),
.A2(n_724),
.B(n_686),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_863),
.B(n_682),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_883),
.A2(n_680),
.B1(n_751),
.B2(n_828),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_923),
.B(n_824),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_927),
.B(n_824),
.Y(n_1008)
);

INVx11_ASAP7_75t_L g1009 ( 
.A(n_961),
.Y(n_1009)
);

OAI321xp33_ASAP7_75t_L g1010 ( 
.A1(n_852),
.A2(n_977),
.A3(n_960),
.B1(n_835),
.B2(n_914),
.C(n_901),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_895),
.B(n_879),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_879),
.A2(n_724),
.B(n_686),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_830),
.A2(n_754),
.B1(n_680),
.B2(n_804),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_939),
.B(n_770),
.Y(n_1014)
);

AO21x1_ASAP7_75t_L g1015 ( 
.A1(n_859),
.A2(n_755),
.B(n_753),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_836),
.B(n_811),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_935),
.A2(n_724),
.B(n_686),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_850),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_889),
.A2(n_795),
.B(n_775),
.Y(n_1019)
);

CKINVDCx10_ASAP7_75t_R g1020 ( 
.A(n_891),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_956),
.B(n_770),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_900),
.B(n_705),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_832),
.B(n_705),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_889),
.A2(n_753),
.B(n_776),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_859),
.A2(n_795),
.B(n_701),
.Y(n_1025)
);

AND2x2_ASAP7_75t_SL g1026 ( 
.A(n_917),
.B(n_817),
.Y(n_1026)
);

AOI21x1_ASAP7_75t_L g1027 ( 
.A1(n_928),
.A2(n_774),
.B(n_776),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_895),
.B(n_777),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_899),
.B(n_827),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_961),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_913),
.B(n_761),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_833),
.B(n_793),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_846),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_854),
.B(n_761),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_837),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_865),
.A2(n_795),
.B(n_701),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_937),
.B(n_793),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_986),
.A2(n_821),
.B(n_805),
.C(n_798),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_857),
.B(n_771),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_865),
.A2(n_795),
.B(n_701),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_855),
.B(n_818),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_931),
.A2(n_764),
.B(n_774),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_920),
.A2(n_718),
.B(n_808),
.Y(n_1043)
);

INVxp67_ASAP7_75t_SL g1044 ( 
.A(n_850),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_977),
.A2(n_798),
.B(n_808),
.C(n_805),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_853),
.A2(n_718),
.B(n_825),
.C(n_253),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_882),
.A2(n_415),
.B1(n_412),
.B2(n_410),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_905),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_971),
.B(n_677),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_872),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_L g1051 ( 
.A(n_907),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_931),
.A2(n_963),
.B(n_938),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_869),
.B(n_799),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_938),
.B(n_787),
.Y(n_1054)
);

BUFx8_ASAP7_75t_SL g1055 ( 
.A(n_969),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_963),
.A2(n_764),
.B(n_799),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_888),
.A2(n_787),
.B(n_672),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_973),
.A2(n_764),
.B(n_799),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_973),
.A2(n_764),
.B(n_799),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_838),
.A2(n_787),
.B1(n_797),
.B2(n_253),
.Y(n_1060)
);

AOI21x1_ASAP7_75t_L g1061 ( 
.A1(n_888),
.A2(n_672),
.B(n_797),
.Y(n_1061)
);

OA22x2_ASAP7_75t_L g1062 ( 
.A1(n_861),
.A2(n_747),
.B1(n_410),
.B2(n_602),
.Y(n_1062)
);

NAND3x1_ASAP7_75t_L g1063 ( 
.A(n_962),
.B(n_992),
.C(n_910),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_878),
.A2(n_826),
.B(n_401),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_905),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_914),
.A2(n_826),
.B(n_721),
.C(n_677),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_993),
.A2(n_972),
.B1(n_975),
.B2(n_954),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_919),
.A2(n_260),
.B(n_262),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_873),
.B(n_260),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_919),
.A2(n_401),
.B(n_270),
.Y(n_1070)
);

AOI22x1_ASAP7_75t_L g1071 ( 
.A1(n_834),
.A2(n_262),
.B1(n_439),
.B2(n_437),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_965),
.A2(n_402),
.B(n_271),
.C(n_437),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_868),
.B(n_721),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_922),
.A2(n_332),
.B(n_432),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_969),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_922),
.A2(n_991),
.B(n_926),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_970),
.B(n_270),
.Y(n_1077)
);

AO22x1_ASAP7_75t_L g1078 ( 
.A1(n_967),
.A2(n_400),
.B1(n_432),
.B2(n_430),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_872),
.Y(n_1079)
);

NAND2xp33_ASAP7_75t_L g1080 ( 
.A(n_902),
.B(n_812),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_908),
.Y(n_1081)
);

OAI22x1_ASAP7_75t_L g1082 ( 
.A1(n_979),
.A2(n_809),
.B1(n_812),
.B2(n_430),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_874),
.B(n_271),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_837),
.A2(n_153),
.B(n_95),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_983),
.A2(n_332),
.B(n_424),
.Y(n_1085)
);

BUFx8_ASAP7_75t_L g1086 ( 
.A(n_891),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_891),
.B(n_812),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_915),
.A2(n_424),
.B(n_417),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_898),
.B(n_274),
.Y(n_1089)
);

OAI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_911),
.A2(n_926),
.B(n_896),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_912),
.B(n_274),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_911),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_968),
.A2(n_330),
.B(n_327),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_933),
.B(n_9),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_940),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_974),
.A2(n_231),
.B(n_194),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_988),
.B(n_12),
.C(n_13),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_908),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_976),
.A2(n_182),
.B(n_178),
.Y(n_1099)
);

OR2x6_ASAP7_75t_L g1100 ( 
.A(n_884),
.B(n_14),
.Y(n_1100)
);

AO21x1_ASAP7_75t_L g1101 ( 
.A1(n_876),
.A2(n_15),
.B(n_16),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_982),
.A2(n_171),
.B(n_162),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_981),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_SL g1104 ( 
.A(n_918),
.B(n_159),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_915),
.A2(n_154),
.B(n_152),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_993),
.A2(n_15),
.B(n_17),
.C(n_19),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_845),
.A2(n_143),
.B(n_136),
.Y(n_1107)
);

OAI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_845),
.A2(n_132),
.B(n_130),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_870),
.B(n_20),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_987),
.A2(n_128),
.B(n_125),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_851),
.A2(n_118),
.B(n_106),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_989),
.A2(n_102),
.B(n_101),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_916),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_917),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_990),
.A2(n_100),
.B(n_98),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_L g1116 ( 
.A(n_864),
.B(n_24),
.C(n_26),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_851),
.A2(n_90),
.B(n_29),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_981),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_945),
.A2(n_27),
.B(n_33),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_887),
.B(n_78),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_944),
.B(n_36),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_SL g1122 ( 
.A(n_925),
.B(n_36),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_950),
.B(n_37),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_946),
.A2(n_38),
.B(n_39),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_947),
.A2(n_38),
.B(n_40),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_949),
.A2(n_40),
.B(n_41),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_890),
.B(n_41),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_964),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_840),
.B(n_44),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_943),
.B(n_76),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_955),
.A2(n_47),
.B(n_48),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_839),
.A2(n_50),
.B(n_51),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_844),
.A2(n_51),
.B(n_53),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_942),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_841),
.B(n_54),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_985),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_881),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_843),
.A2(n_54),
.B(n_55),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_847),
.B(n_56),
.Y(n_1139)
);

NAND3xp33_ASAP7_75t_SL g1140 ( 
.A(n_957),
.B(n_63),
.C(n_64),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_984),
.A2(n_66),
.B(n_67),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_932),
.B(n_66),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_964),
.A2(n_67),
.B(n_68),
.C(n_70),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_902),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_881),
.A2(n_70),
.B(n_73),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_984),
.A2(n_897),
.B(n_978),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_936),
.B(n_75),
.Y(n_1147)
);

AND2x2_ASAP7_75t_SL g1148 ( 
.A(n_941),
.B(n_75),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_902),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_924),
.B(n_862),
.Y(n_1150)
);

OAI321xp33_ASAP7_75t_L g1151 ( 
.A1(n_885),
.A2(n_980),
.A3(n_994),
.B1(n_930),
.B2(n_948),
.C(n_860),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_858),
.A2(n_886),
.B1(n_866),
.B2(n_867),
.Y(n_1152)
);

O2A1O1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_953),
.A2(n_875),
.B(n_880),
.C(n_966),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_892),
.B(n_978),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_893),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_893),
.B(n_966),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_953),
.A2(n_907),
.B1(n_958),
.B2(n_951),
.Y(n_1157)
);

OAI21xp33_ASAP7_75t_L g1158 ( 
.A1(n_907),
.A2(n_909),
.B(n_929),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_SL g1159 ( 
.A(n_839),
.B(n_842),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_842),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_902),
.B(n_848),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_848),
.A2(n_871),
.B(n_877),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_871),
.B(n_877),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_907),
.A2(n_831),
.B(n_921),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_894),
.B(n_694),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_831),
.A2(n_921),
.B(n_835),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_961),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_906),
.B(n_694),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_934),
.A2(n_750),
.B(n_921),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_835),
.A2(n_690),
.B1(n_934),
.B2(n_906),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_850),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_959),
.B(n_849),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_903),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_934),
.A2(n_750),
.B(n_921),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_995),
.A2(n_1166),
.B(n_1170),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1008),
.B(n_1031),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1168),
.B(n_1041),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1148),
.A2(n_1120),
.B1(n_1109),
.B2(n_1067),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1137),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_1146),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_998),
.A2(n_1017),
.B(n_1004),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1067),
.A2(n_1164),
.B1(n_1166),
.B2(n_1145),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1029),
.B(n_999),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1014),
.A2(n_1021),
.B(n_1012),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1010),
.A2(n_1164),
.B(n_1068),
.C(n_1151),
.Y(n_1186)
);

OAI22x1_ASAP7_75t_L g1187 ( 
.A1(n_1073),
.A2(n_1142),
.B1(n_1147),
.B2(n_1049),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1153),
.A2(n_1024),
.B(n_996),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1152),
.B(n_1095),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1145),
.A2(n_1117),
.B1(n_1051),
.B2(n_1063),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1076),
.A2(n_1038),
.B(n_1024),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1117),
.A2(n_1051),
.B1(n_1068),
.B2(n_1121),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_1079),
.B(n_1098),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1015),
.A2(n_1101),
.A3(n_1072),
.B(n_1127),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1055),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_1000),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1048),
.B(n_1065),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1037),
.B(n_1016),
.Y(n_1198)
);

NAND2x1p5_ASAP7_75t_L g1199 ( 
.A(n_1000),
.B(n_1018),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1000),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1044),
.A2(n_1161),
.B(n_1090),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1092),
.B(n_1173),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1090),
.A2(n_1036),
.B(n_1025),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1018),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1010),
.A2(n_1151),
.B(n_1158),
.C(n_1001),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1076),
.A2(n_1043),
.B(n_1045),
.Y(n_1206)
);

AOI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1027),
.A2(n_1104),
.B(n_1019),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_SL g1208 ( 
.A1(n_1107),
.A2(n_1108),
.B(n_1111),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1005),
.B(n_1023),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1136),
.B(n_1079),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1129),
.A2(n_1141),
.A3(n_1013),
.B(n_1094),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1043),
.A2(n_1084),
.B(n_1052),
.Y(n_1212)
);

AO21x1_ASAP7_75t_L g1213 ( 
.A1(n_1122),
.A2(n_1143),
.B(n_1128),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1154),
.A2(n_1156),
.B(n_1057),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1114),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1086),
.Y(n_1216)
);

AO21x1_ASAP7_75t_L g1217 ( 
.A1(n_1122),
.A2(n_1111),
.B(n_1108),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1018),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1040),
.A2(n_1053),
.B(n_1163),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1137),
.B(n_1035),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1033),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1022),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1056),
.A2(n_1059),
.B(n_1058),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1080),
.A2(n_1159),
.B(n_1162),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1042),
.A2(n_1061),
.B(n_1155),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_1171),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1150),
.A2(n_1039),
.B(n_1034),
.Y(n_1227)
);

NOR2x1_ASAP7_75t_L g1228 ( 
.A(n_1167),
.B(n_997),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1079),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1136),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1144),
.A2(n_1149),
.B(n_1107),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1130),
.B(n_1077),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1054),
.A2(n_1002),
.B(n_1011),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1050),
.B(n_1081),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1157),
.A2(n_1123),
.B(n_1066),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1077),
.B(n_1100),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1171),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1081),
.B(n_1118),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1171),
.Y(n_1239)
);

NAND2x1_ASAP7_75t_L g1240 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1105),
.A2(n_1002),
.B(n_1160),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1118),
.B(n_1098),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1103),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1103),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1088),
.A2(n_1102),
.B(n_1112),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1144),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1096),
.A2(n_1110),
.B(n_1115),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1030),
.B(n_1087),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1100),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_SL g1250 ( 
.A1(n_1149),
.A2(n_1134),
.B(n_1113),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1099),
.A2(n_1083),
.B(n_1091),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1046),
.A2(n_1070),
.B(n_1074),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1009),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1069),
.A2(n_1089),
.B(n_1032),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1097),
.A2(n_1116),
.B1(n_1113),
.B2(n_1139),
.Y(n_1255)
);

AO21x1_ASAP7_75t_L g1256 ( 
.A1(n_1106),
.A2(n_1124),
.B(n_1119),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1064),
.A2(n_1135),
.B(n_1165),
.Y(n_1257)
);

BUFx8_ASAP7_75t_L g1258 ( 
.A(n_1020),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1134),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1028),
.A2(n_1006),
.B(n_1003),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1132),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1138),
.B(n_1060),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1125),
.A2(n_1131),
.B(n_1126),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1133),
.A2(n_1071),
.B(n_1093),
.Y(n_1264)
);

AND2x6_ASAP7_75t_L g1265 ( 
.A(n_1134),
.B(n_1087),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1140),
.A2(n_1085),
.B(n_1047),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1047),
.A2(n_1082),
.A3(n_1078),
.B(n_1062),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1062),
.A2(n_1026),
.B(n_1086),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1100),
.B(n_1075),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1137),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1137),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_750),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_995),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1172),
.A2(n_1148),
.B1(n_1109),
.B2(n_1120),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1172),
.A2(n_1010),
.B(n_904),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1117),
.A2(n_1145),
.B(n_1108),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1095),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1117),
.A2(n_1145),
.B(n_1108),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1168),
.B(n_863),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_750),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1000),
.B(n_1018),
.Y(n_1283)
);

AOI221x1_ASAP7_75t_L g1284 ( 
.A1(n_1170),
.A2(n_1172),
.B1(n_999),
.B2(n_1174),
.C(n_1169),
.Y(n_1284)
);

INVx3_ASAP7_75t_L g1285 ( 
.A(n_1000),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_998),
.A2(n_1146),
.B(n_1017),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_SL g1287 ( 
.A(n_999),
.B(n_1172),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1000),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1166),
.A2(n_1076),
.B(n_1164),
.Y(n_1289)
);

INVx5_ASAP7_75t_L g1290 ( 
.A(n_1144),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_995),
.A2(n_1166),
.B(n_1170),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_750),
.Y(n_1292)
);

OAI33xp33_ASAP7_75t_L g1293 ( 
.A1(n_1047),
.A2(n_815),
.A3(n_745),
.B1(n_852),
.B2(n_1067),
.B3(n_906),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_998),
.A2(n_1146),
.B(n_1017),
.Y(n_1294)
);

AOI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1172),
.A2(n_904),
.B1(n_999),
.B2(n_849),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1000),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1168),
.B(n_863),
.Y(n_1298)
);

OAI22x1_ASAP7_75t_L g1299 ( 
.A1(n_1073),
.A2(n_906),
.B1(n_849),
.B2(n_855),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1172),
.A2(n_904),
.B(n_849),
.C(n_959),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_750),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1023),
.Y(n_1302)
);

INVx4_ASAP7_75t_L g1303 ( 
.A(n_1000),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1015),
.A2(n_1170),
.A3(n_1174),
.B(n_1169),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_998),
.A2(n_1146),
.B(n_1017),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_995),
.A2(n_1174),
.B(n_1169),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1137),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_998),
.A2(n_1146),
.B(n_1017),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1169),
.A2(n_1174),
.B(n_750),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1015),
.A2(n_1170),
.A3(n_1174),
.B(n_1169),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1137),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1315)
);

BUFx12f_ASAP7_75t_L g1316 ( 
.A(n_1086),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_995),
.A2(n_1166),
.B(n_1170),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1033),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1137),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_998),
.A2(n_1146),
.B(n_1017),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_995),
.A2(n_1174),
.B(n_1169),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1000),
.B(n_1018),
.Y(n_1324)
);

OA22x2_ASAP7_75t_L g1325 ( 
.A1(n_1100),
.A2(n_906),
.B1(n_1172),
.B2(n_1067),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1172),
.A2(n_904),
.B(n_849),
.C(n_959),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1172),
.B(n_492),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_995),
.A2(n_1166),
.B(n_1170),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_998),
.A2(n_1146),
.B(n_1017),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1172),
.B(n_1007),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1215),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1302),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_SL g1334 ( 
.A(n_1190),
.B(n_1300),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1193),
.B(n_1229),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1221),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1195),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1280),
.B(n_1298),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1259),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1278),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1176),
.B(n_1271),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1244),
.B(n_1209),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1327),
.B(n_1176),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1318),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1222),
.B(n_1253),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1224),
.A2(n_1203),
.B(n_1185),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1179),
.A2(n_1190),
.B1(n_1325),
.B2(n_1255),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1253),
.B(n_1232),
.Y(n_1348)
);

CKINVDCx11_ASAP7_75t_R g1349 ( 
.A(n_1316),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1271),
.B(n_1282),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1326),
.A2(n_1295),
.B(n_1276),
.C(n_1205),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1282),
.B(n_1297),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1297),
.B(n_1304),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1304),
.B(n_1305),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1265),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1275),
.B(n_1305),
.Y(n_1356)
);

INVx4_ASAP7_75t_SL g1357 ( 
.A(n_1265),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1310),
.B(n_1315),
.Y(n_1359)
);

AND2x4_ASAP7_75t_L g1360 ( 
.A(n_1236),
.B(n_1230),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1273),
.A2(n_1281),
.B(n_1292),
.Y(n_1361)
);

A2O1A1Ixp33_ASAP7_75t_L g1362 ( 
.A1(n_1276),
.A2(n_1186),
.B(n_1179),
.C(n_1266),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1242),
.B(n_1210),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1290),
.B(n_1246),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1200),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1180),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1301),
.A2(n_1312),
.B(n_1188),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1249),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1270),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_SL g1370 ( 
.A1(n_1263),
.A2(n_1183),
.B(n_1192),
.C(n_1287),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1320),
.B(n_1322),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1200),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1242),
.Y(n_1373)
);

NAND2x1_ASAP7_75t_L g1374 ( 
.A(n_1265),
.B(n_1246),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1330),
.B(n_1320),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1231),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1322),
.A2(n_1330),
.B1(n_1189),
.B2(n_1183),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1325),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1308),
.A2(n_1323),
.B(n_1251),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1272),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1189),
.A2(n_1177),
.B1(n_1184),
.B2(n_1192),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1269),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1177),
.B(n_1184),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1219),
.A2(n_1191),
.B(n_1208),
.Y(n_1384)
);

BUFx12f_ASAP7_75t_L g1385 ( 
.A(n_1258),
.Y(n_1385)
);

INVx5_ASAP7_75t_L g1386 ( 
.A(n_1265),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1191),
.A2(n_1175),
.B(n_1328),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1266),
.A2(n_1254),
.B(n_1235),
.C(n_1255),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1263),
.B(n_1235),
.C(n_1262),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1197),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1268),
.B(n_1290),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1202),
.B(n_1299),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1293),
.B(n_1248),
.Y(n_1393)
);

AOI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1291),
.A2(n_1317),
.B(n_1206),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1234),
.B(n_1238),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1269),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1291),
.A2(n_1206),
.B(n_1227),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1259),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1290),
.B(n_1228),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1234),
.B(n_1238),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1262),
.B(n_1309),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1187),
.B(n_1267),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1314),
.B(n_1319),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1267),
.B(n_1237),
.Y(n_1404)
);

INVx3_ASAP7_75t_SL g1405 ( 
.A(n_1216),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1259),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1257),
.A2(n_1260),
.B(n_1252),
.C(n_1201),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1267),
.B(n_1237),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1285),
.B(n_1288),
.Y(n_1409)
);

OR2x6_ASAP7_75t_L g1410 ( 
.A(n_1250),
.B(n_1240),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1257),
.A2(n_1252),
.B(n_1264),
.C(n_1233),
.Y(n_1411)
);

OR2x6_ASAP7_75t_L g1412 ( 
.A(n_1246),
.B(n_1218),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1258),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1217),
.B(n_1213),
.Y(n_1414)
);

AOI222xp33_ASAP7_75t_L g1415 ( 
.A1(n_1277),
.A2(n_1279),
.B1(n_1265),
.B2(n_1220),
.C1(n_1261),
.C2(n_1196),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1200),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1196),
.B(n_1226),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1194),
.B(n_1211),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1241),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1226),
.B(n_1303),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1284),
.A2(n_1289),
.B(n_1247),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1199),
.Y(n_1422)
);

OR2x6_ASAP7_75t_L g1423 ( 
.A(n_1204),
.B(n_1239),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1204),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1283),
.Y(n_1425)
);

O2A1O1Ixp5_ASAP7_75t_SL g1426 ( 
.A1(n_1256),
.A2(n_1274),
.B(n_1181),
.C(n_1245),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1218),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1324),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1239),
.Y(n_1429)
);

BUFx5_ASAP7_75t_L g1430 ( 
.A(n_1212),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1239),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1296),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1296),
.A2(n_1324),
.B1(n_1214),
.B2(n_1225),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1194),
.B(n_1211),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1211),
.B(n_1194),
.Y(n_1435)
);

AO21x1_ASAP7_75t_L g1436 ( 
.A1(n_1207),
.A2(n_1223),
.B(n_1321),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1306),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1182),
.A2(n_1286),
.B(n_1294),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1313),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1307),
.A2(n_1311),
.B(n_1329),
.Y(n_1440)
);

AND2x6_ASAP7_75t_L g1441 ( 
.A(n_1313),
.B(n_1246),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1195),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1302),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1176),
.B(n_1271),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1225),
.A2(n_1294),
.B(n_1286),
.Y(n_1445)
);

BUFx6f_ASAP7_75t_L g1446 ( 
.A(n_1200),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1278),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1302),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1198),
.B(n_694),
.Y(n_1449)
);

BUFx2_ASAP7_75t_L g1450 ( 
.A(n_1302),
.Y(n_1450)
);

NAND2xp33_ASAP7_75t_L g1451 ( 
.A(n_1300),
.B(n_1172),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1278),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1179),
.A2(n_1172),
.B1(n_1122),
.B2(n_1148),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1300),
.A2(n_1172),
.B1(n_1326),
.B2(n_1275),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1327),
.B(n_1176),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1186),
.A2(n_1183),
.B(n_1276),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1259),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1300),
.A2(n_1172),
.B1(n_1326),
.B2(n_1275),
.Y(n_1459)
);

NAND2x1p5_ASAP7_75t_L g1460 ( 
.A(n_1290),
.B(n_1193),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1193),
.B(n_1243),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1259),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1176),
.B(n_1271),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1278),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1224),
.A2(n_1174),
.B(n_1169),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1193),
.B(n_1243),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1278),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1302),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1179),
.A2(n_1148),
.B1(n_1293),
.B2(n_1172),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1215),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1259),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1224),
.A2(n_1174),
.B(n_1169),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1224),
.A2(n_1174),
.B(n_1169),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1179),
.A2(n_1148),
.B1(n_1073),
.B2(n_1122),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1300),
.A2(n_1172),
.B(n_1326),
.C(n_694),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1225),
.A2(n_1294),
.B(n_1286),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1176),
.B(n_1271),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1176),
.B(n_1271),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1259),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_L g1480 ( 
.A(n_1300),
.B(n_1172),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_SL g1481 ( 
.A1(n_1263),
.A2(n_855),
.B(n_849),
.C(n_838),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1316),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1193),
.B(n_1243),
.Y(n_1483)
);

INVx6_ASAP7_75t_L g1484 ( 
.A(n_1355),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1474),
.A2(n_1454),
.B1(n_1334),
.B2(n_1347),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1454),
.A2(n_1334),
.B1(n_1469),
.B2(n_1455),
.Y(n_1486)
);

AND2x4_ASAP7_75t_L g1487 ( 
.A(n_1357),
.B(n_1355),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1470),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1340),
.Y(n_1490)
);

INVx6_ASAP7_75t_L g1491 ( 
.A(n_1355),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1344),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1377),
.B(n_1381),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1447),
.Y(n_1494)
);

INVx3_ASAP7_75t_L g1495 ( 
.A(n_1386),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1336),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1452),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1455),
.A2(n_1459),
.B1(n_1480),
.B2(n_1451),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1378),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1467),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1354),
.B(n_1371),
.Y(n_1501)
);

NAND2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1341),
.B(n_1350),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1421),
.A2(n_1379),
.B(n_1407),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1357),
.B(n_1410),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1341),
.A2(n_1463),
.B1(n_1359),
.B2(n_1353),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1459),
.A2(n_1389),
.B1(n_1449),
.B2(n_1457),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1331),
.Y(n_1508)
);

AO21x2_ASAP7_75t_L g1509 ( 
.A1(n_1438),
.A2(n_1440),
.B(n_1376),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1367),
.A2(n_1361),
.B(n_1465),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1429),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1333),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1350),
.A2(n_1463),
.B1(n_1477),
.B2(n_1359),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1373),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1453),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1366),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1441),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1369),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1393),
.A2(n_1389),
.B1(n_1402),
.B2(n_1338),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1374),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1380),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1445),
.A2(n_1476),
.B(n_1472),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1473),
.A2(n_1426),
.B(n_1346),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1353),
.B(n_1444),
.Y(n_1524)
);

BUFx2_ASAP7_75t_R g1525 ( 
.A(n_1413),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1390),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1384),
.A2(n_1436),
.B(n_1419),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1370),
.A2(n_1397),
.B(n_1433),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1441),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1395),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1408),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1414),
.A2(n_1457),
.B1(n_1377),
.B2(n_1456),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1403),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1395),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1443),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1343),
.A2(n_1342),
.B1(n_1387),
.B2(n_1394),
.Y(n_1536)
);

AOI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1435),
.A2(n_1381),
.B(n_1392),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1335),
.Y(n_1538)
);

OAI21xp33_ASAP7_75t_L g1539 ( 
.A1(n_1388),
.A2(n_1478),
.B(n_1477),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1404),
.B(n_1437),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1441),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1444),
.A2(n_1478),
.B1(n_1382),
.B2(n_1396),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1383),
.B(n_1352),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1342),
.A2(n_1375),
.B1(n_1450),
.B2(n_1448),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1410),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1410),
.B(n_1360),
.Y(n_1546)
);

CKINVDCx6p67_ASAP7_75t_R g1547 ( 
.A(n_1385),
.Y(n_1547)
);

AO21x2_ASAP7_75t_L g1548 ( 
.A1(n_1411),
.A2(n_1481),
.B(n_1362),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1348),
.A2(n_1360),
.B1(n_1368),
.B2(n_1468),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1441),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1383),
.Y(n_1551)
);

CKINVDCx6p67_ASAP7_75t_R g1552 ( 
.A(n_1405),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1439),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1418),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1363),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1363),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1400),
.B(n_1351),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1409),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1422),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1434),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1475),
.B(n_1401),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1335),
.B(n_1348),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1428),
.Y(n_1563)
);

CKINVDCx11_ASAP7_75t_R g1564 ( 
.A(n_1349),
.Y(n_1564)
);

INVx4_ASAP7_75t_SL g1565 ( 
.A(n_1423),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1423),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1337),
.A2(n_1442),
.B1(n_1482),
.B2(n_1345),
.Y(n_1567)
);

INVx4_ASAP7_75t_L g1568 ( 
.A(n_1412),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1415),
.A2(n_1430),
.B(n_1425),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1399),
.B(n_1420),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1430),
.Y(n_1571)
);

CKINVDCx5p33_ASAP7_75t_R g1572 ( 
.A(n_1332),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1460),
.A2(n_1412),
.B1(n_1432),
.B2(n_1416),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1461),
.A2(n_1483),
.B1(n_1466),
.B2(n_1339),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1412),
.A2(n_1364),
.B1(n_1339),
.B2(n_1462),
.Y(n_1575)
);

AO21x1_ASAP7_75t_L g1576 ( 
.A1(n_1415),
.A2(n_1430),
.B(n_1417),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_SL g1577 ( 
.A1(n_1479),
.A2(n_1471),
.B1(n_1462),
.B2(n_1398),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1417),
.A2(n_1420),
.B1(n_1471),
.B2(n_1398),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_SL g1579 ( 
.A1(n_1427),
.A2(n_1430),
.B(n_1479),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1406),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1431),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1406),
.B(n_1458),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1365),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1365),
.A2(n_1372),
.B1(n_1424),
.B2(n_1446),
.Y(n_1584)
);

AO21x1_ASAP7_75t_L g1585 ( 
.A1(n_1372),
.A2(n_1424),
.B(n_1446),
.Y(n_1585)
);

CKINVDCx20_ASAP7_75t_R g1586 ( 
.A(n_1424),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1464),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1378),
.Y(n_1588)
);

CKINVDCx11_ASAP7_75t_R g1589 ( 
.A(n_1385),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1474),
.A2(n_1148),
.B1(n_1454),
.B2(n_1122),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1474),
.A2(n_1148),
.B1(n_1454),
.B2(n_1122),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1474),
.B(n_1454),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1378),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1464),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1470),
.Y(n_1598)
);

CKINVDCx20_ASAP7_75t_R g1599 ( 
.A(n_1337),
.Y(n_1599)
);

BUFx10_ASAP7_75t_L g1600 ( 
.A(n_1345),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1344),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1474),
.A2(n_1172),
.B1(n_1275),
.B2(n_1454),
.Y(n_1602)
);

BUFx3_ASAP7_75t_L g1603 ( 
.A(n_1470),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1464),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1464),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_SL g1606 ( 
.A1(n_1334),
.A2(n_1148),
.B1(n_1122),
.B2(n_1073),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1464),
.Y(n_1607)
);

INVx6_ASAP7_75t_L g1608 ( 
.A(n_1355),
.Y(n_1608)
);

BUFx2_ASAP7_75t_R g1609 ( 
.A(n_1413),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1464),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1464),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1464),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1464),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1464),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1445),
.A2(n_1476),
.B(n_1438),
.Y(n_1615)
);

BUFx12f_ASAP7_75t_L g1616 ( 
.A(n_1349),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1355),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1354),
.B(n_1371),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1355),
.Y(n_1619)
);

CKINVDCx5p33_ASAP7_75t_R g1620 ( 
.A(n_1337),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1378),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1464),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1421),
.A2(n_1379),
.B(n_1407),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1358),
.B(n_1356),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1464),
.Y(n_1625)
);

NAND2x1_ASAP7_75t_L g1626 ( 
.A(n_1410),
.B(n_1231),
.Y(n_1626)
);

CKINVDCx11_ASAP7_75t_R g1627 ( 
.A(n_1385),
.Y(n_1627)
);

BUFx6f_ASAP7_75t_L g1628 ( 
.A(n_1355),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1355),
.B(n_1386),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1464),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1554),
.B(n_1560),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1492),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1500),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1554),
.B(n_1560),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1505),
.B(n_1555),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1601),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1512),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1599),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1537),
.Y(n_1639)
);

NAND2x1_ASAP7_75t_L g1640 ( 
.A(n_1545),
.B(n_1505),
.Y(n_1640)
);

NAND2x1_ASAP7_75t_L g1641 ( 
.A(n_1545),
.B(n_1505),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1617),
.Y(n_1642)
);

BUFx5_ASAP7_75t_L g1643 ( 
.A(n_1526),
.Y(n_1643)
);

HB1xp67_ASAP7_75t_L g1644 ( 
.A(n_1556),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1626),
.B(n_1545),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1556),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1606),
.A2(n_1592),
.B1(n_1590),
.B2(n_1591),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1531),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1488),
.B(n_1594),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1489),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1615),
.A2(n_1522),
.B(n_1527),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1530),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1514),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1493),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1496),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1530),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1493),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1540),
.Y(n_1658)
);

OA21x2_ASAP7_75t_L g1659 ( 
.A1(n_1523),
.A2(n_1528),
.B(n_1576),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1551),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1540),
.Y(n_1661)
);

BUFx12f_ASAP7_75t_L g1662 ( 
.A(n_1564),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1551),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1555),
.B(n_1546),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1571),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1501),
.B(n_1618),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1599),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1539),
.A2(n_1513),
.B(n_1506),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1571),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1555),
.B(n_1546),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1489),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1617),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1546),
.B(n_1487),
.Y(n_1673)
);

INVxp33_ASAP7_75t_L g1674 ( 
.A(n_1562),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1502),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1499),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1517),
.Y(n_1677)
);

BUFx12f_ASAP7_75t_L g1678 ( 
.A(n_1564),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1529),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1529),
.Y(n_1680)
);

INVxp67_ASAP7_75t_SL g1681 ( 
.A(n_1558),
.Y(n_1681)
);

OAI21x1_ASAP7_75t_SL g1682 ( 
.A1(n_1579),
.A2(n_1498),
.B(n_1585),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1541),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1541),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1598),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1550),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1550),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1504),
.A2(n_1623),
.B(n_1579),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1490),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1624),
.B(n_1503),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1624),
.B(n_1503),
.Y(n_1693)
);

HB1xp67_ASAP7_75t_L g1694 ( 
.A(n_1499),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1524),
.B(n_1543),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1519),
.B(n_1548),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1494),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1534),
.B(n_1557),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1588),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1497),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1502),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1588),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1557),
.B(n_1507),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1569),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_1620),
.Y(n_1705)
);

NAND2xp33_ASAP7_75t_R g1706 ( 
.A(n_1620),
.B(n_1572),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1548),
.B(n_1532),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1548),
.B(n_1536),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1504),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1510),
.A2(n_1561),
.B(n_1623),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1593),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1593),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1576),
.Y(n_1713)
);

OA21x2_ASAP7_75t_L g1714 ( 
.A1(n_1486),
.A2(n_1592),
.B(n_1485),
.Y(n_1714)
);

CKINVDCx6p67_ASAP7_75t_R g1715 ( 
.A(n_1616),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1621),
.B(n_1607),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1621),
.B(n_1613),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1553),
.B(n_1602),
.Y(n_1718)
);

INVxp67_ASAP7_75t_L g1719 ( 
.A(n_1533),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1622),
.B(n_1587),
.Y(n_1720)
);

AO21x2_ASAP7_75t_L g1721 ( 
.A1(n_1509),
.A2(n_1510),
.B(n_1604),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1598),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1553),
.B(n_1622),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1510),
.Y(n_1724)
);

CKINVDCx20_ASAP7_75t_R g1725 ( 
.A(n_1589),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1630),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1487),
.B(n_1565),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1595),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1605),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1610),
.B(n_1612),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1611),
.B(n_1625),
.Y(n_1731)
);

BUFx3_ASAP7_75t_L g1732 ( 
.A(n_1650),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1638),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1690),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1690),
.Y(n_1735)
);

BUFx12f_ASAP7_75t_L g1736 ( 
.A(n_1662),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1697),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1713),
.B(n_1509),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1713),
.B(n_1515),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1650),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1676),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1695),
.B(n_1508),
.Y(n_1742)
);

OAI211xp5_ASAP7_75t_L g1743 ( 
.A1(n_1647),
.A2(n_1542),
.B(n_1544),
.C(n_1549),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1694),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1695),
.B(n_1614),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1696),
.B(n_1535),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1727),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1699),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1696),
.B(n_1559),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1698),
.B(n_1521),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1692),
.B(n_1563),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1692),
.B(n_1516),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1693),
.B(n_1631),
.Y(n_1753)
);

NOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1671),
.B(n_1686),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1700),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1658),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1693),
.B(n_1518),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1658),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1706),
.Y(n_1759)
);

INVx3_ASAP7_75t_L g1760 ( 
.A(n_1640),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1702),
.Y(n_1761)
);

INVx3_ASAP7_75t_L g1762 ( 
.A(n_1640),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1708),
.B(n_1566),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1708),
.B(n_1566),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1714),
.A2(n_1574),
.B1(n_1538),
.B2(n_1616),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1631),
.B(n_1580),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1649),
.B(n_1495),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1634),
.Y(n_1768)
);

OR2x2_ASAP7_75t_SL g1769 ( 
.A(n_1714),
.B(n_1718),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1649),
.B(n_1495),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1634),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1674),
.B(n_1572),
.Y(n_1772)
);

NAND2xp33_ASAP7_75t_L g1773 ( 
.A(n_1703),
.B(n_1628),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1648),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1636),
.B(n_1538),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1683),
.B(n_1619),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1643),
.Y(n_1777)
);

AOI31xp33_ASAP7_75t_L g1778 ( 
.A1(n_1718),
.A2(n_1629),
.A3(n_1570),
.B(n_1577),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1707),
.B(n_1582),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1691),
.B(n_1520),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1642),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1653),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1661),
.B(n_1565),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1654),
.B(n_1520),
.Y(n_1784)
);

BUFx3_ASAP7_75t_L g1785 ( 
.A(n_1671),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1654),
.B(n_1520),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1703),
.B(n_1570),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1657),
.B(n_1583),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1641),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1666),
.B(n_1573),
.Y(n_1790)
);

NAND2x1_ASAP7_75t_L g1791 ( 
.A(n_1645),
.B(n_1484),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1707),
.B(n_1583),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1716),
.B(n_1568),
.Y(n_1793)
);

NOR2xp33_ASAP7_75t_L g1794 ( 
.A(n_1638),
.B(n_1603),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1717),
.B(n_1665),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1681),
.B(n_1578),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1714),
.A2(n_1484),
.B1(n_1491),
.B2(n_1608),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1669),
.B(n_1711),
.Y(n_1798)
);

AND2x4_ASAP7_75t_SL g1799 ( 
.A(n_1727),
.B(n_1600),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1668),
.B(n_1603),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1719),
.B1(n_1632),
.B2(n_1637),
.C(n_1655),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1743),
.B(n_1710),
.C(n_1714),
.Y(n_1802)
);

OAI22xp5_ASAP7_75t_L g1803 ( 
.A1(n_1765),
.A2(n_1667),
.B1(n_1722),
.B2(n_1715),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1734),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1782),
.B(n_1712),
.Y(n_1805)
);

OAI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1778),
.A2(n_1645),
.B1(n_1641),
.B2(n_1715),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1741),
.B(n_1644),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1744),
.B(n_1646),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1753),
.B(n_1704),
.Y(n_1809)
);

AOI21xp33_ASAP7_75t_L g1810 ( 
.A1(n_1746),
.A2(n_1797),
.B(n_1779),
.Y(n_1810)
);

NAND3xp33_ASAP7_75t_L g1811 ( 
.A(n_1746),
.B(n_1790),
.C(n_1796),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1748),
.B(n_1726),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1761),
.B(n_1726),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1768),
.B(n_1771),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1768),
.B(n_1729),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1771),
.B(n_1728),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1734),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1798),
.B(n_1728),
.Y(n_1818)
);

OA21x2_ASAP7_75t_L g1819 ( 
.A1(n_1777),
.A2(n_1689),
.B(n_1651),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1773),
.A2(n_1662),
.B1(n_1678),
.B2(n_1673),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1735),
.Y(n_1821)
);

NAND4xp25_ASAP7_75t_L g1822 ( 
.A(n_1739),
.B(n_1723),
.C(n_1731),
.D(n_1730),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1795),
.B(n_1677),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1798),
.B(n_1679),
.Y(n_1824)
);

AOI211xp5_ASAP7_75t_SL g1825 ( 
.A1(n_1773),
.A2(n_1687),
.B(n_1688),
.C(n_1685),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1787),
.A2(n_1552),
.B1(n_1547),
.B2(n_1645),
.C(n_1687),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1793),
.B(n_1680),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1745),
.B(n_1742),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1735),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1793),
.B(n_1684),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1767),
.B(n_1685),
.Y(n_1831)
);

AOI221xp5_ASAP7_75t_L g1832 ( 
.A1(n_1750),
.A2(n_1688),
.B1(n_1720),
.B2(n_1633),
.C(n_1682),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1772),
.A2(n_1733),
.B1(n_1791),
.B2(n_1775),
.C(n_1794),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1763),
.A2(n_1552),
.B1(n_1547),
.B2(n_1645),
.C(n_1584),
.Y(n_1834)
);

OAI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1759),
.A2(n_1791),
.B1(n_1736),
.B2(n_1678),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1745),
.B(n_1643),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1759),
.A2(n_1667),
.B1(n_1491),
.B2(n_1484),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1788),
.B(n_1720),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1754),
.B(n_1664),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1788),
.B(n_1652),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1736),
.B(n_1705),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1770),
.B(n_1652),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1738),
.B(n_1659),
.C(n_1724),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1770),
.B(n_1656),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1737),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1783),
.A2(n_1673),
.B1(n_1727),
.B2(n_1682),
.Y(n_1846)
);

OAI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1769),
.A2(n_1484),
.B1(n_1491),
.B2(n_1608),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1776),
.B(n_1659),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1780),
.B(n_1659),
.Y(n_1849)
);

NOR3xp33_ASAP7_75t_L g1850 ( 
.A(n_1781),
.B(n_1672),
.C(n_1675),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1774),
.B(n_1660),
.Y(n_1851)
);

NAND4xp25_ASAP7_75t_L g1852 ( 
.A(n_1749),
.B(n_1792),
.C(n_1763),
.D(n_1764),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1752),
.A2(n_1757),
.B1(n_1751),
.B2(n_1786),
.C(n_1784),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1756),
.B(n_1721),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1756),
.B(n_1721),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1738),
.B(n_1724),
.C(n_1639),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1732),
.B(n_1705),
.Y(n_1857)
);

AND2x2_ASAP7_75t_SL g1858 ( 
.A(n_1799),
.B(n_1673),
.Y(n_1858)
);

NAND2xp33_ASAP7_75t_SL g1859 ( 
.A(n_1747),
.B(n_1725),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1766),
.B(n_1663),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1764),
.A2(n_1670),
.B1(n_1635),
.B2(n_1701),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1758),
.B(n_1721),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1854),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1804),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1849),
.B(n_1760),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1804),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1817),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1817),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1829),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1852),
.B(n_1769),
.Y(n_1870)
);

BUFx3_ASAP7_75t_L g1871 ( 
.A(n_1854),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1848),
.B(n_1809),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1821),
.Y(n_1873)
);

BUFx2_ASAP7_75t_L g1874 ( 
.A(n_1855),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1843),
.B(n_1792),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1845),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1855),
.B(n_1709),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1833),
.B(n_1732),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1845),
.Y(n_1879)
);

NAND2x1p5_ASAP7_75t_L g1880 ( 
.A(n_1839),
.B(n_1760),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1819),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1862),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1814),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1819),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1819),
.Y(n_1885)
);

INVx5_ASAP7_75t_L g1886 ( 
.A(n_1862),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1815),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1816),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1812),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1813),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1851),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1831),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1824),
.Y(n_1893)
);

BUFx2_ASAP7_75t_L g1894 ( 
.A(n_1858),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1818),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1850),
.B(n_1760),
.Y(n_1896)
);

INVx3_ASAP7_75t_L g1897 ( 
.A(n_1858),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1839),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1840),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1860),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1856),
.B(n_1755),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1811),
.Y(n_1902)
);

OAI22xp5_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1834),
.B1(n_1820),
.B2(n_1802),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1894),
.B(n_1823),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1875),
.B(n_1807),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1894),
.B(n_1823),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1875),
.B(n_1808),
.Y(n_1907)
);

NOR2x1_ASAP7_75t_L g1908 ( 
.A(n_1878),
.B(n_1835),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1875),
.B(n_1822),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1864),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1864),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1894),
.B(n_1827),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1864),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1869),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1897),
.B(n_1827),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1867),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1902),
.B(n_1853),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1869),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1897),
.B(n_1830),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1898),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1867),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1897),
.B(n_1762),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1889),
.B(n_1805),
.Y(n_1923)
);

O2A1O1Ixp33_ASAP7_75t_L g1924 ( 
.A1(n_1870),
.A2(n_1803),
.B(n_1806),
.C(n_1826),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1869),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1889),
.B(n_1828),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1890),
.B(n_1832),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1890),
.B(n_1838),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1900),
.B(n_1830),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1870),
.B(n_1842),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1897),
.B(n_1824),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1900),
.B(n_1836),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1880),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1878),
.B(n_1841),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1897),
.B(n_1898),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1887),
.Y(n_1936)
);

AND2x2_ASAP7_75t_L g1937 ( 
.A(n_1872),
.B(n_1847),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1866),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1870),
.B(n_1859),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1867),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1876),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1872),
.B(n_1810),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1867),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1866),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1876),
.Y(n_1945)
);

OR2x2_ASAP7_75t_L g1946 ( 
.A(n_1877),
.B(n_1892),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1872),
.B(n_1762),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1868),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1873),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1865),
.B(n_1762),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1876),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1898),
.B(n_1859),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1879),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1877),
.B(n_1844),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1895),
.B(n_1899),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1865),
.B(n_1789),
.Y(n_1956)
);

BUFx2_ASAP7_75t_L g1957 ( 
.A(n_1880),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1879),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1879),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1938),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1935),
.B(n_1865),
.Y(n_1961)
);

OAI21xp33_ASAP7_75t_SL g1962 ( 
.A1(n_1939),
.A2(n_1883),
.B(n_1893),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1952),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1944),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1935),
.B(n_1865),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1927),
.B(n_1895),
.Y(n_1966)
);

INVxp67_ASAP7_75t_L g1967 ( 
.A(n_1917),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1910),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1948),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1910),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1909),
.B(n_1899),
.Y(n_1971)
);

NAND2x1p5_ASAP7_75t_L g1972 ( 
.A(n_1957),
.B(n_1896),
.Y(n_1972)
);

NOR2x2_ASAP7_75t_L g1973 ( 
.A(n_1908),
.B(n_1892),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1923),
.B(n_1887),
.Y(n_1974)
);

HB1xp67_ASAP7_75t_L g1975 ( 
.A(n_1911),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1911),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1913),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1942),
.B(n_1883),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1948),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1913),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1916),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1909),
.B(n_1930),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1916),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1935),
.B(n_1947),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1942),
.B(n_1888),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1921),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1934),
.B(n_1857),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1947),
.B(n_1865),
.Y(n_1988)
);

NAND2x1p5_ASAP7_75t_L g1989 ( 
.A(n_1957),
.B(n_1896),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1903),
.B(n_1905),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1905),
.B(n_1888),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1914),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1914),
.Y(n_1993)
);

INVxp67_ASAP7_75t_L g1994 ( 
.A(n_1907),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1950),
.B(n_1865),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1918),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1907),
.B(n_1891),
.Y(n_1997)
);

NOR2x1p5_ASAP7_75t_SL g1998 ( 
.A(n_1921),
.B(n_1881),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1936),
.B(n_1926),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1930),
.B(n_1891),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1922),
.B(n_1896),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1922),
.B(n_1950),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1956),
.B(n_1874),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1928),
.B(n_1932),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1940),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1956),
.B(n_1874),
.Y(n_2006)
);

OAI21xp33_ASAP7_75t_L g2007 ( 
.A1(n_1924),
.A2(n_1846),
.B(n_1880),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1918),
.Y(n_2008)
);

OR2x2_ASAP7_75t_L g2009 ( 
.A(n_1954),
.B(n_1901),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1922),
.B(n_1896),
.Y(n_2010)
);

AOI22xp5_ASAP7_75t_L g2011 ( 
.A1(n_1937),
.A2(n_1837),
.B1(n_1896),
.B2(n_1783),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1937),
.B(n_1874),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1954),
.B(n_1892),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_1955),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1929),
.B(n_1892),
.Y(n_2015)
);

O2A1O1Ixp33_ASAP7_75t_L g2016 ( 
.A1(n_1933),
.A2(n_1880),
.B(n_1801),
.C(n_1901),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1984),
.B(n_1920),
.Y(n_2017)
);

INVx3_ASAP7_75t_L g2018 ( 
.A(n_1972),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1975),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1984),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1975),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1969),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1982),
.B(n_1946),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1967),
.B(n_1912),
.Y(n_2024)
);

HB1xp67_ASAP7_75t_L g2025 ( 
.A(n_2012),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2012),
.B(n_1912),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1973),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1990),
.A2(n_1896),
.B1(n_1670),
.B2(n_1886),
.Y(n_2028)
);

OAI21xp5_ASAP7_75t_SL g2029 ( 
.A1(n_2016),
.A2(n_1825),
.B(n_1861),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1973),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1968),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_1963),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1966),
.B(n_1904),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1970),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2003),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1969),
.Y(n_2036)
);

CKINVDCx16_ASAP7_75t_R g2037 ( 
.A(n_1987),
.Y(n_2037)
);

OAI31xp33_ASAP7_75t_SL g2038 ( 
.A1(n_2007),
.A2(n_1906),
.A3(n_1904),
.B(n_1931),
.Y(n_2038)
);

INVx2_ASAP7_75t_SL g2039 ( 
.A(n_1979),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1976),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2002),
.B(n_1906),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2002),
.B(n_1931),
.Y(n_2042)
);

NOR2x1_ASAP7_75t_L g2043 ( 
.A(n_1979),
.B(n_1925),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2014),
.B(n_1915),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1978),
.B(n_1946),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1977),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1980),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1992),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1987),
.B(n_1589),
.Y(n_2049)
);

INVx1_ASAP7_75t_SL g2050 ( 
.A(n_1971),
.Y(n_2050)
);

AND2x4_ASAP7_75t_L g2051 ( 
.A(n_2002),
.B(n_1925),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1961),
.B(n_1915),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_1972),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1993),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1996),
.Y(n_2055)
);

OR2x2_ASAP7_75t_L g2056 ( 
.A(n_1985),
.B(n_1901),
.Y(n_2056)
);

INVx1_ASAP7_75t_SL g2057 ( 
.A(n_1999),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1981),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2019),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2019),
.Y(n_2060)
);

OAI32xp33_ASAP7_75t_L g2061 ( 
.A1(n_2027),
.A2(n_1962),
.A3(n_1989),
.B1(n_1994),
.B2(n_2009),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2021),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2053),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2037),
.B(n_2004),
.Y(n_2064)
);

BUFx3_ASAP7_75t_L g2065 ( 
.A(n_2022),
.Y(n_2065)
);

O2A1O1Ixp33_ASAP7_75t_L g2066 ( 
.A1(n_2030),
.A2(n_1989),
.B(n_2000),
.C(n_1997),
.Y(n_2066)
);

OAI221xp5_ASAP7_75t_L g2067 ( 
.A1(n_2038),
.A2(n_2029),
.B1(n_2030),
.B2(n_2050),
.C(n_2057),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2021),
.Y(n_2068)
);

OAI32xp33_ASAP7_75t_L g2069 ( 
.A1(n_2037),
.A2(n_2009),
.A3(n_2003),
.B1(n_2006),
.B2(n_1991),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2031),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_2053),
.Y(n_2071)
);

OAI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2030),
.A2(n_2028),
.B1(n_2032),
.B2(n_2024),
.C(n_2020),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2031),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_2049),
.B(n_1627),
.Y(n_2074)
);

OAI31xp33_ASAP7_75t_SL g2075 ( 
.A1(n_2043),
.A2(n_2010),
.A3(n_2001),
.B(n_1961),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_2033),
.B(n_1627),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2053),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2026),
.B(n_1965),
.Y(n_2078)
);

INVx1_ASAP7_75t_SL g2079 ( 
.A(n_2025),
.Y(n_2079)
);

AOI311xp33_ASAP7_75t_L g2080 ( 
.A1(n_2034),
.A2(n_2047),
.A3(n_2046),
.B(n_2055),
.C(n_2054),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2034),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_2020),
.Y(n_2082)
);

AOI211xp5_ASAP7_75t_L g2083 ( 
.A1(n_2018),
.A2(n_2001),
.B(n_2010),
.C(n_1965),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2026),
.B(n_2041),
.Y(n_2084)
);

AOI21xp33_ASAP7_75t_L g2085 ( 
.A1(n_2018),
.A2(n_1974),
.B(n_1964),
.Y(n_2085)
);

OAI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2018),
.A2(n_2011),
.B1(n_1886),
.B2(n_1871),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2041),
.B(n_1960),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2042),
.B(n_2001),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_2017),
.A2(n_2010),
.B1(n_2006),
.B2(n_1995),
.Y(n_2089)
);

AOI21xp33_ASAP7_75t_L g2090 ( 
.A1(n_2018),
.A2(n_2008),
.B(n_1983),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2084),
.B(n_2017),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2065),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2079),
.B(n_2035),
.Y(n_2093)
);

INVxp33_ASAP7_75t_L g2094 ( 
.A(n_2074),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2084),
.B(n_2042),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_2075),
.B(n_2023),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2082),
.B(n_2035),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_2065),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2088),
.B(n_2051),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2081),
.Y(n_2100)
);

INVx1_ASAP7_75t_SL g2101 ( 
.A(n_2064),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2088),
.B(n_2051),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2081),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2059),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_2063),
.B(n_2022),
.Y(n_2105)
);

INVxp33_ASAP7_75t_L g2106 ( 
.A(n_2076),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2063),
.B(n_2071),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2087),
.B(n_2036),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2059),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2071),
.B(n_2039),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2078),
.B(n_2051),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2078),
.B(n_2051),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2077),
.B(n_2039),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2104),
.Y(n_2114)
);

AOI211xp5_ASAP7_75t_SL g2115 ( 
.A1(n_2092),
.A2(n_2067),
.B(n_2072),
.C(n_2086),
.Y(n_2115)
);

OAI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_2096),
.A2(n_2061),
.B(n_2066),
.Y(n_2116)
);

AOI221x1_ASAP7_75t_L g2117 ( 
.A1(n_2092),
.A2(n_2060),
.B1(n_2068),
.B2(n_2062),
.C(n_2077),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_2106),
.A2(n_2061),
.B(n_2069),
.Y(n_2118)
);

NAND3xp33_ASAP7_75t_L g2119 ( 
.A(n_2098),
.B(n_2080),
.C(n_2083),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2098),
.B(n_2062),
.Y(n_2120)
);

AOI211xp5_ASAP7_75t_L g2121 ( 
.A1(n_2094),
.A2(n_2069),
.B(n_2085),
.C(n_2090),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_2091),
.A2(n_2089),
.B1(n_2044),
.B2(n_2036),
.Y(n_2122)
);

OAI211xp5_ASAP7_75t_SL g2123 ( 
.A1(n_2101),
.A2(n_2073),
.B(n_2070),
.C(n_2036),
.Y(n_2123)
);

AOI21xp33_ASAP7_75t_L g2124 ( 
.A1(n_2093),
.A2(n_2023),
.B(n_2056),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2104),
.Y(n_2125)
);

NAND3xp33_ASAP7_75t_SL g2126 ( 
.A(n_2097),
.B(n_2056),
.C(n_2045),
.Y(n_2126)
);

OAI221xp5_ASAP7_75t_L g2127 ( 
.A1(n_2107),
.A2(n_2113),
.B1(n_2110),
.B2(n_2091),
.C(n_2095),
.Y(n_2127)
);

AOI222xp33_ASAP7_75t_L g2128 ( 
.A1(n_2095),
.A2(n_2043),
.B1(n_1998),
.B2(n_2048),
.C1(n_2054),
.C2(n_2040),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2118),
.B(n_2099),
.Y(n_2129)
);

NOR3x1_ASAP7_75t_L g2130 ( 
.A(n_2119),
.B(n_2109),
.C(n_2108),
.Y(n_2130)
);

NOR3xp33_ASAP7_75t_L g2131 ( 
.A(n_2127),
.B(n_2109),
.C(n_2103),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2116),
.A2(n_2099),
.B1(n_2102),
.B2(n_2111),
.Y(n_2132)
);

AND4x1_ASAP7_75t_L g2133 ( 
.A(n_2115),
.B(n_2102),
.C(n_2112),
.D(n_2111),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_2128),
.B(n_2121),
.Y(n_2134)
);

OAI322xp33_ASAP7_75t_L g2135 ( 
.A1(n_2120),
.A2(n_2108),
.A3(n_2103),
.B1(n_2100),
.B2(n_2112),
.C1(n_2047),
.C2(n_2046),
.Y(n_2135)
);

AO22x2_ASAP7_75t_L g2136 ( 
.A1(n_2117),
.A2(n_2100),
.B1(n_2105),
.B2(n_2048),
.Y(n_2136)
);

NAND5xp2_ASAP7_75t_SL g2137 ( 
.A(n_2122),
.B(n_2105),
.C(n_2052),
.D(n_1995),
.E(n_1988),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_2124),
.Y(n_2138)
);

NOR2xp33_ASAP7_75t_L g2139 ( 
.A(n_2126),
.B(n_2105),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_2123),
.B(n_2045),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2114),
.Y(n_2141)
);

NOR3xp33_ASAP7_75t_L g2142 ( 
.A(n_2134),
.B(n_2125),
.C(n_1511),
.Y(n_2142)
);

NOR3xp33_ASAP7_75t_L g2143 ( 
.A(n_2138),
.B(n_1511),
.C(n_1567),
.Y(n_2143)
);

NOR4xp25_ASAP7_75t_L g2144 ( 
.A(n_2129),
.B(n_2058),
.C(n_2055),
.D(n_2040),
.Y(n_2144)
);

AOI221x1_ASAP7_75t_L g2145 ( 
.A1(n_2136),
.A2(n_2131),
.B1(n_2141),
.B2(n_2139),
.C(n_2132),
.Y(n_2145)
);

NAND5xp2_ASAP7_75t_L g2146 ( 
.A(n_2133),
.B(n_2052),
.C(n_1609),
.D(n_1525),
.E(n_1988),
.Y(n_2146)
);

NOR3xp33_ASAP7_75t_L g2147 ( 
.A(n_2135),
.B(n_1511),
.C(n_2058),
.Y(n_2147)
);

NOR3x1_ASAP7_75t_L g2148 ( 
.A(n_2140),
.B(n_2130),
.C(n_2137),
.Y(n_2148)
);

NOR3xp33_ASAP7_75t_L g2149 ( 
.A(n_2136),
.B(n_2058),
.C(n_1983),
.Y(n_2149)
);

NOR3xp33_ASAP7_75t_L g2150 ( 
.A(n_2134),
.B(n_1986),
.C(n_1981),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2149),
.Y(n_2151)
);

NOR2x1_ASAP7_75t_L g2152 ( 
.A(n_2146),
.B(n_1581),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2145),
.Y(n_2153)
);

AOI22xp5_ASAP7_75t_L g2154 ( 
.A1(n_2143),
.A2(n_1586),
.B1(n_2005),
.B2(n_1986),
.Y(n_2154)
);

NAND3xp33_ASAP7_75t_L g2155 ( 
.A(n_2142),
.B(n_2005),
.C(n_1886),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2148),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2150),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2144),
.B(n_1919),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2147),
.Y(n_2159)
);

NAND3xp33_ASAP7_75t_SL g2160 ( 
.A(n_2153),
.B(n_1586),
.C(n_2013),
.Y(n_2160)
);

NAND4xp75_ASAP7_75t_L g2161 ( 
.A(n_2151),
.B(n_1919),
.C(n_1945),
.D(n_1941),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2156),
.B(n_2015),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_2158),
.B(n_1893),
.Y(n_2163)
);

INVxp33_ASAP7_75t_SL g2164 ( 
.A(n_2157),
.Y(n_2164)
);

OAI22x1_ASAP7_75t_L g2165 ( 
.A1(n_2154),
.A2(n_1886),
.B1(n_1945),
.B2(n_1941),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2152),
.A2(n_1886),
.B1(n_1949),
.B2(n_1943),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2162),
.B(n_2154),
.Y(n_2167)
);

XNOR2x1_ASAP7_75t_L g2168 ( 
.A(n_2166),
.B(n_2159),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2160),
.A2(n_2155),
.B(n_1943),
.Y(n_2169)
);

XNOR2xp5_ASAP7_75t_L g2170 ( 
.A(n_2164),
.B(n_2161),
.Y(n_2170)
);

XNOR2x1_ASAP7_75t_L g2171 ( 
.A(n_2170),
.B(n_2163),
.Y(n_2171)
);

AOI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_2167),
.A2(n_2165),
.B1(n_1959),
.B2(n_1958),
.Y(n_2172)
);

INVx4_ASAP7_75t_L g2173 ( 
.A(n_2171),
.Y(n_2173)
);

NAND4xp75_ASAP7_75t_L g2174 ( 
.A(n_2172),
.B(n_2169),
.C(n_2168),
.D(n_1959),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2173),
.Y(n_2175)
);

OAI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2174),
.A2(n_1940),
.B1(n_1949),
.B2(n_1951),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2175),
.Y(n_2177)
);

INVxp67_ASAP7_75t_L g2178 ( 
.A(n_2176),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2177),
.A2(n_1953),
.B(n_1951),
.Y(n_2179)
);

AOI22xp33_ASAP7_75t_SL g2180 ( 
.A1(n_2178),
.A2(n_1886),
.B1(n_1871),
.B2(n_1863),
.Y(n_2180)
);

AOI221xp5_ASAP7_75t_L g2181 ( 
.A1(n_2179),
.A2(n_1958),
.B1(n_1953),
.B2(n_1884),
.C(n_1881),
.Y(n_2181)
);

AOI322xp5_ASAP7_75t_L g2182 ( 
.A1(n_2181),
.A2(n_2180),
.A3(n_1882),
.B1(n_1884),
.B2(n_1871),
.C1(n_1863),
.C2(n_1886),
.Y(n_2182)
);

AOI221xp5_ASAP7_75t_L g2183 ( 
.A1(n_2182),
.A2(n_1884),
.B1(n_1881),
.B2(n_1885),
.C(n_1740),
.Y(n_2183)
);

AOI211xp5_ASAP7_75t_L g2184 ( 
.A1(n_2183),
.A2(n_1575),
.B(n_1628),
.C(n_1785),
.Y(n_2184)
);


endmodule