module fake_jpeg_5615_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx4_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_5),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_9),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_7),
.B(n_9),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_5),
.B(n_7),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_14),
.A2(n_1),
.B1(n_4),
.B2(n_8),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_21),
.A2(n_23),
.B1(n_19),
.B2(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_14),
.A2(n_16),
.B1(n_17),
.B2(n_13),
.Y(n_23)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_1),
.CI(n_8),
.CON(n_24),
.SN(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_20),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_13),
.B1(n_17),
.B2(n_10),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_34),
.B1(n_12),
.B2(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_15),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_27),
.C(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_46),
.B1(n_31),
.B2(n_30),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_22),
.C(n_24),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_10),
.C(n_11),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_33),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_36),
.Y(n_58)
);

XOR2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_31),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_54),
.C(n_43),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_24),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_45),
.C(n_36),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_47),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_57),
.B(n_61),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_59),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_43),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.C(n_62),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_70),
.B2(n_71),
.Y(n_74)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);


endmodule