module real_jpeg_26366_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_352, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_352;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_61),
.B1(n_66),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_1),
.A2(n_30),
.B1(n_33),
.B2(n_61),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_1),
.A2(n_61),
.B1(n_83),
.B2(n_94),
.Y(n_263)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_4),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_4),
.A2(n_30),
.B1(n_33),
.B2(n_77),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_77),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_77),
.B1(n_83),
.B2(n_93),
.Y(n_230)
);

INVx8_ASAP7_75t_SL g90 ( 
.A(n_5),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_80),
.B1(n_92),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_6),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_6),
.A2(n_66),
.B1(n_69),
.B2(n_98),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_98),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_30),
.B1(n_33),
.B2(n_98),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_8),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_8),
.B(n_95),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_8),
.B(n_30),
.C(n_44),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_84),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_75),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_29),
.B1(n_37),
.B2(n_170),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_9),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_9),
.A2(n_34),
.B1(n_66),
.B2(n_69),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_9),
.A2(n_34),
.B1(n_94),
.B2(n_285),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_10),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_40),
.B1(n_66),
.B2(n_69),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g284 ( 
.A1(n_10),
.A2(n_40),
.B1(n_86),
.B2(n_285),
.Y(n_284)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_13),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_13),
.A2(n_68),
.B1(n_83),
.B2(n_93),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_13),
.A2(n_30),
.B1(n_33),
.B2(n_68),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_14),
.A2(n_30),
.B1(n_33),
.B2(n_49),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_14),
.A2(n_49),
.B1(n_66),
.B2(n_69),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_14),
.A2(n_49),
.B1(n_81),
.B2(n_93),
.Y(n_302)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_345),
.C(n_350),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_343),
.B(n_348),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_330),
.B(n_342),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_297),
.A3(n_323),
.B1(n_328),
.B2(n_329),
.C(n_352),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_271),
.B(n_296),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_247),
.B(n_270),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_134),
.B(n_221),
.C(n_246),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_118),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_24),
.B(n_118),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_99),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_26),
.B(n_56),
.C(n_99),
.Y(n_222)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_28),
.B(n_41),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_29),
.A2(n_32),
.B1(n_37),
.B2(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_29),
.B(n_39),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_29),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_29),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_29),
.A2(n_163),
.B1(n_170),
.B2(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_29),
.A2(n_37),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g132 ( 
.A(n_31),
.Y(n_132)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_31),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_33),
.B(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_36),
.A2(n_157),
.B(n_161),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_38),
.B(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_50),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_42),
.A2(n_53),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_42),
.A2(n_53),
.B1(n_146),
.B2(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_42),
.B(n_84),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_42),
.A2(n_46),
.B1(n_53),
.B2(n_242),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_42),
.A2(n_53),
.B(n_59),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_48),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_47),
.B(n_66),
.C(n_73),
.Y(n_189)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_48),
.B(n_142),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_48),
.A2(n_72),
.B(n_188),
.C(n_189),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_50),
.B(n_211),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_52),
.A2(n_63),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_59),
.B(n_62),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_53),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_53),
.A2(n_62),
.B(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.C(n_78),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_57),
.A2(n_58),
.B1(n_64),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_60),
.B(n_63),
.Y(n_211)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_65),
.Y(n_127)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_69),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_85),
.B(n_89),
.C(n_116),
.Y(n_115)
);

HAxp5_ASAP7_75t_SL g188 ( 
.A(n_66),
.B(n_84),
.CON(n_188),
.SN(n_188)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_86),
.C(n_90),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_70),
.A2(n_75),
.B1(n_126),
.B2(n_188),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_70),
.B(n_235),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_70),
.A2(n_75),
.B1(n_291),
.B2(n_292),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_70),
.A2(n_75),
.B(n_110),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_108),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_71),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_75),
.B(n_235),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_78),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_87),
.B1(n_95),
.B2(n_96),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B(n_85),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_84),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_84),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_87),
.A2(n_95),
.B1(n_105),
.B2(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_87),
.B(n_284),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_87),
.A2(n_95),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_87),
.A2(n_321),
.B(n_337),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_87),
.A2(n_95),
.B(n_263),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_88),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_88),
.A2(n_302),
.B(n_303),
.Y(n_301)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_94),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_95),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_95),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_111),
.B2(n_117),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_102),
.B(n_106),
.C(n_117),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_103),
.A2(n_261),
.B(n_262),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_103),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_108),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_108),
.A2(n_234),
.B(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_109),
.B(n_266),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_115),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_119),
.B(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_122),
.B(n_123),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.C(n_130),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_124),
.B(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_133),
.B(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_220),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_215),
.B(n_219),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_200),
.B(n_214),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_184),
.B(n_199),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_158),
.B(n_183),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_152),
.C(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_157),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_167),
.B(n_182),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_165),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_176),
.B(n_181),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_171),
.Y(n_168)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_198),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_198),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_194),
.C(n_197),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_192),
.Y(n_208)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_201),
.B(n_202),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_209),
.C(n_212),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_218),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_223),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_245),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_224)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_229),
.C(n_231),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_243),
.C(n_245),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_269),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_257),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_257),
.C(n_269),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_253),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_252),
.A2(n_277),
.B(n_281),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_255),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_255),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_267),
.B2(n_268),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_264),
.C(n_268),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_262),
.B(n_303),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_272),
.B(n_273),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_295),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_287),
.B2(n_288),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_287),
.C(n_295),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_286),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_283),
.Y(n_337)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_294),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_294),
.A2(n_299),
.B1(n_310),
.B2(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_312),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_312),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_310),
.C(n_311),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_304),
.B2(n_309),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_301),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_301),
.B(n_305),
.C(n_308),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_301),
.B(n_315),
.C(n_322),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_302),
.Y(n_320)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_307),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_308),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_317),
.C(n_319),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_332),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_340),
.B2(n_341),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_335),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_336),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_338),
.C(n_340),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_345),
.Y(n_349)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_347),
.B(n_349),
.Y(n_348)
);


endmodule