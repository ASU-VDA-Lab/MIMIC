module fake_aes_8640_n_710 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_710);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_710;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_599;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_135;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_466;
wire n_302;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_565;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_446;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_17), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_42), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_49), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_62), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_46), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_8), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_22), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_47), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_45), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_15), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_50), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_23), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_55), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_39), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_7), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_67), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_73), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_29), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_31), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_61), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_77), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_64), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_4), .B(n_35), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_16), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_15), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_5), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_56), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
BUFx6f_ASAP7_75t_SL g113 ( .A(n_13), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_44), .Y(n_114) );
INVx4_ASAP7_75t_R g115 ( .A(n_66), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_80), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_24), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_21), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_54), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_71), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_18), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_52), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_65), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_68), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_6), .Y(n_127) );
INVxp33_ASAP7_75t_SL g128 ( .A(n_3), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_74), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_27), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_122), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_122), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_109), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_122), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_109), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_83), .B(n_0), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_97), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_109), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_113), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_112), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_129), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_97), .B(n_100), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_94), .B(n_1), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_130), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_130), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_104), .B(n_1), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_130), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
NOR2xp67_ASAP7_75t_L g153 ( .A(n_118), .B(n_2), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_81), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_84), .Y(n_155) );
BUFx3_ASAP7_75t_L g156 ( .A(n_84), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_86), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_113), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_92), .Y(n_160) );
BUFx2_ASAP7_75t_L g161 ( .A(n_82), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_98), .B(n_2), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_113), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_98), .B(n_3), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_110), .B(n_4), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_108), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_88), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_95), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_113), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_95), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_99), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_87), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_96), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_99), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_161), .Y(n_176) );
INVx4_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_175), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_161), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_142), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_159), .B(n_85), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_142), .Y(n_184) );
INVx6_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
OR2x2_ASAP7_75t_L g188 ( .A(n_168), .B(n_88), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_147), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_144), .B(n_93), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_131), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_161), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_144), .A2(n_128), .B1(n_127), .B2(n_110), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_147), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_175), .Y(n_195) );
OR2x2_ASAP7_75t_L g196 ( .A(n_168), .B(n_93), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_173), .Y(n_197) );
INVx5_ASAP7_75t_L g198 ( .A(n_175), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
INVx6_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_131), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_144), .A2(n_127), .B1(n_119), .B2(n_89), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_131), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_167), .B(n_119), .Y(n_205) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_137), .B(n_126), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_147), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_175), .Y(n_208) );
INVx1_ASAP7_75t_SL g209 ( .A(n_167), .Y(n_209) );
OR2x6_ASAP7_75t_L g210 ( .A(n_137), .B(n_126), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_167), .B(n_125), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_134), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_156), .B(n_125), .Y(n_213) );
AND2x4_ASAP7_75t_L g214 ( .A(n_137), .B(n_89), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_175), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
OAI22xp33_ASAP7_75t_SL g218 ( .A1(n_162), .A2(n_90), .B1(n_91), .B2(n_121), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_152), .B(n_111), .Y(n_219) );
OR2x6_ASAP7_75t_L g220 ( .A(n_136), .B(n_111), .Y(n_220) );
INVx5_ASAP7_75t_L g221 ( .A(n_132), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_147), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_154), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_132), .Y(n_224) );
AND2x6_ASAP7_75t_L g225 ( .A(n_146), .B(n_101), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_170), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_152), .B(n_116), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_146), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_157), .B(n_116), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_154), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_134), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_157), .B(n_90), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_158), .A2(n_101), .B1(n_106), .B2(n_121), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_155), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_158), .B(n_124), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_136), .B(n_103), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_155), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_149), .Y(n_239) );
AND2x6_ASAP7_75t_L g240 ( .A(n_146), .B(n_103), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_149), .Y(n_241) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_150), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_169), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_174), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_242), .B(n_150), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_228), .B(n_150), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_176), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_242), .B(n_160), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_228), .B(n_153), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_237), .B(n_160), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_180), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_180), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_178), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_232), .B(n_163), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_209), .B(n_163), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_221), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_211), .B(n_171), .Y(n_258) );
NOR3xp33_ASAP7_75t_SL g259 ( .A(n_197), .B(n_166), .C(n_165), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g260 ( .A(n_209), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_211), .B(n_171), .Y(n_261) );
BUFx6f_ASAP7_75t_L g262 ( .A(n_221), .Y(n_262) );
OR2x2_ASAP7_75t_SL g263 ( .A(n_179), .B(n_166), .Y(n_263) );
NOR3xp33_ASAP7_75t_SL g264 ( .A(n_203), .B(n_165), .C(n_162), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_195), .Y(n_265) );
XOR2xp5_ASAP7_75t_L g266 ( .A(n_244), .B(n_5), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_224), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_208), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_179), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_220), .B(n_153), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_224), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_221), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_221), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_220), .B(n_172), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_220), .B(n_172), .Y(n_275) );
INVx1_ASAP7_75t_SL g276 ( .A(n_192), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g277 ( .A1(n_190), .A2(n_172), .B1(n_169), .B2(n_102), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_188), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_215), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_185), .Y(n_280) );
CKINVDCx6p67_ASAP7_75t_R g281 ( .A(n_210), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_216), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_214), .B(n_169), .Y(n_283) );
BUFx6f_ASAP7_75t_L g284 ( .A(n_186), .Y(n_284) );
INVx3_ASAP7_75t_SL g285 ( .A(n_210), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_186), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_223), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_225), .B(n_132), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_190), .A2(n_105), .B1(n_120), .B2(n_107), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_225), .B(n_132), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_230), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_214), .B(n_143), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_206), .B(n_143), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_225), .B(n_143), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_233), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_232), .A2(n_106), .B1(n_117), .B2(n_143), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_235), .Y(n_297) );
NOR3xp33_ASAP7_75t_SL g298 ( .A(n_203), .B(n_114), .C(n_123), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_238), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_243), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_225), .B(n_143), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_186), .Y(n_302) );
INVx5_ASAP7_75t_L g303 ( .A(n_185), .Y(n_303) );
CKINVDCx16_ASAP7_75t_R g304 ( .A(n_210), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_187), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_191), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_240), .B(n_206), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_240), .B(n_140), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_240), .B(n_140), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_202), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_196), .B(n_133), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_205), .Y(n_312) );
BUFx4f_ASAP7_75t_L g313 ( .A(n_240), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_213), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_213), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_185), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_201), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_218), .A2(n_151), .B1(n_149), .B2(n_145), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_255), .A2(n_236), .B(n_227), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_253), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_SL g321 ( .A1(n_255), .A2(n_229), .B(n_227), .C(n_117), .Y(n_321) );
AOI21x1_ASAP7_75t_L g322 ( .A1(n_274), .A2(n_229), .B(n_184), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_256), .B(n_193), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_293), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_253), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_247), .B(n_226), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_256), .B(n_218), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_247), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_260), .A2(n_226), .B1(n_200), .B2(n_177), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_254), .Y(n_330) );
BUFx10_ASAP7_75t_L g331 ( .A(n_246), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_269), .B(n_219), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_257), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_265), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_276), .B(n_234), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_314), .A2(n_219), .B(n_183), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_293), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_292), .Y(n_339) );
BUFx4_ASAP7_75t_SL g340 ( .A(n_260), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_304), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_257), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_313), .B(n_177), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_292), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_278), .B(n_234), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_280), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_283), .Y(n_347) );
NOR2xp33_ASAP7_75t_R g348 ( .A(n_281), .B(n_200), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g349 ( .A(n_269), .B(n_182), .C(n_133), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_283), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_246), .A2(n_201), .B1(n_181), .B2(n_231), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_250), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_245), .B(n_212), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_265), .Y(n_354) );
INVx5_ASAP7_75t_L g355 ( .A(n_257), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_311), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_313), .B(n_198), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_246), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_258), .A2(n_198), .B(n_204), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_257), .Y(n_360) );
BUFx2_ASAP7_75t_SL g361 ( .A(n_312), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_280), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_311), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_281), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_262), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_268), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_248), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_315), .B(n_198), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_248), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_285), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_261), .B(n_201), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_275), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_261), .B(n_198), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_356), .Y(n_377) );
INVx6_ASAP7_75t_L g378 ( .A(n_355), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_352), .A2(n_318), .B1(n_249), .B2(n_291), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_320), .Y(n_380) );
BUFx3_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
AO31x2_ASAP7_75t_L g382 ( .A1(n_320), .A2(n_145), .A3(n_138), .B(n_141), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_330), .A2(n_285), .B1(n_245), .B2(n_307), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_340), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_326), .Y(n_385) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_323), .A2(n_270), .B(n_249), .C(n_289), .Y(n_386) );
OR2x6_ASAP7_75t_L g387 ( .A(n_361), .B(n_249), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_325), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_332), .B(n_264), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_319), .A2(n_268), .B(n_279), .Y(n_390) );
OR2x6_ASAP7_75t_L g391 ( .A(n_372), .B(n_288), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_326), .A2(n_259), .B1(n_298), .B2(n_277), .Y(n_393) );
AOI21xp5_ASAP7_75t_SL g394 ( .A1(n_325), .A2(n_294), .B(n_301), .Y(n_394) );
OAI22xp5_ASAP7_75t_SL g395 ( .A1(n_341), .A2(n_266), .B1(n_263), .B2(n_290), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_345), .A2(n_263), .B1(n_296), .B2(n_282), .Y(n_396) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_345), .A2(n_299), .B1(n_295), .B2(n_287), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_326), .A2(n_309), .B1(n_308), .B2(n_267), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_332), .B(n_282), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_369), .A2(n_297), .B1(n_300), .B2(n_279), .Y(n_400) );
OAI21xp5_ASAP7_75t_L g401 ( .A1(n_336), .A2(n_359), .B(n_375), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_371), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_353), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_321), .A2(n_145), .B(n_148), .Y(n_404) );
BUFx4f_ASAP7_75t_L g405 ( .A(n_343), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_353), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_324), .Y(n_407) );
CKINVDCx6p67_ASAP7_75t_R g408 ( .A(n_341), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_322), .A2(n_297), .B(n_300), .Y(n_409) );
AOI221xp5_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_344), .B1(n_339), .B2(n_327), .C(n_335), .Y(n_410) );
NAND3xp33_ASAP7_75t_L g411 ( .A(n_401), .B(n_321), .C(n_328), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_403), .B(n_374), .Y(n_412) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_397), .A2(n_335), .B1(n_373), .B2(n_368), .Y(n_414) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_381), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_395), .A2(n_349), .B1(n_358), .B2(n_337), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_393), .B(n_365), .Y(n_417) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_390), .A2(n_354), .B(n_368), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_397), .A2(n_358), .B1(n_347), .B2(n_350), .Y(n_419) );
OR2x2_ASAP7_75t_SL g420 ( .A(n_376), .B(n_348), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_399), .B(n_334), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_380), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_385), .B(n_334), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_380), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_409), .A2(n_370), .B(n_354), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_386), .A2(n_329), .B(n_348), .C(n_351), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_379), .A2(n_135), .B1(n_138), .B2(n_141), .Y(n_427) );
AOI211xp5_ASAP7_75t_L g428 ( .A1(n_396), .A2(n_365), .B(n_370), .C(n_135), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_406), .B(n_333), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_388), .B(n_331), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_409), .A2(n_148), .B(n_217), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_388), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_379), .A2(n_271), .B(n_251), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_377), .A2(n_392), .B1(n_402), .B2(n_387), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_400), .B(n_331), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_387), .A2(n_331), .B1(n_267), .B2(n_363), .Y(n_436) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_383), .A2(n_343), .B1(n_252), .B2(n_267), .C(n_362), .Y(n_437) );
OAI22xp33_ASAP7_75t_L g438 ( .A1(n_387), .A2(n_338), .B1(n_360), .B2(n_355), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_400), .B(n_306), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_421), .B(n_382), .Y(n_441) );
OAI33xp33_ASAP7_75t_L g442 ( .A1(n_414), .A2(n_407), .A3(n_384), .B1(n_357), .B2(n_11), .B3(n_12), .Y(n_442) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_428), .B(n_151), .C(n_149), .Y(n_443) );
INVx4_ASAP7_75t_L g444 ( .A(n_415), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_422), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_414), .B(n_382), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_417), .B(n_384), .C(n_398), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_432), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_424), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_410), .A2(n_391), .B1(n_405), .B2(n_408), .Y(n_450) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_416), .A2(n_394), .B(n_381), .C(n_273), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_412), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_426), .A2(n_391), .B(n_404), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_419), .B(n_391), .Y(n_454) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_428), .A2(n_405), .B1(n_149), .B2(n_151), .C(n_404), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_420), .A2(n_378), .B1(n_360), .B2(n_355), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_413), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_421), .B(n_382), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_420), .A2(n_378), .B1(n_360), .B2(n_355), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_432), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_424), .B(n_382), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_435), .B(n_360), .Y(n_463) );
NOR2x2_ASAP7_75t_L g464 ( .A(n_438), .B(n_378), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_360), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_435), .A2(n_338), .B1(n_366), .B2(n_363), .Y(n_466) );
INVxp67_ASAP7_75t_SL g467 ( .A(n_423), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_437), .A2(n_366), .B1(n_362), .B2(n_346), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_430), .B(n_367), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_415), .B(n_367), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
NOR4xp25_ASAP7_75t_SL g473 ( .A(n_437), .B(n_357), .C(n_115), .D(n_10), .Y(n_473) );
INVx3_ASAP7_75t_L g474 ( .A(n_415), .Y(n_474) );
INVxp67_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g476 ( .A(n_415), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_476), .B(n_415), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_468), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_447), .A2(n_411), .B1(n_434), .B2(n_427), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_468), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_440), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_442), .A2(n_427), .B1(n_411), .B2(n_429), .C(n_436), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_441), .B(n_415), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_441), .B(n_439), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_459), .B(n_433), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_444), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_458), .A2(n_429), .B1(n_439), .B2(n_149), .C(n_151), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_472), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_472), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
OAI221xp5_ASAP7_75t_L g493 ( .A1(n_450), .A2(n_433), .B1(n_418), .B2(n_425), .C(n_346), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_448), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_448), .Y(n_495) );
BUFx2_ASAP7_75t_L g496 ( .A(n_444), .Y(n_496) );
AOI33xp33_ASAP7_75t_L g497 ( .A1(n_452), .A2(n_6), .A3(n_9), .B1(n_10), .B2(n_11), .B3(n_13), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_461), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_465), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_449), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_459), .B(n_433), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_462), .B(n_431), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_462), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_475), .B(n_465), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_446), .B(n_431), .Y(n_508) );
AOI33xp33_ASAP7_75t_L g509 ( .A1(n_473), .A2(n_9), .A3(n_14), .B1(n_16), .B2(n_17), .B3(n_310), .Y(n_509) );
NAND3xp33_ASAP7_75t_L g510 ( .A(n_453), .B(n_149), .C(n_151), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_457), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_457), .B(n_418), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_454), .B(n_151), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_474), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_470), .B(n_151), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_470), .B(n_14), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_474), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_443), .A2(n_306), .B(n_310), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_446), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_444), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_474), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_471), .Y(n_522) );
NAND2x1_ASAP7_75t_SL g523 ( .A(n_463), .B(n_333), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_456), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_471), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
AOI31xp33_ASAP7_75t_L g527 ( .A1(n_460), .A2(n_115), .A3(n_20), .B(n_25), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_463), .Y(n_528) );
AND2x4_ASAP7_75t_L g529 ( .A(n_463), .B(n_367), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_504), .B(n_455), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_479), .A2(n_469), .B1(n_466), .B2(n_464), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_499), .B(n_464), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_481), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_507), .B(n_451), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_502), .B(n_333), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_484), .B(n_19), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_490), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_484), .B(n_26), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_488), .Y(n_540) );
NOR2xp33_ASAP7_75t_R g541 ( .A(n_488), .B(n_342), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_491), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_496), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_484), .B(n_28), .Y(n_544) );
OAI31xp33_ASAP7_75t_L g545 ( .A1(n_516), .A2(n_273), .A3(n_272), .B(n_36), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_487), .B(n_33), .Y(n_546) );
NAND2xp33_ASAP7_75t_SL g547 ( .A(n_496), .B(n_338), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_506), .B(n_342), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_483), .B(n_342), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_516), .B(n_342), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_481), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_483), .B(n_34), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_520), .Y(n_553) );
AO21x1_ASAP7_75t_L g554 ( .A1(n_527), .A2(n_317), .B(n_40), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_491), .Y(n_555) );
CKINVDCx16_ASAP7_75t_R g556 ( .A(n_483), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_510), .A2(n_317), .B(n_303), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_505), .B(n_38), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_505), .B(n_41), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_486), .B(n_189), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_487), .B(n_43), .Y(n_562) );
INVxp33_ASAP7_75t_SL g563 ( .A(n_477), .Y(n_563) );
CKINVDCx8_ASAP7_75t_R g564 ( .A(n_529), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_486), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_528), .B(n_48), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_520), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_515), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_492), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_511), .B(n_51), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_513), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_494), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_494), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_489), .A2(n_317), .B(n_303), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_511), .B(n_53), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_495), .B(n_57), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_478), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_503), .B(n_58), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_524), .A2(n_273), .B1(n_272), .B2(n_262), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_519), .A2(n_199), .B1(n_189), .B2(n_187), .C(n_194), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_503), .B(n_59), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_523), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_478), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_528), .B(n_60), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_480), .B(n_63), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_540), .B(n_523), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_543), .B(n_508), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_533), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_551), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_556), .B(n_525), .Y(n_591) );
AND2x4_ASAP7_75t_L g592 ( .A(n_553), .B(n_525), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_559), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_531), .A2(n_482), .B1(n_525), .B2(n_526), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_565), .Y(n_595) );
INVx1_ASAP7_75t_SL g596 ( .A(n_567), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_563), .B(n_529), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_532), .B(n_522), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_537), .Y(n_599) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_568), .A2(n_521), .B1(n_493), .B2(n_529), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_534), .A2(n_497), .B(n_509), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_554), .A2(n_508), .B1(n_512), .B2(n_514), .Y(n_602) );
OAI22xp33_ASAP7_75t_L g603 ( .A1(n_564), .A2(n_500), .B1(n_501), .B2(n_517), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_572), .Y(n_605) );
OAI21xp33_ASAP7_75t_SL g606 ( .A1(n_536), .A2(n_501), .B(n_500), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_573), .B(n_512), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_541), .Y(n_608) );
AOI211xp5_ASAP7_75t_L g609 ( .A1(n_547), .A2(n_517), .B(n_518), .C(n_222), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_577), .B(n_207), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_547), .A2(n_581), .B(n_545), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_578), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_577), .B(n_207), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_584), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_571), .B(n_207), .Y(n_615) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_541), .Y(n_616) );
OAI31xp33_ASAP7_75t_L g617 ( .A1(n_536), .A2(n_272), .A3(n_72), .B(n_75), .Y(n_617) );
OAI322xp33_ASAP7_75t_L g618 ( .A1(n_571), .A2(n_222), .A3(n_199), .B1(n_241), .B2(n_239), .C1(n_187), .C2(n_189), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_537), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_546), .B(n_69), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_538), .Y(n_621) );
NOR3xp33_ASAP7_75t_SL g622 ( .A(n_530), .B(n_76), .C(n_78), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_568), .B(n_79), .Y(n_623) );
OA21x2_ASAP7_75t_L g624 ( .A1(n_538), .A2(n_194), .B(n_199), .Y(n_624) );
XNOR2x2_ASAP7_75t_L g625 ( .A(n_539), .B(n_303), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_539), .A2(n_194), .B1(n_222), .B2(n_239), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_542), .Y(n_627) );
AOI21xp33_ASAP7_75t_SL g628 ( .A1(n_544), .A2(n_303), .B(n_262), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_546), .B(n_241), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_542), .B(n_241), .Y(n_630) );
NOR2xp33_ASAP7_75t_SL g631 ( .A(n_564), .B(n_303), .Y(n_631) );
NOR2xp67_ASAP7_75t_SL g632 ( .A(n_558), .B(n_262), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_555), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_588), .B(n_555), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_596), .Y(n_635) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_601), .A2(n_583), .B(n_579), .Y(n_636) );
NAND2x1_ASAP7_75t_L g637 ( .A(n_632), .B(n_582), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_606), .A2(n_562), .B(n_560), .C(n_552), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_607), .B(n_562), .Y(n_639) );
XNOR2x2_ASAP7_75t_L g640 ( .A(n_625), .B(n_576), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_599), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_598), .B(n_549), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_589), .B(n_586), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_590), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_619), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_602), .A2(n_580), .B1(n_535), .B2(n_550), .C(n_575), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_593), .B(n_586), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_608), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_621), .Y(n_649) );
NOR3xp33_ASAP7_75t_SL g650 ( .A(n_611), .B(n_561), .C(n_574), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_595), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_604), .B(n_548), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_627), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_605), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_633), .B(n_570), .Y(n_655) );
NOR3xp33_ASAP7_75t_L g656 ( .A(n_618), .B(n_566), .C(n_585), .Y(n_656) );
AOI21xp5_ASAP7_75t_SL g657 ( .A1(n_616), .A2(n_557), .B(n_286), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_612), .Y(n_658) );
BUFx2_ASAP7_75t_L g659 ( .A(n_592), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_614), .Y(n_660) );
XNOR2x1_ASAP7_75t_L g661 ( .A(n_591), .B(n_284), .Y(n_661) );
XNOR2xp5_ASAP7_75t_L g662 ( .A(n_594), .B(n_284), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g663 ( .A(n_592), .B(n_284), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_609), .B(n_286), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_644), .Y(n_665) );
XNOR2xp5_ASAP7_75t_L g666 ( .A(n_635), .B(n_620), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_641), .Y(n_667) );
XNOR2x1_ASAP7_75t_L g668 ( .A(n_640), .B(n_600), .Y(n_668) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_648), .B(n_617), .C(n_622), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_651), .Y(n_670) );
NOR2x1_ASAP7_75t_L g671 ( .A(n_657), .B(n_603), .Y(n_671) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_664), .B(n_624), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_659), .Y(n_673) );
XOR2x2_ASAP7_75t_L g674 ( .A(n_638), .B(n_597), .Y(n_674) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_637), .A2(n_628), .B(n_623), .C(n_587), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_654), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_648), .B(n_615), .Y(n_677) );
NAND4xp25_ASAP7_75t_SL g678 ( .A(n_636), .B(n_626), .C(n_631), .D(n_629), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_642), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_639), .A2(n_610), .B1(n_613), .B2(n_630), .Y(n_680) );
XNOR2x1_ASAP7_75t_L g681 ( .A(n_661), .B(n_302), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_668), .A2(n_650), .B1(n_634), .B2(n_646), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g683 ( .A(n_671), .B(n_650), .C(n_662), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_678), .A2(n_656), .B(n_663), .C(n_647), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_666), .B(n_658), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_674), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g687 ( .A(n_671), .B(n_656), .C(n_660), .Y(n_687) );
OAI32xp33_ASAP7_75t_L g688 ( .A1(n_669), .A2(n_643), .A3(n_655), .B1(n_652), .B2(n_649), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_673), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_677), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_665), .Y(n_691) );
INVx1_ASAP7_75t_SL g692 ( .A(n_681), .Y(n_692) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_675), .B(n_645), .Y(n_693) );
AND3x4_ASAP7_75t_L g694 ( .A(n_672), .B(n_653), .C(n_641), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_670), .A2(n_305), .B1(n_676), .B2(n_679), .C(n_667), .Y(n_695) );
NAND4xp75_ASAP7_75t_L g696 ( .A(n_680), .B(n_671), .C(n_672), .D(n_650), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_668), .A2(n_674), .B1(n_669), .B2(n_673), .Y(n_697) );
OA22x2_ASAP7_75t_L g698 ( .A1(n_697), .A2(n_692), .B1(n_694), .B2(n_682), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_689), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_686), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_690), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_691), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_698), .B(n_683), .C(n_687), .D(n_692), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_698), .A2(n_696), .B1(n_684), .B2(n_693), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_700), .Y(n_705) );
BUFx2_ASAP7_75t_L g706 ( .A(n_705), .Y(n_706) );
NAND2x1_ASAP7_75t_L g707 ( .A(n_704), .B(n_701), .Y(n_707) );
AND2x2_ASAP7_75t_L g708 ( .A(n_706), .B(n_699), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_703), .B1(n_707), .B2(n_700), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_709), .A2(n_688), .B1(n_702), .B2(n_695), .C(n_685), .Y(n_710) );
endmodule