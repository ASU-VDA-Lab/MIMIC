module real_jpeg_25540_n_29 (n_17, n_8, n_0, n_21, n_168, n_2, n_10, n_9, n_12, n_24, n_165, n_166, n_6, n_159, n_28, n_161, n_162, n_167, n_23, n_11, n_14, n_160, n_25, n_163, n_7, n_22, n_18, n_3, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_164, n_158, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_168;
input n_2;
input n_10;
input n_9;
input n_12;
input n_24;
input n_165;
input n_166;
input n_6;
input n_159;
input n_28;
input n_161;
input n_162;
input n_167;
input n_23;
input n_11;
input n_14;
input n_160;
input n_25;
input n_163;
input n_7;
input n_22;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_164;
input n_158;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_0),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_1),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_2),
.A2(n_32),
.B(n_36),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_2),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_2),
.B(n_39),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_3),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_5),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_5),
.B(n_113),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_7),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_7),
.B(n_61),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_8),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_9),
.B(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_10),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_11),
.A2(n_30),
.B(n_156),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_11),
.B(n_33),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_12),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_13),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_13),
.B(n_124),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_14),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_15),
.B(n_96),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_17),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_17),
.B(n_68),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_18),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_18),
.B(n_145),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_19),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_20),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_21),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_22),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_22),
.B(n_130),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_23),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_24),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_66),
.C(n_141),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_27),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_28),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_37),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_34),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_34),
.B(n_151),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_35),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_35),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_35),
.B(n_103),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_35),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B(n_155),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_57),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_45),
.B(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_52),
.B(n_146),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_54),
.Y(n_143)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_55),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_55),
.B(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_154),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_148),
.B(n_153),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_144),
.B(n_147),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B(n_140),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_134),
.B(n_139),
.Y(n_70)
);

OAI321xp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_123),
.A3(n_129),
.B1(n_132),
.B2(n_133),
.C(n_158),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_117),
.B(n_122),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_112),
.B(n_116),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_106),
.B(n_111),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B(n_105),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_99),
.B(n_104),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_95),
.B(n_98),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_89),
.B(n_94),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_88),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_101),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_107),
.B(n_108),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_118),
.B(n_119),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_138),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_159),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_160),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_161),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_162),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_163),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_164),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_165),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_166),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_167),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_168),
.Y(n_131)
);


endmodule