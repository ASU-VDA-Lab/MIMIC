module fake_netlist_6_4400_n_2289 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2289);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2289;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_2209;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_182),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_127),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_60),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_78),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_65),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_16),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_130),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_15),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_89),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_164),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_168),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_46),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_80),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_105),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_9),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_81),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_167),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_68),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_101),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_91),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_173),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_205),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_24),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_149),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_95),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_98),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_40),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_41),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_189),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_185),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_141),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_57),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_55),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_145),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_51),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_52),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_23),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_128),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_177),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_4),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_131),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_48),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_121),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_162),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_12),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_136),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_181),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_204),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_61),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_183),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_8),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_132),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_15),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_27),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_22),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_99),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_92),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_106),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_193),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_77),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_51),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_78),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_71),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_115),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_174),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_186),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_176),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_112),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_27),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_184),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_152),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_67),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_100),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_23),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_188),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_125),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_14),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_50),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_75),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_200),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_13),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_26),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_199),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_203),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_139),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g320 ( 
.A(n_118),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_120),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_82),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_116),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_40),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_114),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_30),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_150),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_221),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_18),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_80),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_143),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_58),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_169),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_72),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_117),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_122),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_70),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_137),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_146),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_6),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_12),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_60),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_66),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_17),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_47),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_24),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_218),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_54),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_34),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_133),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_25),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_179),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_30),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_194),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_55),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_77),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_109),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_11),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_153),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_20),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_82),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_161),
.Y(n_362)
);

BUFx3_ASAP7_75t_L g363 ( 
.A(n_208),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_4),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_28),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_42),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_43),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_160),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_210),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_159),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_111),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_158),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_163),
.Y(n_373)
);

BUFx2_ASAP7_75t_SL g374 ( 
.A(n_212),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_74),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_144),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_88),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_41),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_64),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_13),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_214),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_10),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_73),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_32),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_129),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_198),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_84),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_45),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_20),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_62),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_157),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_85),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_62),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_196),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_47),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_75),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_180),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_66),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_96),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_58),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_11),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_172),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_14),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_138),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_220),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_154),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_64),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_76),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_31),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_53),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_170),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_135),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_70),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_140),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_71),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_192),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_190),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_9),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_38),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_74),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_107),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_191),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_213),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_123),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_175),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_72),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_56),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_102),
.Y(n_428)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_217),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_54),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_219),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_5),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_63),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_87),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_49),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_34),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_59),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_209),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_230),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_268),
.B(n_0),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_306),
.B(n_0),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_223),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_264),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_259),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_230),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_234),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_267),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_409),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_268),
.B(n_1),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_264),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_271),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_319),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_415),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_227),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_234),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_235),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_235),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_228),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_281),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_240),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_R g462 ( 
.A(n_331),
.B(n_86),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_240),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_248),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_306),
.B(n_1),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_231),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_338),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_350),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_238),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_239),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_233),
.B(n_250),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_415),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_411),
.Y(n_474)
);

NOR2xp67_ASAP7_75t_L g475 ( 
.A(n_268),
.B(n_2),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_241),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_373),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_248),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_368),
.B(n_2),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_376),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_242),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_367),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_244),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_406),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_255),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_368),
.B(n_3),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_255),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_263),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_414),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_263),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_251),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_256),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_367),
.Y(n_493)
);

INVx4_ASAP7_75t_R g494 ( 
.A(n_319),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_274),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_274),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_261),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_275),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_275),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_262),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_428),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_R g502 ( 
.A(n_429),
.B(n_90),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_277),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_277),
.Y(n_504)
);

INVxp33_ASAP7_75t_SL g505 ( 
.A(n_435),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_284),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_377),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_278),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_377),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_278),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_287),
.Y(n_511)
);

INVxp33_ASAP7_75t_SL g512 ( 
.A(n_435),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_285),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_287),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_293),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_294),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_320),
.B(n_3),
.Y(n_518)
);

BUFx2_ASAP7_75t_SL g519 ( 
.A(n_270),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_288),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_304),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_224),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_268),
.B(n_6),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_288),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_412),
.Y(n_525)
);

INVxp33_ASAP7_75t_L g526 ( 
.A(n_233),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_340),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_R g528 ( 
.A(n_225),
.B(n_93),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_307),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_310),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_R g531 ( 
.A(n_229),
.B(n_94),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_257),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_311),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_232),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_291),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_312),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_291),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_319),
.B(n_7),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_324),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_298),
.Y(n_540)
);

NOR2xp67_ASAP7_75t_L g541 ( 
.A(n_270),
.B(n_7),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_237),
.Y(n_542)
);

CKINVDCx14_ASAP7_75t_R g543 ( 
.A(n_340),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_243),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_247),
.Y(n_546)
);

INVxp33_ASAP7_75t_SL g547 ( 
.A(n_326),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_329),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_340),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_330),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_332),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_415),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_226),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_334),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_249),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_342),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_335),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_525),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_454),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_525),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_468),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_517),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_453),
.B(n_341),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_473),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_447),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_453),
.B(n_438),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_442),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_544),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_544),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_519),
.B(n_341),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_552),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_552),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_439),
.B(n_253),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_547),
.B(n_309),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_553),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_553),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_446),
.B(n_254),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_472),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_457),
.Y(n_590)
);

OA21x2_ASAP7_75t_L g591 ( 
.A1(n_458),
.A2(n_364),
.B(n_226),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_461),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_463),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_449),
.Y(n_595)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_305),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_478),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_526),
.B(n_341),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_485),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_487),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_488),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_490),
.Y(n_602)
);

BUFx8_ASAP7_75t_L g603 ( 
.A(n_443),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_521),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_505),
.A2(n_292),
.B1(n_295),
.B2(n_273),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_495),
.B(n_258),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_522),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_498),
.B(n_260),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_499),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_503),
.B(n_269),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_450),
.B(n_335),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_507),
.B(n_532),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_504),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_508),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_510),
.B(n_272),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_509),
.B(n_303),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_511),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_514),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_475),
.B(n_335),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_520),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_524),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_317),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_535),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_537),
.B(n_540),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_538),
.B(n_279),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_443),
.B(n_305),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_465),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_441),
.B(n_283),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_518),
.B(n_363),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_486),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_529),
.B(n_363),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_512),
.A2(n_390),
.B1(n_379),
.B2(n_361),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_455),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_462),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_528),
.B(n_289),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_451),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_449),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_455),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_482),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_459),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_531),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_459),
.Y(n_648)
);

NAND3xp33_ASAP7_75t_L g649 ( 
.A(n_633),
.B(n_246),
.C(n_298),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_563),
.Y(n_650)
);

INVx5_ASAP7_75t_L g651 ( 
.A(n_558),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_591),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_558),
.Y(n_653)
);

AND2x6_ASAP7_75t_L g654 ( 
.A(n_630),
.B(n_246),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_563),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_558),
.Y(n_656)
);

NAND2x1p5_ASAP7_75t_L g657 ( 
.A(n_591),
.B(n_363),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_563),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_558),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_613),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_582),
.B(n_549),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_568),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_558),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_591),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_568),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_568),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_633),
.B(n_466),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_579),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_576),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_591),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_558),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_579),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_561),
.Y(n_674)
);

INVx5_ASAP7_75t_L g675 ( 
.A(n_561),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_585),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_579),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_585),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_576),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_559),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_585),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_639),
.B(n_466),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_635),
.A2(n_623),
.B1(n_631),
.B2(n_645),
.Y(n_683)
);

XOR2xp5_ASAP7_75t_L g684 ( 
.A(n_613),
.B(n_444),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_576),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_561),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_630),
.B(n_246),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_598),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_585),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_633),
.B(n_578),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_599),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_578),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_576),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_639),
.B(n_534),
.Y(n_694)
);

INVxp67_ASAP7_75t_SL g695 ( 
.A(n_566),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_561),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_576),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_640),
.B(n_470),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_625),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_640),
.B(n_470),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_599),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_592),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_561),
.Y(n_704)
);

AOI21x1_ASAP7_75t_L g705 ( 
.A1(n_559),
.A2(n_302),
.B(n_299),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_566),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_599),
.Y(n_707)
);

AOI22xp33_ASAP7_75t_L g708 ( 
.A1(n_631),
.A2(n_493),
.B1(n_364),
.B2(n_226),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_599),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_596),
.Y(n_710)
);

AND2x2_ASAP7_75t_SL g711 ( 
.A(n_632),
.B(n_245),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_601),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_601),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_638),
.B(n_471),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_557),
.B(n_299),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_584),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_638),
.B(n_471),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_598),
.Y(n_718)
);

BUFx4f_ASAP7_75t_L g719 ( 
.A(n_638),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_647),
.B(n_542),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_561),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_601),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_635),
.A2(n_364),
.B1(n_420),
.B2(n_252),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_590),
.B(n_327),
.C(n_302),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_560),
.Y(n_725)
);

CKINVDCx6p67_ASAP7_75t_R g726 ( 
.A(n_575),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_647),
.B(n_545),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_625),
.Y(n_728)
);

HB1xp67_ASAP7_75t_L g729 ( 
.A(n_564),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_632),
.B(n_556),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_638),
.B(n_644),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_569),
.Y(n_732)
);

BUFx4f_ASAP7_75t_L g733 ( 
.A(n_638),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_648),
.B(n_546),
.Y(n_734)
);

BUFx4f_ASAP7_75t_L g735 ( 
.A(n_638),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_627),
.B(n_476),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_569),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_564),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_596),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_557),
.B(n_327),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_608),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_644),
.B(n_646),
.Y(n_742)
);

INVx1_ASAP7_75t_SL g743 ( 
.A(n_565),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_627),
.B(n_476),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_648),
.B(n_555),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_569),
.Y(n_747)
);

NAND3xp33_ASAP7_75t_L g748 ( 
.A(n_590),
.B(n_359),
.C(n_347),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_601),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_560),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_562),
.Y(n_751)
);

BUFx10_ASAP7_75t_L g752 ( 
.A(n_644),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_562),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_557),
.B(n_481),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_557),
.B(n_481),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_644),
.B(n_483),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_634),
.A2(n_420),
.B1(n_252),
.B2(n_343),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_567),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_567),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_L g760 ( 
.A(n_593),
.B(n_359),
.C(n_347),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_634),
.B(n_245),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_648),
.B(n_483),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_565),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_644),
.B(n_491),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_569),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_571),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_644),
.B(n_646),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_584),
.Y(n_769)
);

CKINVDCx6p67_ASAP7_75t_R g770 ( 
.A(n_646),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_634),
.A2(n_588),
.B1(n_589),
.B2(n_612),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_569),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_646),
.B(n_491),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_645),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_569),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_610),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_566),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_571),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_592),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_612),
.B(n_492),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_610),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_592),
.Y(n_782)
);

XOR2xp5_ASAP7_75t_L g783 ( 
.A(n_605),
.B(n_448),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_574),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_646),
.B(n_492),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_L g786 ( 
.A1(n_645),
.A2(n_315),
.B1(n_433),
.B2(n_276),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_610),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_646),
.B(n_497),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_610),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_574),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_566),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_618),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_618),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_618),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_612),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_612),
.Y(n_796)
);

INVxp67_ASAP7_75t_SL g797 ( 
.A(n_570),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_620),
.B(n_497),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_603),
.A2(n_543),
.B1(n_527),
.B2(n_605),
.Y(n_799)
);

BUFx10_ASAP7_75t_L g800 ( 
.A(n_634),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_618),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_592),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_SL g803 ( 
.A1(n_603),
.A2(n_469),
.B1(n_489),
.B2(n_452),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_573),
.B(n_604),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_621),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_690),
.B(n_573),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_738),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_738),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_762),
.B(n_604),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_692),
.B(n_771),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_762),
.B(n_620),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_762),
.B(n_620),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_774),
.B(n_588),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_690),
.B(n_641),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_791),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_711),
.B(n_719),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_738),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_711),
.B(n_620),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_729),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_SL g820 ( 
.A(n_741),
.B(n_603),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_804),
.A2(n_617),
.B1(n_595),
.B2(n_572),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_795),
.A2(n_796),
.B(n_733),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_688),
.B(n_572),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_680),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_711),
.A2(n_460),
.B1(n_477),
.B2(n_467),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_680),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_692),
.A2(n_636),
.B1(n_589),
.B2(n_626),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_719),
.B(n_733),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_795),
.B(n_641),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_725),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_699),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_796),
.B(n_626),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_725),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_752),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_736),
.B(n_581),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_744),
.B(n_581),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_715),
.B(n_586),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_699),
.B(n_593),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_699),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_719),
.B(n_412),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_763),
.Y(n_841)
);

O2A1O1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_668),
.A2(n_606),
.B(n_609),
.C(n_586),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_791),
.Y(n_843)
);

AND2x2_ASAP7_75t_SL g844 ( 
.A(n_768),
.B(n_313),
.Y(n_844)
);

INVx6_ASAP7_75t_L g845 ( 
.A(n_752),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_715),
.B(n_606),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_733),
.B(n_412),
.Y(n_847)
);

NAND2xp33_ASAP7_75t_L g848 ( 
.A(n_657),
.B(n_412),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_715),
.A2(n_636),
.B1(n_621),
.B2(n_325),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_715),
.B(n_609),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_740),
.B(n_611),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_740),
.B(n_611),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_735),
.B(n_412),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_728),
.B(n_594),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_728),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_735),
.B(n_412),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_SL g857 ( 
.A(n_743),
.B(n_603),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_740),
.B(n_616),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_735),
.B(n_616),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_752),
.B(n_628),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_710),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_740),
.A2(n_636),
.B1(n_621),
.B2(n_325),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_754),
.B(n_374),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_728),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_752),
.B(n_628),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_652),
.B(n_621),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_654),
.A2(n_313),
.B1(n_391),
.B2(n_387),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_676),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_652),
.B(n_592),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_800),
.B(n_710),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_661),
.B(n_614),
.Y(n_871)
);

BUFx8_ASAP7_75t_L g872 ( 
.A(n_739),
.Y(n_872)
);

AND2x6_ASAP7_75t_SL g873 ( 
.A(n_694),
.B(n_250),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_800),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_750),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_661),
.B(n_665),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_750),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_800),
.B(n_643),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_676),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_678),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_678),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_751),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_751),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_681),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_L g885 ( 
.A(n_657),
.B(n_387),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_730),
.B(n_391),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_800),
.B(n_643),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_665),
.B(n_614),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_753),
.Y(n_889)
);

NAND2x1_ASAP7_75t_L g890 ( 
.A(n_671),
.B(n_570),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_739),
.B(n_595),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_654),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_671),
.B(n_614),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_718),
.B(n_614),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_SL g895 ( 
.A1(n_783),
.A2(n_484),
.B1(n_501),
.B2(n_480),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_682),
.B(n_500),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_681),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_698),
.B(n_500),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_683),
.B(n_614),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_657),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_726),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_753),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_734),
.B(n_642),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_755),
.Y(n_904)
);

NAND3xp33_ASAP7_75t_L g905 ( 
.A(n_683),
.B(n_513),
.C(n_506),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_689),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_764),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_691),
.B(n_506),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_691),
.B(n_513),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_758),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_702),
.B(n_515),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_770),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_702),
.B(n_515),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_707),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_780),
.A2(n_402),
.B1(n_424),
.B2(n_392),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_700),
.B(n_516),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_731),
.B(n_742),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_798),
.B(n_318),
.Y(n_918)
);

INVx8_ASAP7_75t_L g919 ( 
.A(n_654),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_707),
.B(n_516),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_654),
.A2(n_431),
.B1(n_424),
.B2(n_392),
.Y(n_921)
);

OR2x6_ASAP7_75t_L g922 ( 
.A(n_714),
.B(n_374),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_758),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_662),
.B(n_530),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_709),
.B(n_530),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_709),
.B(n_421),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_712),
.B(n_533),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_720),
.B(n_533),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_788),
.A2(n_539),
.B1(n_554),
.B2(n_551),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_654),
.A2(n_394),
.B1(n_431),
.B2(n_397),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_712),
.B(n_713),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_713),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_727),
.B(n_536),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_770),
.A2(n_757),
.B1(n_717),
.B2(n_756),
.Y(n_934)
);

NAND2x1_ASAP7_75t_L g935 ( 
.A(n_659),
.B(n_570),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_759),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_746),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_765),
.B(n_536),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_708),
.B(n_642),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_722),
.B(n_422),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_695),
.A2(n_570),
.B(n_587),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_773),
.B(n_539),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_722),
.B(n_548),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_785),
.A2(n_394),
.B1(n_417),
.B2(n_397),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_684),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_749),
.B(n_776),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_660),
.B(n_548),
.Y(n_947)
);

AND2x6_ASAP7_75t_SL g948 ( 
.A(n_684),
.B(n_265),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_749),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_776),
.B(n_550),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_654),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_781),
.B(n_550),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_759),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_781),
.B(n_551),
.Y(n_954)
);

AOI22xp33_ASAP7_75t_L g955 ( 
.A1(n_654),
.A2(n_402),
.B1(n_405),
.B2(n_417),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_767),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_787),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_787),
.B(n_554),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_786),
.B(n_556),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_789),
.B(n_577),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_789),
.B(n_577),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_792),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_792),
.B(n_580),
.Y(n_963)
);

INVxp33_ASAP7_75t_L g964 ( 
.A(n_783),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_793),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_793),
.B(n_580),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_794),
.B(n_801),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_794),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_791),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_649),
.B(n_405),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_801),
.B(n_587),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_767),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_724),
.Y(n_973)
);

AOI22xp33_ASAP7_75t_L g974 ( 
.A1(n_687),
.A2(n_649),
.B1(n_784),
.B2(n_778),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_805),
.B(n_587),
.Y(n_975)
);

AOI22xp33_ASAP7_75t_L g976 ( 
.A1(n_687),
.A2(n_629),
.B1(n_622),
.B2(n_624),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_835),
.B(n_805),
.Y(n_977)
);

O2A1O1Ixp5_ASAP7_75t_L g978 ( 
.A1(n_816),
.A2(n_705),
.B(n_784),
.C(n_778),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_828),
.A2(n_797),
.B(n_706),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_814),
.B(n_836),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_834),
.B(n_791),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_876),
.A2(n_871),
.B(n_869),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_842),
.A2(n_724),
.B(n_760),
.C(n_748),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_806),
.B(n_687),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_868),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_900),
.A2(n_723),
.B1(n_799),
.B2(n_790),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_828),
.A2(n_802),
.B(n_703),
.Y(n_987)
);

AO21x1_ASAP7_75t_L g988 ( 
.A1(n_816),
.A2(n_705),
.B(n_703),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_834),
.A2(n_802),
.B(n_703),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_841),
.B(n_687),
.Y(n_990)
);

OR2x2_ASAP7_75t_L g991 ( 
.A(n_907),
.B(n_637),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_824),
.Y(n_992)
);

OAI21xp5_ASAP7_75t_L g993 ( 
.A1(n_888),
.A2(n_687),
.B(n_790),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_903),
.B(n_629),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_834),
.A2(n_802),
.B(n_703),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_819),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_848),
.A2(n_802),
.B(n_693),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_824),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_823),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_809),
.A2(n_597),
.B(n_600),
.C(n_594),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_826),
.Y(n_1001)
);

NAND2xp33_ASAP7_75t_L g1002 ( 
.A(n_874),
.B(n_687),
.Y(n_1002)
);

CKINVDCx8_ASAP7_75t_R g1003 ( 
.A(n_948),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_837),
.B(n_679),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_848),
.A2(n_693),
.B(n_670),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_893),
.A2(n_866),
.B(n_885),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_885),
.A2(n_693),
.B(n_670),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_811),
.A2(n_693),
.B(n_670),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_829),
.B(n_687),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_811),
.A2(n_670),
.B(n_745),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_809),
.A2(n_600),
.B(n_602),
.C(n_597),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_826),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_812),
.A2(n_779),
.B(n_745),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_810),
.A2(n_748),
.B(n_760),
.C(n_637),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_864),
.B(n_602),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_937),
.B(n_803),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_830),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_812),
.A2(n_779),
.B(n_745),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_899),
.A2(n_615),
.B(n_607),
.C(n_619),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_830),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_813),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_L g1022 ( 
.A(n_905),
.B(n_290),
.C(n_236),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_822),
.A2(n_782),
.B(n_779),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_833),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_833),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_875),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_956),
.B(n_782),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_939),
.B(n_726),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_810),
.A2(n_959),
.B(n_928),
.C(n_933),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_875),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_879),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_956),
.B(n_659),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_917),
.A2(n_656),
.B(n_653),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_831),
.B(n_659),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_938),
.A2(n_380),
.B(n_378),
.C(n_437),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_846),
.A2(n_656),
.B(n_653),
.Y(n_1036)
);

INVx6_ASAP7_75t_L g1037 ( 
.A(n_872),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_864),
.B(n_607),
.Y(n_1038)
);

AO21x1_ASAP7_75t_L g1039 ( 
.A1(n_818),
.A2(n_685),
.B(n_679),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_899),
.A2(n_619),
.B(n_624),
.C(n_615),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_808),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_877),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_839),
.B(n_659),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_973),
.A2(n_769),
.B(n_761),
.C(n_716),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_855),
.B(n_664),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_850),
.A2(n_852),
.B(n_851),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_818),
.A2(n_685),
.B(n_679),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_943),
.A2(n_761),
.B(n_716),
.C(n_769),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_858),
.B(n_685),
.Y(n_1049)
);

NAND2x1p5_ASAP7_75t_L g1050 ( 
.A(n_874),
.B(n_697),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_859),
.A2(n_772),
.B(n_701),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_859),
.A2(n_701),
.B(n_697),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_808),
.B(n_622),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_880),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_838),
.B(n_854),
.Y(n_1055)
);

OAI21xp33_ASAP7_75t_L g1056 ( 
.A1(n_827),
.A2(n_346),
.B(n_345),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_838),
.B(n_854),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_838),
.B(n_664),
.Y(n_1058)
);

NAND2xp33_ASAP7_75t_L g1059 ( 
.A(n_874),
.B(n_772),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_874),
.B(n_697),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_844),
.A2(n_656),
.B(n_653),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_881),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_877),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_884),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_844),
.A2(n_656),
.B(n_653),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_815),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_815),
.Y(n_1067)
);

AND2x6_ASAP7_75t_L g1068 ( 
.A(n_892),
.B(n_772),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_919),
.A2(n_672),
.B(n_653),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_919),
.A2(n_686),
.B(n_672),
.Y(n_1070)
);

BUFx4f_ASAP7_75t_L g1071 ( 
.A(n_922),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_904),
.A2(n_701),
.B1(n_674),
.B2(n_696),
.Y(n_1072)
);

AO21x1_ASAP7_75t_L g1073 ( 
.A1(n_840),
.A2(n_266),
.B(n_265),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_931),
.A2(n_761),
.B(n_716),
.Y(n_1074)
);

NAND2x1_ASAP7_75t_L g1075 ( 
.A(n_845),
.B(n_664),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_919),
.A2(n_686),
.B(n_672),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_890),
.A2(n_673),
.B(n_669),
.Y(n_1077)
);

AO21x1_ASAP7_75t_L g1078 ( 
.A1(n_840),
.A2(n_282),
.B(n_266),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_919),
.A2(n_686),
.B(n_672),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_886),
.A2(n_358),
.B1(n_432),
.B2(n_353),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_860),
.A2(n_686),
.B(n_672),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_854),
.B(n_664),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_897),
.Y(n_1083)
);

INVx11_ASAP7_75t_L g1084 ( 
.A(n_872),
.Y(n_1084)
);

OAI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_946),
.A2(n_769),
.B(n_673),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_894),
.B(n_674),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_906),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_860),
.A2(n_721),
.B(n_686),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_891),
.B(n_674),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_896),
.A2(n_622),
.B(n_669),
.C(n_677),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_815),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_914),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_865),
.A2(n_775),
.B(n_721),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_847),
.A2(n_398),
.B(n_419),
.C(n_426),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_943),
.A2(n_954),
.B(n_918),
.C(n_934),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_865),
.A2(n_775),
.B(n_721),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_967),
.A2(n_677),
.B(n_650),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_832),
.A2(n_853),
.B(n_847),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_843),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_932),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_853),
.A2(n_775),
.B(n_721),
.Y(n_1101)
);

INVx2_ASAP7_75t_SL g1102 ( 
.A(n_861),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_807),
.B(n_674),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_901),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_843),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_825),
.B(n_891),
.C(n_947),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_882),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_856),
.A2(n_775),
.B(n_721),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_924),
.B(n_351),
.C(n_348),
.Y(n_1109)
);

AO21x1_ASAP7_75t_L g1110 ( 
.A1(n_856),
.A2(n_286),
.B(n_282),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_817),
.B(n_696),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_949),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_870),
.A2(n_704),
.B(n_696),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_870),
.A2(n_912),
.B(n_971),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_843),
.A2(n_969),
.B(n_941),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_957),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_845),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_962),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_912),
.A2(n_845),
.B(n_908),
.Y(n_1119)
);

A2O1A1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_886),
.A2(n_344),
.B(n_426),
.C(n_337),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_912),
.A2(n_704),
.B(n_696),
.Y(n_1121)
);

INVxp67_ASAP7_75t_L g1122 ( 
.A(n_954),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_976),
.B(n_704),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_898),
.A2(n_732),
.B(n_766),
.C(n_747),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_849),
.B(n_732),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_916),
.A2(n_732),
.B1(n_766),
.B2(n_747),
.Y(n_1126)
);

AOI21x1_ASAP7_75t_L g1127 ( 
.A1(n_975),
.A2(n_935),
.B(n_960),
.Y(n_1127)
);

INVx11_ASAP7_75t_L g1128 ( 
.A(n_872),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_862),
.B(n_732),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_909),
.B(n_737),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_911),
.B(n_737),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_942),
.B(n_340),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_913),
.B(n_737),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_970),
.A2(n_337),
.B1(n_322),
.B2(n_316),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_975),
.A2(n_963),
.B(n_961),
.Y(n_1135)
);

OAI21xp33_ASAP7_75t_L g1136 ( 
.A1(n_821),
.A2(n_356),
.B(n_355),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_969),
.B(n_737),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_920),
.A2(n_766),
.B(n_747),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_882),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_L g1140 ( 
.A(n_922),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_892),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_925),
.B(n_747),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_927),
.A2(n_766),
.B(n_675),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_950),
.B(n_655),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_952),
.A2(n_675),
.B(n_651),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_965),
.Y(n_1146)
);

CKINVDCx6p67_ASAP7_75t_R g1147 ( 
.A(n_922),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_958),
.B(n_655),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_968),
.B(n_658),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_883),
.B(n_658),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_918),
.B(n_360),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_969),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_974),
.A2(n_650),
.B(n_663),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_878),
.B(n_366),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_820),
.B(n_296),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_951),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_889),
.B(n_663),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_889),
.B(n_666),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_966),
.A2(n_675),
.B(n_651),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_926),
.A2(n_343),
.B(n_280),
.C(n_666),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_878),
.B(n_375),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_902),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_926),
.A2(n_280),
.B(n_322),
.C(n_419),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_902),
.B(n_777),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_940),
.A2(n_384),
.B(n_301),
.C(n_316),
.Y(n_1165)
);

AND2x2_ASAP7_75t_SL g1166 ( 
.A(n_921),
.B(n_286),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_895),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_L g1168 ( 
.A(n_980),
.B(n_887),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1046),
.A2(n_997),
.B(n_1005),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_994),
.B(n_929),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1029),
.A2(n_944),
.B(n_915),
.C(n_922),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_1104),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1002),
.A2(n_951),
.B(n_867),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1007),
.A2(n_955),
.B(n_930),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1141),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1141),
.Y(n_1176)
);

AOI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1106),
.A2(n_863),
.B1(n_887),
.B2(n_940),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_996),
.Y(n_1178)
);

NOR2xp67_ASAP7_75t_SL g1179 ( 
.A(n_1117),
.B(n_910),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_1102),
.Y(n_1180)
);

INVx5_ASAP7_75t_L g1181 ( 
.A(n_1068),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1029),
.A2(n_863),
.B(n_970),
.C(n_972),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_SL g1183 ( 
.A(n_1167),
.B(n_857),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1037),
.B(n_945),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1055),
.A2(n_863),
.B1(n_972),
.B2(n_953),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1162),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1006),
.A2(n_923),
.B(n_910),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_984),
.A2(n_936),
.B(n_923),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_985),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_977),
.B(n_936),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_982),
.A2(n_953),
.B(n_863),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1031),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_992),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_999),
.B(n_964),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1054),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1106),
.A2(n_970),
.B1(n_964),
.B2(n_303),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1021),
.B(n_297),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1037),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_1141),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1141),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1057),
.A2(n_1122),
.B1(n_999),
.B2(n_1156),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1014),
.A2(n_970),
.B(n_398),
.C(n_301),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_977),
.B(n_667),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_998),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_991),
.B(n_583),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1095),
.A2(n_344),
.B(n_349),
.C(n_353),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1037),
.B(n_349),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1062),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1001),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1021),
.B(n_300),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1051),
.A2(n_650),
.B(n_667),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1156),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1115),
.A2(n_1077),
.B(n_1033),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1122),
.B(n_873),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1064),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1012),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1009),
.A2(n_675),
.B(n_651),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1156),
.A2(n_328),
.B1(n_308),
.B2(n_314),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1152),
.B(n_583),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1152),
.B(n_777),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1008),
.A2(n_675),
.B(n_651),
.Y(n_1221)
);

AOI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1060),
.A2(n_378),
.B(n_358),
.Y(n_1222)
);

AO21x1_ASAP7_75t_L g1223 ( 
.A1(n_1098),
.A2(n_365),
.B(n_380),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1109),
.A2(n_303),
.B1(n_321),
.B2(n_323),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1016),
.B(n_382),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1017),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1144),
.B(n_777),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1156),
.A2(n_352),
.B1(n_333),
.B2(n_336),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1148),
.B(n_777),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1020),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1151),
.A2(n_365),
.B(n_384),
.C(n_430),
.Y(n_1231)
);

AO22x1_ASAP7_75t_L g1232 ( 
.A1(n_1016),
.A2(n_389),
.B1(n_388),
.B2(n_436),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1083),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_993),
.A2(n_675),
.B(n_651),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1087),
.B(n_777),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1024),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1109),
.A2(n_303),
.B1(n_339),
.B2(n_362),
.Y(n_1237)
);

BUFx4f_ASAP7_75t_L g1238 ( 
.A(n_1147),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1092),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1071),
.B(n_354),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1154),
.B(n_383),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1028),
.B(n_393),
.Y(n_1242)
);

BUFx12f_ASAP7_75t_L g1243 ( 
.A(n_1015),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1036),
.A2(n_651),
.B(n_777),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1100),
.B(n_357),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1112),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1116),
.B(n_369),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_1151),
.A2(n_418),
.B1(n_395),
.B2(n_407),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1154),
.A2(n_437),
.B(n_430),
.C(n_432),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_L g1250 ( 
.A1(n_1161),
.A2(n_434),
.B(n_371),
.C(n_425),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1118),
.B(n_370),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1161),
.B(n_396),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1146),
.B(n_372),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_981),
.A2(n_381),
.B(n_423),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1080),
.B(n_385),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1071),
.B(n_386),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1025),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1117),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_981),
.A2(n_399),
.B(n_416),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1026),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_990),
.A2(n_404),
.B1(n_413),
.B2(n_410),
.Y(n_1261)
);

NOR2xp67_ASAP7_75t_SL g1262 ( 
.A(n_1119),
.B(n_427),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1030),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_989),
.A2(n_156),
.B(n_103),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_995),
.A2(n_1059),
.B(n_1010),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1140),
.B(n_400),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1042),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1080),
.B(n_401),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1140),
.B(n_1015),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1061),
.A2(n_155),
.B(n_104),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1066),
.B(n_408),
.Y(n_1271)
);

NAND3xp33_ASAP7_75t_SL g1272 ( 
.A(n_1022),
.B(n_403),
.C(n_10),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1066),
.B(n_1067),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1063),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1107),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_SL g1276 ( 
.A1(n_1120),
.A2(n_222),
.B(n_216),
.C(n_215),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1053),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_978),
.A2(n_211),
.B(n_202),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1065),
.A2(n_201),
.B(n_195),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1041),
.B(n_8),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_1041),
.Y(n_1281)
);

AND2x2_ASAP7_75t_SL g1282 ( 
.A(n_1166),
.B(n_16),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_987),
.A2(n_171),
.B(n_166),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1067),
.B(n_151),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1123),
.A2(n_147),
.B1(n_142),
.B2(n_126),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_978),
.A2(n_124),
.B(n_113),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_986),
.A2(n_110),
.B1(n_108),
.B2(n_97),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1086),
.A2(n_83),
.B(n_18),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1091),
.B(n_17),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1091),
.B(n_19),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1139),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1099),
.B(n_1105),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1099),
.Y(n_1293)
);

OAI22x1_ASAP7_75t_L g1294 ( 
.A1(n_1132),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_1294)
);

INVx3_ASAP7_75t_L g1295 ( 
.A(n_1105),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1069),
.A2(n_83),
.B(n_25),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1070),
.A2(n_81),
.B(n_26),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1038),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1068),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1038),
.B(n_21),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1130),
.B(n_28),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_R g1302 ( 
.A(n_1003),
.B(n_79),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1053),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1125),
.A2(n_29),
.B(n_31),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1155),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1131),
.B(n_1133),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1068),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1076),
.A2(n_29),
.B(n_32),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1142),
.B(n_33),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1136),
.B(n_33),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1079),
.A2(n_79),
.B(n_36),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1075),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1050),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1089),
.B(n_35),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1058),
.B(n_35),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1155),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1149),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1050),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_1068),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1120),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1150),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1157),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1089),
.B(n_1004),
.Y(n_1323)
);

O2A1O1Ixp5_ASAP7_75t_L g1324 ( 
.A1(n_988),
.A2(n_1114),
.B(n_1039),
.C(n_983),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1004),
.A2(n_76),
.B(n_39),
.Y(n_1325)
);

AOI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1022),
.A2(n_37),
.B1(n_39),
.B2(n_42),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1049),
.A2(n_43),
.B(n_44),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_1056),
.Y(n_1328)
);

INVx3_ASAP7_75t_L g1329 ( 
.A(n_1068),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1082),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1049),
.A2(n_44),
.B(n_45),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1084),
.B(n_46),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1035),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1013),
.A2(n_52),
.B(n_53),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1166),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1213),
.A2(n_1052),
.B(n_1047),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1281),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1211),
.A2(n_1023),
.B(n_1113),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1205),
.B(n_1134),
.Y(n_1339)
);

OAI22x1_ASAP7_75t_L g1340 ( 
.A1(n_1241),
.A2(n_1072),
.B1(n_1126),
.B2(n_1060),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1317),
.B(n_1027),
.Y(n_1341)
);

AOI221x1_ASAP7_75t_L g1342 ( 
.A1(n_1304),
.A2(n_1252),
.B1(n_1334),
.B2(n_1278),
.C(n_1286),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1194),
.B(n_1011),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1189),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1192),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1170),
.B(n_1134),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1169),
.A2(n_1018),
.B(n_979),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1265),
.A2(n_1074),
.B(n_1085),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1180),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1243),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1174),
.A2(n_1097),
.B(n_1129),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1195),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1208),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1322),
.B(n_1040),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1215),
.Y(n_1355)
);

O2A1O1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1225),
.A2(n_1035),
.B(n_1000),
.C(n_1165),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1214),
.B(n_1305),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1172),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1306),
.A2(n_1124),
.B(n_1093),
.Y(n_1359)
);

AOI221x1_ASAP7_75t_L g1360 ( 
.A1(n_1334),
.A2(n_1090),
.B1(n_1138),
.B2(n_1160),
.C(n_1096),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1191),
.A2(n_1168),
.B(n_1306),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1233),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1239),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1303),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1324),
.A2(n_1153),
.B(n_1088),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1223),
.A2(n_1073),
.A3(n_1110),
.B(n_1078),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1182),
.A2(n_1044),
.B(n_1081),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1321),
.B(n_1019),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1173),
.A2(n_1158),
.B(n_1143),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_SL g1370 ( 
.A(n_1178),
.B(n_1163),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1246),
.Y(n_1371)
);

CKINVDCx20_ASAP7_75t_R g1372 ( 
.A(n_1316),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1186),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1257),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1188),
.A2(n_1187),
.B(n_1221),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1219),
.B(n_1032),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1219),
.B(n_1103),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1193),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1323),
.A2(n_1121),
.B(n_1137),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_SL g1380 ( 
.A1(n_1206),
.A2(n_1164),
.B(n_1137),
.C(n_1045),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1323),
.A2(n_1048),
.B(n_1135),
.Y(n_1381)
);

INVxp67_ASAP7_75t_L g1382 ( 
.A(n_1280),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1181),
.A2(n_1101),
.B(n_1108),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1181),
.A2(n_1145),
.B(n_1111),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1204),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_SL g1386 ( 
.A1(n_1314),
.A2(n_1164),
.B(n_1043),
.C(n_1034),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1330),
.B(n_1127),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1330),
.B(n_1159),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1234),
.A2(n_1094),
.B(n_1128),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1175),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1184),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1181),
.A2(n_1094),
.B(n_63),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1209),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1269),
.B(n_61),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1181),
.A2(n_65),
.B(n_68),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1171),
.A2(n_69),
.B(n_1314),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1217),
.A2(n_69),
.B(n_1244),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1227),
.A2(n_1229),
.B(n_1185),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_1310),
.B(n_1224),
.C(n_1237),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1177),
.A2(n_1202),
.B(n_1328),
.C(n_1287),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1249),
.A2(n_1231),
.B(n_1268),
.C(n_1325),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1284),
.A2(n_1250),
.B(n_1290),
.C(n_1289),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1203),
.A2(n_1190),
.B(n_1222),
.Y(n_1403)
);

XOR2xp5_ASAP7_75t_L g1404 ( 
.A(n_1201),
.B(n_1240),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1203),
.A2(n_1190),
.B(n_1284),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_1299),
.B(n_1307),
.Y(n_1406)
);

AO32x2_ASAP7_75t_L g1407 ( 
.A1(n_1285),
.A2(n_1261),
.A3(n_1307),
.B1(n_1299),
.B2(n_1319),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1216),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1226),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1301),
.A2(n_1309),
.B(n_1227),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_1315),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1270),
.A2(n_1279),
.B(n_1283),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1229),
.A2(n_1319),
.B(n_1264),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1183),
.A2(n_1242),
.B1(n_1282),
.B2(n_1266),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1196),
.B(n_1315),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1301),
.A2(n_1309),
.B(n_1292),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1273),
.A2(n_1292),
.B(n_1220),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1268),
.A2(n_1255),
.B(n_1331),
.C(n_1327),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1260),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1273),
.A2(n_1258),
.B(n_1312),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1258),
.A2(n_1312),
.B(n_1210),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1276),
.A2(n_1255),
.B(n_1271),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1198),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1230),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1272),
.A2(n_1300),
.B(n_1320),
.C(n_1333),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1298),
.Y(n_1426)
);

OR2x2_ASAP7_75t_L g1427 ( 
.A(n_1271),
.B(n_1184),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1184),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1267),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1330),
.B(n_1263),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1327),
.A2(n_1331),
.B(n_1290),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1275),
.Y(n_1432)
);

O2A1O1Ixp5_ASAP7_75t_L g1433 ( 
.A1(n_1262),
.A2(n_1256),
.B(n_1297),
.C(n_1308),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1236),
.B(n_1274),
.Y(n_1434)
);

AOI21xp33_ASAP7_75t_L g1435 ( 
.A1(n_1248),
.A2(n_1289),
.B(n_1335),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1175),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1296),
.A2(n_1311),
.B(n_1288),
.C(n_1326),
.Y(n_1437)
);

INVx5_ASAP7_75t_L g1438 ( 
.A(n_1175),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1179),
.A2(n_1259),
.B(n_1254),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1245),
.B(n_1247),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1220),
.A2(n_1329),
.B(n_1313),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1291),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1207),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1207),
.Y(n_1444)
);

AO31x2_ASAP7_75t_L g1445 ( 
.A1(n_1294),
.A2(n_1235),
.A3(n_1253),
.B(n_1251),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1207),
.Y(n_1446)
);

OR2x6_ASAP7_75t_L g1447 ( 
.A(n_1277),
.B(n_1176),
.Y(n_1447)
);

NOR4xp25_ASAP7_75t_L g1448 ( 
.A(n_1245),
.B(n_1247),
.C(n_1253),
.D(n_1251),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1232),
.B(n_1197),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1238),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1199),
.B(n_1295),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1199),
.B(n_1295),
.Y(n_1452)
);

AOI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1235),
.A2(n_1228),
.B(n_1218),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1332),
.B(n_1277),
.C(n_1293),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1277),
.B(n_1293),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1176),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1329),
.A2(n_1313),
.B(n_1318),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1318),
.A2(n_1176),
.B(n_1200),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1200),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1200),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1212),
.A2(n_1238),
.B(n_1302),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1212),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1212),
.A2(n_733),
.B(n_719),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1213),
.A2(n_1211),
.B(n_1051),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1324),
.A2(n_1046),
.B(n_1029),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1324),
.A2(n_1046),
.B(n_1029),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1241),
.B(n_937),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1213),
.A2(n_1211),
.B(n_1051),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1213),
.A2(n_1211),
.B(n_1051),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1213),
.A2(n_1211),
.B(n_1051),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_SL g1471 ( 
.A1(n_1206),
.A2(n_1029),
.B(n_1014),
.C(n_1120),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1223),
.A2(n_1206),
.A3(n_1191),
.B(n_1039),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1194),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1282),
.A2(n_980),
.B1(n_1029),
.B2(n_1080),
.Y(n_1474)
);

A2O1A1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1241),
.A2(n_1029),
.B(n_1252),
.C(n_1095),
.Y(n_1475)
);

A2O1A1Ixp33_ASAP7_75t_L g1476 ( 
.A1(n_1241),
.A2(n_1029),
.B(n_1252),
.C(n_1095),
.Y(n_1476)
);

A2O1A1Ixp33_ASAP7_75t_L g1477 ( 
.A1(n_1241),
.A2(n_1029),
.B(n_1252),
.C(n_1095),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1324),
.A2(n_1046),
.B(n_1029),
.Y(n_1478)
);

BUFx2_ASAP7_75t_L g1479 ( 
.A(n_1281),
.Y(n_1479)
);

O2A1O1Ixp33_ASAP7_75t_SL g1480 ( 
.A1(n_1206),
.A2(n_1029),
.B(n_1014),
.C(n_1120),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1317),
.B(n_980),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1169),
.A2(n_733),
.B(n_719),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1169),
.A2(n_733),
.B(n_719),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1189),
.Y(n_1484)
);

AO31x2_ASAP7_75t_L g1485 ( 
.A1(n_1223),
.A2(n_1206),
.A3(n_1191),
.B(n_1039),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1170),
.B(n_994),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1317),
.B(n_980),
.Y(n_1487)
);

O2A1O1Ixp33_ASAP7_75t_SL g1488 ( 
.A1(n_1206),
.A2(n_1029),
.B(n_1014),
.C(n_1120),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1169),
.A2(n_733),
.B(n_719),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1169),
.A2(n_733),
.B(n_719),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1170),
.B(n_994),
.Y(n_1491)
);

CKINVDCx8_ASAP7_75t_R g1492 ( 
.A(n_1172),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1324),
.A2(n_1191),
.B(n_1213),
.Y(n_1493)
);

INVx3_ASAP7_75t_SL g1494 ( 
.A(n_1172),
.Y(n_1494)
);

BUFx12f_ASAP7_75t_L g1495 ( 
.A(n_1172),
.Y(n_1495)
);

AO22x2_ASAP7_75t_L g1496 ( 
.A1(n_1304),
.A2(n_1106),
.B1(n_1314),
.B2(n_1286),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1189),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1182),
.A2(n_1202),
.B(n_1327),
.Y(n_1498)
);

BUFx2_ASAP7_75t_L g1499 ( 
.A(n_1281),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1317),
.B(n_980),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1213),
.A2(n_1211),
.B(n_1051),
.Y(n_1501)
);

AOI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1191),
.A2(n_828),
.B(n_1187),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1194),
.B(n_980),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1189),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1241),
.A2(n_1252),
.B1(n_1225),
.B2(n_928),
.Y(n_1505)
);

CKINVDCx20_ASAP7_75t_R g1506 ( 
.A(n_1172),
.Y(n_1506)
);

AOI31xp67_ASAP7_75t_L g1507 ( 
.A1(n_1177),
.A2(n_816),
.A3(n_828),
.B(n_859),
.Y(n_1507)
);

BUFx5_ASAP7_75t_L g1508 ( 
.A(n_1322),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1194),
.B(n_980),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1170),
.B(n_994),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1317),
.B(n_980),
.Y(n_1511)
);

AO31x2_ASAP7_75t_L g1512 ( 
.A1(n_1223),
.A2(n_1206),
.A3(n_1191),
.B(n_1039),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1467),
.A2(n_1399),
.B1(n_1474),
.B2(n_1505),
.Y(n_1513)
);

INVx6_ASAP7_75t_L g1514 ( 
.A(n_1438),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1353),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1484),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1474),
.A2(n_1435),
.B1(n_1396),
.B2(n_1440),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1506),
.Y(n_1518)
);

BUFx12f_ASAP7_75t_L g1519 ( 
.A(n_1358),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1492),
.Y(n_1520)
);

BUFx2_ASAP7_75t_SL g1521 ( 
.A(n_1349),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1344),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_L g1523 ( 
.A1(n_1475),
.A2(n_1477),
.B(n_1476),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1486),
.B(n_1491),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1345),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1435),
.A2(n_1396),
.B1(n_1415),
.B2(n_1404),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1449),
.A2(n_1496),
.B1(n_1510),
.B2(n_1346),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1372),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1348),
.A2(n_1361),
.B(n_1482),
.Y(n_1529)
);

INVx2_ASAP7_75t_SL g1530 ( 
.A(n_1438),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1496),
.A2(n_1394),
.B1(n_1503),
.B2(n_1509),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1414),
.A2(n_1357),
.B1(n_1382),
.B2(n_1411),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1423),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1496),
.A2(n_1394),
.B1(n_1343),
.B2(n_1339),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1438),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1406),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1411),
.A2(n_1473),
.B1(n_1427),
.B2(n_1498),
.Y(n_1537)
);

CKINVDCx6p67_ASAP7_75t_R g1538 ( 
.A(n_1494),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1443),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1370),
.A2(n_1428),
.B1(n_1391),
.B2(n_1431),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1479),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1431),
.A2(n_1446),
.B1(n_1444),
.B2(n_1511),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1447),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1481),
.A2(n_1511),
.B1(n_1487),
.B2(n_1500),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1406),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1481),
.A2(n_1500),
.B1(n_1487),
.B2(n_1342),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1352),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1459),
.Y(n_1548)
);

BUFx4_ASAP7_75t_SL g1549 ( 
.A(n_1462),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1495),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1461),
.A2(n_1454),
.B1(n_1465),
.B2(n_1466),
.Y(n_1551)
);

BUFx4_ASAP7_75t_SL g1552 ( 
.A(n_1426),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1461),
.A2(n_1478),
.B1(n_1465),
.B2(n_1466),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1478),
.A2(n_1508),
.B1(n_1499),
.B2(n_1340),
.Y(n_1554)
);

BUFx2_ASAP7_75t_SL g1555 ( 
.A(n_1450),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1508),
.A2(n_1364),
.B1(n_1337),
.B2(n_1422),
.Y(n_1556)
);

BUFx4f_ASAP7_75t_L g1557 ( 
.A(n_1459),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1508),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1508),
.Y(n_1559)
);

CKINVDCx11_ASAP7_75t_R g1560 ( 
.A(n_1350),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1400),
.A2(n_1337),
.B1(n_1364),
.B2(n_1341),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1508),
.A2(n_1422),
.B1(n_1354),
.B2(n_1410),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1355),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1362),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1354),
.A2(n_1410),
.B1(n_1388),
.B2(n_1368),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1363),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1388),
.A2(n_1368),
.B1(n_1395),
.B2(n_1424),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1401),
.A2(n_1418),
.B1(n_1448),
.B2(n_1455),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1457),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1378),
.A2(n_1408),
.B1(n_1409),
.B2(n_1393),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1371),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1385),
.A2(n_1419),
.B1(n_1432),
.B2(n_1374),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1429),
.A2(n_1442),
.B1(n_1430),
.B2(n_1341),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1497),
.Y(n_1574)
);

OAI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1377),
.A2(n_1376),
.B1(n_1504),
.B2(n_1430),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1456),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1377),
.A2(n_1416),
.B1(n_1373),
.B2(n_1376),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1434),
.Y(n_1578)
);

BUFx3_ASAP7_75t_L g1579 ( 
.A(n_1459),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_SL g1580 ( 
.A1(n_1392),
.A2(n_1425),
.B1(n_1361),
.B2(n_1412),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1447),
.Y(n_1581)
);

CKINVDCx11_ASAP7_75t_R g1582 ( 
.A(n_1447),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1416),
.A2(n_1421),
.B1(n_1434),
.B2(n_1387),
.Y(n_1583)
);

BUFx10_ASAP7_75t_L g1584 ( 
.A(n_1460),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1471),
.A2(n_1480),
.B1(n_1488),
.B2(n_1367),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1403),
.Y(n_1586)
);

INVx6_ASAP7_75t_L g1587 ( 
.A(n_1390),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1367),
.A2(n_1387),
.B1(n_1365),
.B2(n_1356),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1451),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1441),
.Y(n_1590)
);

INVx8_ASAP7_75t_L g1591 ( 
.A(n_1390),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1417),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1451),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1452),
.A2(n_1379),
.B1(n_1381),
.B2(n_1351),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1452),
.A2(n_1420),
.B1(n_1453),
.B2(n_1413),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1398),
.A2(n_1436),
.B1(n_1381),
.B2(n_1360),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1458),
.Y(n_1597)
);

BUFx4f_ASAP7_75t_SL g1598 ( 
.A(n_1507),
.Y(n_1598)
);

BUFx8_ASAP7_75t_SL g1599 ( 
.A(n_1439),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1365),
.A2(n_1359),
.B1(n_1405),
.B2(n_1369),
.Y(n_1600)
);

CKINVDCx11_ASAP7_75t_R g1601 ( 
.A(n_1445),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1397),
.A2(n_1493),
.B1(n_1389),
.B2(n_1347),
.Y(n_1602)
);

BUFx8_ASAP7_75t_SL g1603 ( 
.A(n_1502),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1437),
.A2(n_1482),
.B1(n_1483),
.B2(n_1463),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1493),
.B(n_1336),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1483),
.A2(n_1490),
.B1(n_1489),
.B2(n_1384),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1347),
.A2(n_1383),
.B(n_1445),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1445),
.B(n_1402),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1380),
.A2(n_1386),
.B1(n_1375),
.B2(n_1338),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1407),
.A2(n_1433),
.B1(n_1512),
.B2(n_1485),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1366),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1366),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1472),
.B(n_1512),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1472),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1366),
.Y(n_1615)
);

AO22x1_ASAP7_75t_L g1616 ( 
.A1(n_1407),
.A2(n_1485),
.B1(n_1512),
.B2(n_1469),
.Y(n_1616)
);

OAI22x1_ASAP7_75t_SL g1617 ( 
.A1(n_1407),
.A2(n_1464),
.B1(n_1468),
.B2(n_1470),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1501),
.A2(n_1241),
.B1(n_1252),
.B2(n_1282),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1337),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1505),
.A2(n_1241),
.B1(n_1252),
.B2(n_1225),
.Y(n_1621)
);

CKINVDCx11_ASAP7_75t_R g1622 ( 
.A(n_1492),
.Y(n_1622)
);

OAI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1505),
.A2(n_1467),
.B1(n_1414),
.B2(n_1399),
.Y(n_1623)
);

CKINVDCx5p33_ASAP7_75t_R g1624 ( 
.A(n_1506),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1625)
);

BUFx10_ASAP7_75t_L g1626 ( 
.A(n_1358),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1438),
.Y(n_1631)
);

CKINVDCx11_ASAP7_75t_R g1632 ( 
.A(n_1492),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1353),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1353),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_1349),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1353),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1638)
);

INVx6_ASAP7_75t_L g1639 ( 
.A(n_1438),
.Y(n_1639)
);

INVx4_ASAP7_75t_L g1640 ( 
.A(n_1438),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1358),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1353),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1479),
.Y(n_1643)
);

INVx5_ASAP7_75t_L g1644 ( 
.A(n_1447),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1353),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1406),
.Y(n_1646)
);

INVx8_ASAP7_75t_L g1647 ( 
.A(n_1438),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1506),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1438),
.Y(n_1651)
);

BUFx12f_ASAP7_75t_L g1652 ( 
.A(n_1358),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_SL g1653 ( 
.A1(n_1467),
.A2(n_1241),
.B1(n_1252),
.B2(n_1282),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1353),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1353),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1506),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1353),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1406),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1467),
.A2(n_1241),
.B1(n_1252),
.B2(n_1282),
.Y(n_1662)
);

CKINVDCx11_ASAP7_75t_R g1663 ( 
.A(n_1492),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1505),
.A2(n_1467),
.B1(n_999),
.B2(n_1225),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1353),
.Y(n_1665)
);

BUFx3_ASAP7_75t_L g1666 ( 
.A(n_1349),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1353),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1506),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1337),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1505),
.B(n_1467),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1353),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1505),
.A2(n_1467),
.B1(n_999),
.B2(n_1225),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1438),
.Y(n_1674)
);

CKINVDCx11_ASAP7_75t_R g1675 ( 
.A(n_1492),
.Y(n_1675)
);

BUFx12f_ASAP7_75t_L g1676 ( 
.A(n_1358),
.Y(n_1676)
);

INVx6_ASAP7_75t_L g1677 ( 
.A(n_1438),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1353),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1353),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1505),
.A2(n_1467),
.B1(n_1414),
.B2(n_1399),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1505),
.A2(n_1252),
.B(n_1241),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1486),
.B(n_1491),
.Y(n_1682)
);

CKINVDCx6p67_ASAP7_75t_R g1683 ( 
.A(n_1494),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1353),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1685)
);

OAI21xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1505),
.A2(n_1225),
.B(n_803),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_L g1687 ( 
.A1(n_1505),
.A2(n_1399),
.B1(n_1241),
.B2(n_1252),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1353),
.Y(n_1688)
);

AOI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1616),
.A2(n_1529),
.B(n_1606),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1611),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1612),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1615),
.Y(n_1692)
);

OA21x2_ASAP7_75t_L g1693 ( 
.A1(n_1607),
.A2(n_1608),
.B(n_1600),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1681),
.A2(n_1653),
.B1(n_1662),
.B2(n_1621),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1586),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1620),
.A2(n_1629),
.B1(n_1687),
.B2(n_1685),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1592),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1520),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1569),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1544),
.B(n_1625),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1592),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1569),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1614),
.Y(n_1704)
);

BUFx3_ASAP7_75t_L g1705 ( 
.A(n_1603),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1669),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1613),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1590),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1603),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1590),
.Y(n_1710)
);

CKINVDCx11_ASAP7_75t_R g1711 ( 
.A(n_1520),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1590),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1605),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1584),
.Y(n_1714)
);

HB1xp67_ASAP7_75t_L g1715 ( 
.A(n_1619),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1543),
.Y(n_1716)
);

BUFx2_ASAP7_75t_L g1717 ( 
.A(n_1599),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1569),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1513),
.A2(n_1670),
.B1(n_1656),
.B2(n_1638),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1589),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1527),
.B(n_1523),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1593),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1617),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1598),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1522),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1536),
.B(n_1545),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1525),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1536),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1547),
.Y(n_1729)
);

CKINVDCx6p67_ASAP7_75t_R g1730 ( 
.A(n_1622),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1536),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1561),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1563),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1643),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1564),
.Y(n_1735)
);

INVx2_ASAP7_75t_L g1736 ( 
.A(n_1566),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1571),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1574),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1568),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1516),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1604),
.A2(n_1602),
.B(n_1609),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1543),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1584),
.Y(n_1743)
);

BUFx2_ASAP7_75t_L g1744 ( 
.A(n_1599),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1553),
.B(n_1534),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1628),
.B(n_1630),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1517),
.B(n_1526),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1634),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1644),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1637),
.Y(n_1750)
);

OAI21x1_ASAP7_75t_L g1751 ( 
.A1(n_1594),
.A2(n_1562),
.B(n_1583),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1524),
.B(n_1682),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1541),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1637),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1545),
.Y(n_1755)
);

CKINVDCx14_ASAP7_75t_R g1756 ( 
.A(n_1622),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1655),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1543),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1655),
.B(n_1658),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1658),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1636),
.A2(n_1650),
.B1(n_1660),
.B2(n_1649),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1661),
.A2(n_1673),
.B1(n_1627),
.B2(n_1686),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1665),
.Y(n_1763)
);

OA21x2_ASAP7_75t_L g1764 ( 
.A1(n_1556),
.A2(n_1554),
.B(n_1565),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1678),
.B(n_1679),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1664),
.B(n_1672),
.Y(n_1766)
);

OA21x2_ASAP7_75t_L g1767 ( 
.A1(n_1577),
.A2(n_1531),
.B(n_1567),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1578),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1515),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1541),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1551),
.B(n_1588),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1601),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1644),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1601),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1576),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1633),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1610),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1596),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1642),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1644),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1688),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1645),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1644),
.Y(n_1783)
);

OAI21x1_ASAP7_75t_L g1784 ( 
.A1(n_1540),
.A2(n_1659),
.B(n_1646),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1646),
.B(n_1659),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1654),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1667),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1684),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1671),
.Y(n_1789)
);

OAI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1623),
.A2(n_1680),
.B1(n_1532),
.B2(n_1683),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1542),
.B(n_1537),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1644),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1584),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1597),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1573),
.B(n_1585),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1659),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1575),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1546),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1572),
.B(n_1618),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1514),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1595),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1570),
.B(n_1580),
.Y(n_1802)
);

CKINVDCx20_ASAP7_75t_R g1803 ( 
.A(n_1632),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1530),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1631),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1631),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1651),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1651),
.Y(n_1808)
);

BUFx4f_ASAP7_75t_SL g1809 ( 
.A(n_1519),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1535),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1548),
.B(n_1581),
.Y(n_1811)
);

INVx1_ASAP7_75t_SL g1812 ( 
.A(n_1582),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1535),
.Y(n_1813)
);

BUFx4f_ASAP7_75t_SL g1814 ( 
.A(n_1519),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1581),
.B(n_1528),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1535),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1548),
.B(n_1579),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1579),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1647),
.A2(n_1640),
.B(n_1514),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1548),
.B(n_1582),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1528),
.B(n_1518),
.Y(n_1821)
);

OAI21x1_ASAP7_75t_L g1822 ( 
.A1(n_1647),
.A2(n_1514),
.B(n_1639),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1674),
.Y(n_1823)
);

BUFx12f_ASAP7_75t_L g1824 ( 
.A(n_1711),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1701),
.B(n_1518),
.Y(n_1825)
);

OAI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1746),
.A2(n_1557),
.B(n_1533),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1797),
.B(n_1548),
.Y(n_1827)
);

AOI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1719),
.A2(n_1539),
.B1(n_1560),
.B2(n_1538),
.Y(n_1828)
);

OAI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1694),
.A2(n_1539),
.B1(n_1538),
.B2(n_1683),
.Y(n_1829)
);

OA21x2_ASAP7_75t_L g1830 ( 
.A1(n_1741),
.A2(n_1550),
.B(n_1647),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1719),
.B(n_1624),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1726),
.B(n_1635),
.Y(n_1832)
);

OAI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1741),
.A2(n_1647),
.B(n_1677),
.Y(n_1833)
);

OA21x2_ASAP7_75t_L g1834 ( 
.A1(n_1801),
.A2(n_1550),
.B(n_1639),
.Y(n_1834)
);

AO32x2_ASAP7_75t_L g1835 ( 
.A1(n_1762),
.A2(n_1560),
.A3(n_1555),
.B1(n_1587),
.B2(n_1552),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1803),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1727),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1752),
.B(n_1648),
.Y(n_1838)
);

A2O1A1Ixp33_ASAP7_75t_L g1839 ( 
.A1(n_1761),
.A2(n_1557),
.B(n_1635),
.C(n_1666),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1772),
.B(n_1626),
.Y(n_1840)
);

BUFx4f_ASAP7_75t_SL g1841 ( 
.A(n_1730),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1772),
.B(n_1626),
.Y(n_1842)
);

OR2x6_ASAP7_75t_L g1843 ( 
.A(n_1749),
.B(n_1677),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1774),
.B(n_1753),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1790),
.A2(n_1666),
.B(n_1549),
.C(n_1521),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1774),
.B(n_1753),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1706),
.B(n_1657),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1811),
.B(n_1587),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1745),
.B(n_1657),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1745),
.B(n_1820),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1797),
.B(n_1674),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1820),
.B(n_1624),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1706),
.B(n_1668),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1735),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1737),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1697),
.A2(n_1668),
.B1(n_1674),
.B2(n_1675),
.C(n_1663),
.Y(n_1856)
);

OAI211xp5_ASAP7_75t_SL g1857 ( 
.A1(n_1761),
.A2(n_1663),
.B(n_1675),
.C(n_1652),
.Y(n_1857)
);

AO32x2_ASAP7_75t_L g1858 ( 
.A1(n_1714),
.A2(n_1591),
.A3(n_1641),
.B1(n_1676),
.B2(n_1743),
.Y(n_1858)
);

OAI21x1_ASAP7_75t_SL g1859 ( 
.A1(n_1799),
.A2(n_1676),
.B(n_1591),
.Y(n_1859)
);

AND2x4_ASAP7_75t_L g1860 ( 
.A(n_1726),
.B(n_1785),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1720),
.B(n_1722),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1787),
.B(n_1771),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1766),
.A2(n_1747),
.B(n_1739),
.C(n_1721),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1725),
.B(n_1729),
.Y(n_1864)
);

INVx4_ASAP7_75t_L g1865 ( 
.A(n_1716),
.Y(n_1865)
);

AO32x2_ASAP7_75t_L g1866 ( 
.A1(n_1743),
.A2(n_1793),
.A3(n_1800),
.B1(n_1777),
.B2(n_1798),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1720),
.B(n_1722),
.Y(n_1867)
);

HB1xp67_ASAP7_75t_L g1868 ( 
.A(n_1775),
.Y(n_1868)
);

A2O1A1Ixp33_ASAP7_75t_L g1869 ( 
.A1(n_1739),
.A2(n_1721),
.B(n_1771),
.C(n_1709),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1751),
.A2(n_1732),
.B(n_1802),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1791),
.B(n_1817),
.Y(n_1871)
);

NAND2x1_ASAP7_75t_L g1872 ( 
.A(n_1794),
.B(n_1728),
.Y(n_1872)
);

AO32x2_ASAP7_75t_L g1873 ( 
.A1(n_1793),
.A2(n_1800),
.A3(n_1777),
.B1(n_1798),
.B2(n_1778),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1756),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_L g1875 ( 
.A(n_1815),
.B(n_1821),
.Y(n_1875)
);

O2A1O1Ixp33_ASAP7_75t_SL g1876 ( 
.A1(n_1812),
.A2(n_1723),
.B(n_1734),
.C(n_1770),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_SL g1877 ( 
.A(n_1794),
.B(n_1749),
.Y(n_1877)
);

AO21x2_ASAP7_75t_L g1878 ( 
.A1(n_1689),
.A2(n_1801),
.B(n_1778),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1699),
.B(n_1715),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1768),
.B(n_1794),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1791),
.B(n_1817),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1795),
.A2(n_1723),
.B1(n_1734),
.B2(n_1802),
.C(n_1717),
.Y(n_1882)
);

AOI211xp5_ASAP7_75t_L g1883 ( 
.A1(n_1717),
.A2(n_1744),
.B(n_1709),
.C(n_1705),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1726),
.B(n_1785),
.Y(n_1884)
);

OAI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1744),
.A2(n_1795),
.B(n_1709),
.C(n_1705),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1738),
.Y(n_1886)
);

A2O1A1Ixp33_ASAP7_75t_L g1887 ( 
.A1(n_1705),
.A2(n_1751),
.B(n_1784),
.C(n_1724),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1804),
.B(n_1805),
.Y(n_1888)
);

OAI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1812),
.A2(n_1764),
.B1(n_1730),
.B2(n_1767),
.Y(n_1889)
);

CKINVDCx20_ASAP7_75t_R g1890 ( 
.A(n_1809),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1725),
.B(n_1729),
.Y(n_1891)
);

CKINVDCx5p33_ASAP7_75t_R g1892 ( 
.A(n_1814),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1784),
.A2(n_1724),
.B(n_1822),
.C(n_1819),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1733),
.B(n_1736),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1779),
.A2(n_1788),
.B1(n_1781),
.B2(n_1738),
.C(n_1707),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1726),
.B(n_1785),
.Y(n_1896)
);

O2A1O1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1767),
.A2(n_1764),
.B(n_1724),
.C(n_1781),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1768),
.B(n_1707),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1767),
.A2(n_1764),
.B(n_1689),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1767),
.A2(n_1764),
.B1(n_1758),
.B2(n_1742),
.Y(n_1900)
);

NOR2x1_ASAP7_75t_SL g1901 ( 
.A(n_1749),
.B(n_1773),
.Y(n_1901)
);

OAI21x1_ASAP7_75t_L g1902 ( 
.A1(n_1819),
.A2(n_1822),
.B(n_1700),
.Y(n_1902)
);

AOI221xp5_ASAP7_75t_L g1903 ( 
.A1(n_1779),
.A2(n_1788),
.B1(n_1776),
.B2(n_1789),
.C(n_1769),
.Y(n_1903)
);

A2O1A1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1716),
.A2(n_1758),
.B(n_1742),
.C(n_1792),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1760),
.B(n_1740),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1759),
.B(n_1765),
.Y(n_1906)
);

OAI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1700),
.A2(n_1703),
.B(n_1713),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1690),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_1818),
.Y(n_1909)
);

INVx4_ASAP7_75t_L g1910 ( 
.A(n_1742),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1690),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1691),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1758),
.A2(n_1810),
.B1(n_1813),
.B2(n_1816),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1769),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1740),
.B(n_1750),
.Y(n_1915)
);

OAI211xp5_ASAP7_75t_L g1916 ( 
.A1(n_1782),
.A2(n_1786),
.B(n_1789),
.C(n_1693),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1893),
.B(n_1713),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1871),
.B(n_1693),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1868),
.B(n_1782),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1908),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1911),
.Y(n_1921)
);

INVxp67_ASAP7_75t_L g1922 ( 
.A(n_1881),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1862),
.B(n_1693),
.Y(n_1923)
);

OR2x2_ASAP7_75t_L g1924 ( 
.A(n_1864),
.B(n_1891),
.Y(n_1924)
);

AND2x2_ASAP7_75t_SL g1925 ( 
.A(n_1834),
.B(n_1693),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1912),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1866),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1906),
.B(n_1713),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1828),
.A2(n_1749),
.B1(n_1773),
.B2(n_1780),
.Y(n_1929)
);

OR2x2_ASAP7_75t_L g1930 ( 
.A(n_1880),
.B(n_1708),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1829),
.A2(n_1780),
.B1(n_1749),
.B2(n_1773),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1866),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1837),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1854),
.Y(n_1934)
);

OR2x6_ASAP7_75t_L g1935 ( 
.A(n_1833),
.B(n_1749),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1914),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1855),
.Y(n_1937)
);

INVx4_ASAP7_75t_R g1938 ( 
.A(n_1852),
.Y(n_1938)
);

OAI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1829),
.A2(n_1856),
.B1(n_1831),
.B2(n_1882),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1894),
.Y(n_1940)
);

INVx1_ASAP7_75t_SL g1941 ( 
.A(n_1847),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1850),
.B(n_1710),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1880),
.B(n_1710),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1870),
.B(n_1786),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1886),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1844),
.B(n_1846),
.Y(n_1946)
);

NOR2xp33_ASAP7_75t_L g1947 ( 
.A(n_1825),
.B(n_1785),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1905),
.B(n_1712),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1905),
.B(n_1712),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1870),
.B(n_1786),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1888),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1872),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1860),
.B(n_1718),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1861),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1856),
.A2(n_1780),
.B1(n_1773),
.B2(n_1783),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1884),
.B(n_1718),
.Y(n_1956)
);

OAI222xp33_ASAP7_75t_L g1957 ( 
.A1(n_1889),
.A2(n_1805),
.B1(n_1807),
.B2(n_1808),
.C1(n_1804),
.C2(n_1806),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1896),
.B(n_1718),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1902),
.B(n_1700),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1896),
.B(n_1698),
.Y(n_1960)
);

BUFx4f_ASAP7_75t_SL g1961 ( 
.A(n_1824),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1861),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1863),
.B(n_1789),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1834),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1867),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1889),
.B(n_1696),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1867),
.Y(n_1967)
);

BUFx2_ASAP7_75t_L g1968 ( 
.A(n_1866),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1915),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1873),
.B(n_1698),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1915),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1882),
.B(n_1696),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1857),
.A2(n_1796),
.B1(n_1755),
.B2(n_1731),
.Y(n_1973)
);

AND2x4_ASAP7_75t_L g1974 ( 
.A(n_1964),
.B(n_1901),
.Y(n_1974)
);

OR2x2_ASAP7_75t_L g1975 ( 
.A(n_1918),
.B(n_1878),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1918),
.B(n_1907),
.Y(n_1976)
);

INVxp67_ASAP7_75t_SL g1977 ( 
.A(n_1963),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1952),
.Y(n_1978)
);

OR2x2_ASAP7_75t_L g1979 ( 
.A(n_1924),
.B(n_1878),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1924),
.B(n_1899),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1959),
.Y(n_1981)
);

AOI211xp5_ASAP7_75t_SL g1982 ( 
.A1(n_1939),
.A2(n_1885),
.B(n_1887),
.C(n_1876),
.Y(n_1982)
);

AOI21xp33_ASAP7_75t_L g1983 ( 
.A1(n_1955),
.A2(n_1897),
.B(n_1845),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1923),
.B(n_1946),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1929),
.A2(n_1857),
.B1(n_1849),
.B2(n_1900),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1927),
.B(n_1899),
.Y(n_1986)
);

BUFx3_ASAP7_75t_L g1987 ( 
.A(n_1961),
.Y(n_1987)
);

INVx4_ASAP7_75t_L g1988 ( 
.A(n_1951),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1922),
.B(n_1895),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1936),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1920),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1936),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1964),
.Y(n_1993)
);

INVx1_ASAP7_75t_SL g1994 ( 
.A(n_1941),
.Y(n_1994)
);

INVxp67_ASAP7_75t_L g1995 ( 
.A(n_1919),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1927),
.B(n_1916),
.Y(n_1996)
);

OAI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1931),
.A2(n_1869),
.B(n_1845),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1954),
.B(n_1895),
.Y(n_1998)
);

AOI33xp33_ASAP7_75t_L g1999 ( 
.A1(n_1954),
.A2(n_1883),
.A3(n_1897),
.B1(n_1842),
.B2(n_1840),
.B3(n_1853),
.Y(n_1999)
);

AOI221x1_ASAP7_75t_L g2000 ( 
.A1(n_1972),
.A2(n_1826),
.B1(n_1839),
.B2(n_1913),
.C(n_1879),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1920),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1936),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1953),
.B(n_1830),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1932),
.B(n_1916),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1930),
.Y(n_2005)
);

OAI33xp33_ASAP7_75t_L g2006 ( 
.A1(n_1944),
.A2(n_1827),
.A3(n_1898),
.B1(n_1851),
.B2(n_1692),
.B3(n_1909),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1921),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1932),
.B(n_1830),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1964),
.Y(n_2009)
);

AOI31xp67_ASAP7_75t_L g2010 ( 
.A1(n_1917),
.A2(n_1702),
.A3(n_1704),
.B(n_1695),
.Y(n_2010)
);

INVx2_ASAP7_75t_SL g2011 ( 
.A(n_1951),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1959),
.B(n_1877),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1959),
.B(n_1904),
.Y(n_2013)
);

AOI211xp5_ASAP7_75t_SL g2014 ( 
.A1(n_1957),
.A2(n_1885),
.B(n_1966),
.C(n_1950),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1921),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1956),
.B(n_1873),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_1959),
.B(n_1843),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1958),
.B(n_1873),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1935),
.B(n_1917),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1926),
.Y(n_2020)
);

OAI33xp33_ASAP7_75t_L g2021 ( 
.A1(n_1962),
.A2(n_1827),
.A3(n_1851),
.B1(n_1692),
.B2(n_1754),
.B3(n_1748),
.Y(n_2021)
);

INVxp67_ASAP7_75t_SL g2022 ( 
.A(n_1943),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1947),
.B(n_1875),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1942),
.B(n_1838),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1928),
.B(n_1835),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1965),
.B(n_1903),
.Y(n_2026)
);

OAI221xp5_ASAP7_75t_L g2027 ( 
.A1(n_1973),
.A2(n_1826),
.B1(n_1874),
.B2(n_1865),
.C(n_1910),
.Y(n_2027)
);

NAND4xp25_ASAP7_75t_L g2028 ( 
.A(n_1968),
.B(n_1903),
.C(n_1763),
.D(n_1757),
.Y(n_2028)
);

AOI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1925),
.A2(n_1841),
.B1(n_1832),
.B2(n_1848),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1977),
.B(n_1967),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1998),
.B(n_2026),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1976),
.B(n_1968),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1991),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_2010),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_2010),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1976),
.B(n_2003),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1996),
.B(n_1971),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2003),
.B(n_1925),
.Y(n_2038)
);

INVx3_ASAP7_75t_L g2039 ( 
.A(n_2019),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1996),
.B(n_1971),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1979),
.Y(n_2041)
);

OR2x2_ASAP7_75t_L g2042 ( 
.A(n_2004),
.B(n_1948),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1979),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1993),
.B(n_1925),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1991),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2001),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1990),
.Y(n_2047)
);

AND2x4_ASAP7_75t_L g2048 ( 
.A(n_2019),
.B(n_1917),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1993),
.B(n_1970),
.Y(n_2049)
);

OAI33xp33_ASAP7_75t_L g2050 ( 
.A1(n_2004),
.A2(n_1967),
.A3(n_1934),
.B1(n_1933),
.B2(n_1937),
.B3(n_1945),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_1986),
.B(n_1949),
.Y(n_2051)
);

AND2x2_ASAP7_75t_SL g2052 ( 
.A(n_1999),
.B(n_1917),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1980),
.Y(n_2053)
);

INVxp67_ASAP7_75t_SL g2054 ( 
.A(n_2008),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_2019),
.B(n_2012),
.Y(n_2055)
);

AND2x2_ASAP7_75t_L g2056 ( 
.A(n_2009),
.B(n_1970),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2007),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_2019),
.B(n_1935),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2015),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1986),
.B(n_1949),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2009),
.B(n_1940),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2015),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1980),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1990),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_1975),
.B(n_1969),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2016),
.B(n_2018),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2020),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2016),
.B(n_2018),
.Y(n_2068)
);

INVx1_ASAP7_75t_SL g2069 ( 
.A(n_1978),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1992),
.Y(n_2070)
);

AOI221x1_ASAP7_75t_L g2071 ( 
.A1(n_1997),
.A2(n_1813),
.B1(n_1810),
.B2(n_1816),
.C(n_1823),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_1978),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2002),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1984),
.B(n_1960),
.Y(n_2074)
);

OAI32xp33_ASAP7_75t_L g2075 ( 
.A1(n_2031),
.A2(n_2008),
.A3(n_2069),
.B1(n_2053),
.B2(n_2063),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2055),
.B(n_2066),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2055),
.B(n_2013),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2033),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2031),
.B(n_2014),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_2052),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2042),
.B(n_1975),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2052),
.B(n_1989),
.Y(n_2082)
);

INVx1_ASAP7_75t_SL g2083 ( 
.A(n_2052),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2042),
.B(n_2005),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2052),
.B(n_1994),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2030),
.B(n_1995),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2055),
.B(n_2013),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2033),
.Y(n_2088)
);

NAND2x1_ASAP7_75t_L g2089 ( 
.A(n_2055),
.B(n_1938),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2033),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2034),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2030),
.B(n_2022),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2045),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2034),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2042),
.B(n_2037),
.Y(n_2095)
);

OAI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_2071),
.A2(n_1982),
.B(n_2000),
.Y(n_2096)
);

NOR2x1p5_ASAP7_75t_L g2097 ( 
.A(n_2039),
.B(n_1987),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2055),
.B(n_2013),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2034),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2055),
.B(n_2013),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_2034),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2037),
.B(n_2005),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2074),
.B(n_2025),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_2048),
.B(n_1987),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2066),
.B(n_2025),
.Y(n_2105)
);

AOI32xp33_ASAP7_75t_L g2106 ( 
.A1(n_2044),
.A2(n_1985),
.A3(n_2027),
.B1(n_2023),
.B2(n_2000),
.Y(n_2106)
);

INVx1_ASAP7_75t_SL g2107 ( 
.A(n_2069),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2037),
.B(n_2040),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_2044),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2045),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2074),
.B(n_2024),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2066),
.B(n_2012),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2048),
.B(n_2058),
.Y(n_2113)
);

OAI21xp5_ASAP7_75t_L g2114 ( 
.A1(n_2071),
.A2(n_1983),
.B(n_2029),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2045),
.Y(n_2115)
);

NOR2x1p5_ASAP7_75t_L g2116 ( 
.A(n_2039),
.B(n_1892),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_2048),
.B(n_1890),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2068),
.B(n_2012),
.Y(n_2118)
);

NOR2xp33_ASAP7_75t_SL g2119 ( 
.A(n_2050),
.B(n_2006),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2068),
.B(n_2012),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2068),
.B(n_2017),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2039),
.B(n_2017),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2039),
.B(n_2017),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_2035),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2046),
.Y(n_2125)
);

INVx2_ASAP7_75t_SL g2126 ( 
.A(n_2097),
.Y(n_2126)
);

AOI221x1_ASAP7_75t_L g2127 ( 
.A1(n_2096),
.A2(n_1988),
.B1(n_2028),
.B2(n_2044),
.C(n_2067),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2078),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2091),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2082),
.B(n_2053),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2080),
.B(n_2063),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2091),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2076),
.B(n_2048),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2076),
.B(n_2048),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2078),
.Y(n_2135)
);

INVxp67_ASAP7_75t_SL g2136 ( 
.A(n_2091),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2097),
.B(n_2048),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2088),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2121),
.B(n_2058),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2121),
.B(n_2058),
.Y(n_2140)
);

HB1xp67_ASAP7_75t_L g2141 ( 
.A(n_2107),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2088),
.Y(n_2142)
);

OR2x2_ASAP7_75t_L g2143 ( 
.A(n_2103),
.B(n_2051),
.Y(n_2143)
);

AND3x2_ASAP7_75t_L g2144 ( 
.A(n_2119),
.B(n_2072),
.C(n_2054),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2090),
.Y(n_2145)
);

HB1xp67_ASAP7_75t_L g2146 ( 
.A(n_2095),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2083),
.B(n_2054),
.Y(n_2147)
);

INVxp67_ASAP7_75t_SL g2148 ( 
.A(n_2094),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2112),
.B(n_2058),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2094),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2079),
.B(n_2071),
.C(n_2072),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2094),
.Y(n_2152)
);

INVx1_ASAP7_75t_SL g2153 ( 
.A(n_2085),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2090),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2093),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2095),
.B(n_2051),
.Y(n_2156)
);

AND2x4_ASAP7_75t_L g2157 ( 
.A(n_2112),
.B(n_2058),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2099),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2093),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_2108),
.B(n_2051),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2110),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2119),
.B(n_2032),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2086),
.B(n_2032),
.Y(n_2163)
);

NAND2xp33_ASAP7_75t_L g2164 ( 
.A(n_2106),
.B(n_2029),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2110),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2146),
.Y(n_2166)
);

NAND2x1_ASAP7_75t_L g2167 ( 
.A(n_2126),
.B(n_2113),
.Y(n_2167)
);

OAI22xp5_ASAP7_75t_L g2168 ( 
.A1(n_2162),
.A2(n_2106),
.B1(n_2151),
.B2(n_2114),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_SL g2169 ( 
.A1(n_2127),
.A2(n_2116),
.B(n_2104),
.Y(n_2169)
);

AOI22x1_ASAP7_75t_L g2170 ( 
.A1(n_2141),
.A2(n_2116),
.B1(n_2109),
.B2(n_2075),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2128),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2139),
.B(n_2118),
.Y(n_2172)
);

OAI22xp5_ASAP7_75t_L g2173 ( 
.A1(n_2162),
.A2(n_2089),
.B1(n_2105),
.B2(n_2111),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2144),
.B(n_2105),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_2151),
.B(n_2117),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2139),
.B(n_2118),
.Y(n_2176)
);

AOI22xp5_ASAP7_75t_L g2177 ( 
.A1(n_2164),
.A2(n_2089),
.B1(n_2113),
.B2(n_2100),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2129),
.Y(n_2178)
);

NAND2xp33_ASAP7_75t_SL g2179 ( 
.A(n_2126),
.B(n_1836),
.Y(n_2179)
);

OAI32xp33_ASAP7_75t_L g2180 ( 
.A1(n_2153),
.A2(n_2108),
.A3(n_2081),
.B1(n_2039),
.B2(n_2075),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2128),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2126),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2135),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2135),
.Y(n_2184)
);

OAI211xp5_ASAP7_75t_L g2185 ( 
.A1(n_2127),
.A2(n_2077),
.B(n_2087),
.C(n_2098),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2138),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_L g2187 ( 
.A1(n_2153),
.A2(n_2113),
.B1(n_2120),
.B2(n_2039),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2138),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2142),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2129),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2142),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2145),
.Y(n_2192)
);

OAI22xp5_ASAP7_75t_L g2193 ( 
.A1(n_2163),
.A2(n_2113),
.B1(n_2120),
.B2(n_2058),
.Y(n_2193)
);

AOI31xp33_ASAP7_75t_L g2194 ( 
.A1(n_2130),
.A2(n_2087),
.A3(n_2077),
.B(n_2098),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2167),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_2166),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2182),
.B(n_2130),
.Y(n_2197)
);

AND2x2_ASAP7_75t_L g2198 ( 
.A(n_2172),
.B(n_2137),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_2168),
.B(n_2131),
.Y(n_2199)
);

AOI222xp33_ASAP7_75t_L g2200 ( 
.A1(n_2175),
.A2(n_2147),
.B1(n_2131),
.B2(n_2163),
.C1(n_2137),
.C2(n_2050),
.Y(n_2200)
);

OAI221xp5_ASAP7_75t_L g2201 ( 
.A1(n_2175),
.A2(n_2147),
.B1(n_2156),
.B2(n_2160),
.C(n_2143),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2172),
.B(n_2140),
.Y(n_2202)
);

NAND3x2_ASAP7_75t_L g2203 ( 
.A(n_2170),
.B(n_2156),
.C(n_2160),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_2179),
.A2(n_2157),
.B1(n_2134),
.B2(n_2133),
.Y(n_2204)
);

AND2x2_ASAP7_75t_SL g2205 ( 
.A(n_2174),
.B(n_2133),
.Y(n_2205)
);

AOI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2180),
.A2(n_2165),
.B1(n_2161),
.B2(n_2159),
.C(n_2145),
.Y(n_2206)
);

AOI21xp33_ASAP7_75t_SL g2207 ( 
.A1(n_2170),
.A2(n_2143),
.B(n_2134),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2176),
.B(n_2140),
.Y(n_2208)
);

HB1xp67_ASAP7_75t_L g2209 ( 
.A(n_2167),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2176),
.B(n_2149),
.Y(n_2210)
);

INVx3_ASAP7_75t_SL g2211 ( 
.A(n_2179),
.Y(n_2211)
);

OAI32xp33_ASAP7_75t_L g2212 ( 
.A1(n_2173),
.A2(n_2169),
.A3(n_2187),
.B1(n_2193),
.B2(n_2191),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2177),
.B(n_2149),
.Y(n_2213)
);

INVxp67_ASAP7_75t_L g2214 ( 
.A(n_2171),
.Y(n_2214)
);

INVx1_ASAP7_75t_SL g2215 ( 
.A(n_2181),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2183),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2194),
.B(n_2157),
.Y(n_2217)
);

OAI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2203),
.A2(n_2207),
.B(n_2199),
.Y(n_2218)
);

AO22x2_ASAP7_75t_L g2219 ( 
.A1(n_2215),
.A2(n_2192),
.B1(n_2184),
.B2(n_2189),
.Y(n_2219)
);

NAND2x1p5_ASAP7_75t_L g2220 ( 
.A(n_2204),
.B(n_2178),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2195),
.Y(n_2221)
);

OAI21xp33_ASAP7_75t_L g2222 ( 
.A1(n_2212),
.A2(n_2169),
.B(n_2185),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2209),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2205),
.B(n_2157),
.Y(n_2224)
);

BUFx3_ASAP7_75t_L g2225 ( 
.A(n_2211),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2205),
.B(n_2157),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2196),
.B(n_2186),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2211),
.A2(n_2217),
.B1(n_2200),
.B2(n_2213),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2196),
.Y(n_2229)
);

OAI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2201),
.A2(n_2188),
.B1(n_2092),
.B2(n_2081),
.C(n_2148),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2198),
.B(n_2100),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2197),
.B(n_2178),
.Y(n_2232)
);

OAI211xp5_ASAP7_75t_L g2233 ( 
.A1(n_2222),
.A2(n_2206),
.B(n_2214),
.C(n_2216),
.Y(n_2233)
);

OAI21xp33_ASAP7_75t_SL g2234 ( 
.A1(n_2218),
.A2(n_2208),
.B(n_2202),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2224),
.B(n_2210),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2221),
.B(n_2214),
.Y(n_2236)
);

AOI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2218),
.A2(n_2136),
.B1(n_2148),
.B2(n_2161),
.C(n_2159),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2226),
.B(n_2122),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2219),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2219),
.Y(n_2240)
);

OAI21xp33_ASAP7_75t_L g2241 ( 
.A1(n_2228),
.A2(n_2190),
.B(n_2155),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2223),
.Y(n_2242)
);

NOR2x1_ASAP7_75t_L g2243 ( 
.A(n_2225),
.B(n_2190),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2229),
.B(n_2154),
.Y(n_2244)
);

AOI221xp5_ASAP7_75t_L g2245 ( 
.A1(n_2233),
.A2(n_2230),
.B1(n_2227),
.B2(n_2232),
.C(n_2220),
.Y(n_2245)
);

NOR2x1_ASAP7_75t_L g2246 ( 
.A(n_2239),
.B(n_2227),
.Y(n_2246)
);

NOR4xp25_ASAP7_75t_L g2247 ( 
.A(n_2240),
.B(n_2232),
.C(n_2231),
.D(n_2129),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2234),
.A2(n_2220),
.B(n_2136),
.Y(n_2248)
);

AOI221xp5_ASAP7_75t_L g2249 ( 
.A1(n_2241),
.A2(n_2237),
.B1(n_2236),
.B2(n_2242),
.C(n_2235),
.Y(n_2249)
);

NAND5xp2_ASAP7_75t_L g2250 ( 
.A(n_2238),
.B(n_2165),
.C(n_2154),
.D(n_2155),
.E(n_2122),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2243),
.B(n_2038),
.Y(n_2251)
);

INVxp67_ASAP7_75t_L g2252 ( 
.A(n_2244),
.Y(n_2252)
);

NAND3xp33_ASAP7_75t_L g2253 ( 
.A(n_2244),
.B(n_2150),
.C(n_2132),
.Y(n_2253)
);

OAI221xp5_ASAP7_75t_L g2254 ( 
.A1(n_2245),
.A2(n_2158),
.B1(n_2152),
.B2(n_2150),
.C(n_2132),
.Y(n_2254)
);

OAI21x1_ASAP7_75t_SL g2255 ( 
.A1(n_2248),
.A2(n_2150),
.B(n_2132),
.Y(n_2255)
);

AOI221x1_ASAP7_75t_L g2256 ( 
.A1(n_2253),
.A2(n_2158),
.B1(n_2152),
.B2(n_2101),
.C(n_2099),
.Y(n_2256)
);

NAND3xp33_ASAP7_75t_SL g2257 ( 
.A(n_2249),
.B(n_2158),
.C(n_2152),
.Y(n_2257)
);

NAND5xp2_ASAP7_75t_L g2258 ( 
.A(n_2251),
.B(n_2123),
.C(n_2038),
.D(n_2032),
.E(n_2049),
.Y(n_2258)
);

OAI311xp33_ASAP7_75t_L g2259 ( 
.A1(n_2252),
.A2(n_2084),
.A3(n_2102),
.B1(n_2123),
.C1(n_2038),
.Y(n_2259)
);

OAI211xp5_ASAP7_75t_L g2260 ( 
.A1(n_2246),
.A2(n_2101),
.B(n_2124),
.C(n_2099),
.Y(n_2260)
);

OAI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2247),
.A2(n_1988),
.B1(n_2124),
.B2(n_2101),
.Y(n_2261)
);

NOR3xp33_ASAP7_75t_L g2262 ( 
.A(n_2250),
.B(n_2124),
.C(n_2115),
.Y(n_2262)
);

XNOR2x1_ASAP7_75t_L g2263 ( 
.A(n_2261),
.B(n_2084),
.Y(n_2263)
);

HB1xp67_ASAP7_75t_L g2264 ( 
.A(n_2254),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2262),
.B(n_2036),
.Y(n_2265)
);

OAI322xp33_ASAP7_75t_L g2266 ( 
.A1(n_2259),
.A2(n_2125),
.A3(n_2115),
.B1(n_2041),
.B2(n_2043),
.C1(n_2102),
.C2(n_2011),
.Y(n_2266)
);

NOR2x1_ASAP7_75t_L g2267 ( 
.A(n_2257),
.B(n_2260),
.Y(n_2267)
);

AO22x2_ASAP7_75t_L g2268 ( 
.A1(n_2255),
.A2(n_2125),
.B1(n_2041),
.B2(n_2056),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2258),
.B(n_2043),
.Y(n_2269)
);

OAI211xp5_ASAP7_75t_L g2270 ( 
.A1(n_2264),
.A2(n_2267),
.B(n_2269),
.C(n_2265),
.Y(n_2270)
);

OR3x2_ASAP7_75t_L g2271 ( 
.A(n_2263),
.B(n_2256),
.C(n_2028),
.Y(n_2271)
);

OR3x2_ASAP7_75t_L g2272 ( 
.A(n_2266),
.B(n_2040),
.C(n_2060),
.Y(n_2272)
);

AND4x1_ASAP7_75t_L g2273 ( 
.A(n_2268),
.B(n_2049),
.C(n_2056),
.D(n_2021),
.Y(n_2273)
);

OAI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2268),
.A2(n_2041),
.B(n_2049),
.Y(n_2274)
);

XOR2xp5_ASAP7_75t_L g2275 ( 
.A(n_2271),
.B(n_1832),
.Y(n_2275)
);

NAND5xp2_ASAP7_75t_L g2276 ( 
.A(n_2270),
.B(n_2274),
.C(n_2272),
.D(n_2273),
.E(n_2056),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2275),
.A2(n_2041),
.B1(n_2011),
.B2(n_1988),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2276),
.A2(n_1974),
.B1(n_2036),
.B2(n_2061),
.Y(n_2278)
);

XNOR2xp5_ASAP7_75t_L g2279 ( 
.A(n_2277),
.B(n_1974),
.Y(n_2279)
);

AOI211xp5_ASAP7_75t_L g2280 ( 
.A1(n_2278),
.A2(n_1974),
.B(n_2040),
.C(n_2060),
.Y(n_2280)
);

AOI22x1_ASAP7_75t_L g2281 ( 
.A1(n_2279),
.A2(n_1859),
.B1(n_2073),
.B2(n_2070),
.Y(n_2281)
);

XNOR2xp5_ASAP7_75t_L g2282 ( 
.A(n_2280),
.B(n_1974),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2282),
.B(n_2047),
.Y(n_2283)
);

AOI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2281),
.A2(n_2061),
.B1(n_2036),
.B2(n_1981),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2283),
.A2(n_2064),
.B(n_2047),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_2285),
.A2(n_2284),
.B(n_2064),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2286),
.Y(n_2287)
);

OAI221xp5_ASAP7_75t_R g2288 ( 
.A1(n_2287),
.A2(n_1938),
.B1(n_1835),
.B2(n_2065),
.C(n_1858),
.Y(n_2288)
);

AOI211xp5_ASAP7_75t_L g2289 ( 
.A1(n_2288),
.A2(n_2059),
.B(n_2057),
.C(n_2062),
.Y(n_2289)
);


endmodule