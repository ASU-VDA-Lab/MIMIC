module fake_jpeg_12253_n_41 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_41);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_17;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_7),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_1),
.B1(n_3),
.B2(n_12),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_1),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_16),
.A2(n_15),
.B(n_24),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_31),
.B1(n_28),
.B2(n_23),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_18),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_34),
.B1(n_35),
.B2(n_22),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_38),
.B(n_21),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_30),
.B(n_16),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AOI31xp33_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_25),
.A3(n_17),
.B(n_19),
.Y(n_41)
);


endmodule