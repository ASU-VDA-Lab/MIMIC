module fake_jpeg_17724_n_33 (n_3, n_2, n_1, n_0, n_4, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx5_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_10),
.B(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_12),
.Y(n_17)
);

AND2x2_ASAP7_75t_SL g12 ( 
.A(n_7),
.B(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_4),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_16),
.B1(n_14),
.B2(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

BUFx12f_ASAP7_75t_SL g21 ( 
.A(n_19),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_21),
.B(n_22),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_2),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

OAI21x1_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_21),
.B(n_23),
.Y(n_28)
);

OAI211xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_22),
.B(n_26),
.C(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_18),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_4),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_20),
.B2(n_5),
.Y(n_32)
);

AOI31xp33_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_5),
.A3(n_8),
.B(n_3),
.Y(n_33)
);


endmodule