module real_jpeg_14557_n_6 (n_46, n_5, n_4, n_43, n_0, n_1, n_2, n_45, n_42, n_44, n_3, n_6);

input n_46;
input n_5;
input n_4;
input n_43;
input n_0;
input n_1;
input n_2;
input n_45;
input n_42;
input n_44;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_33;
wire n_38;
wire n_35;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_39;
wire n_40;
wire n_36;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_1),
.B(n_11),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_11),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_2),
.B(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_4),
.B(n_34),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g6 ( 
.A(n_7),
.Y(n_6)
);

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_15),
.B1(n_39),
.B2(n_40),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_9),
.B(n_14),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_13),
.Y(n_11)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_33),
.B(n_38),
.Y(n_15)
);

OA21x2_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_21),
.B(n_32),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_31),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_42),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_43),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_44),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_45),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_46),
.Y(n_35)
);


endmodule