module fake_jpeg_1220_n_81 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_81);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_81;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx5_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_19),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_27),
.A2(n_28),
.B1(n_19),
.B2(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_10),
.B1(n_16),
.B2(n_20),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_22),
.B1(n_17),
.B2(n_15),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_19),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_17),
.C(n_20),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_34),
.C(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_8),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_33),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_49),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_15),
.B1(n_36),
.B2(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVxp33_ASAP7_75t_SL g65 ( 
.A(n_55),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_44),
.B1(n_51),
.B2(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_63),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_60),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_52),
.B(n_47),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_56),
.C(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_60),
.B1(n_59),
.B2(n_65),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_58),
.C(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_65),
.Y(n_77)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_78),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_79),
.A2(n_57),
.B(n_55),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_57),
.B(n_32),
.Y(n_81)
);


endmodule