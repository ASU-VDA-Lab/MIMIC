module fake_jpeg_5168_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_5),
.B(n_1),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx11_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_14),
.Y(n_16)
);

OR2x2_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_0),
.Y(n_13)
);

AOI21xp5_ASAP7_75t_L g15 ( 
.A1(n_13),
.A2(n_6),
.B(n_11),
.Y(n_15)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_12),
.B(n_13),
.C(n_7),
.Y(n_22)
);

NOR4xp25_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_13),
.C(n_12),
.D(n_6),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_23),
.A2(n_22),
.B(n_7),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_19),
.C(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_10),
.Y(n_25)
);

OAI322xp33_ASAP7_75t_L g29 ( 
.A1(n_27),
.A2(n_10),
.A3(n_11),
.B1(n_7),
.B2(n_8),
.C1(n_5),
.C2(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_27),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_26),
.B1(n_8),
.B2(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

XOR2x2_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_33),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_4),
.C(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_0),
.Y(n_38)
);


endmodule