module real_jpeg_24330_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_79),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_1),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_79),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_25),
.B1(n_29),
.B2(n_79),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_2),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_58),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_25),
.B1(n_29),
.B2(n_58),
.Y(n_162)
);

INVx8_ASAP7_75t_SL g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_6),
.A2(n_25),
.B1(n_29),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_70),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_10),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_10),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_10),
.B(n_53),
.C(n_54),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_10),
.B(n_77),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_52),
.B1(n_53),
.B2(n_98),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_10),
.B(n_25),
.C(n_85),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_10),
.A2(n_24),
.B(n_150),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_12),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_61),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_40),
.B1(n_45),
.B2(n_61),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_61),
.Y(n_122)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_14),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_125),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_102),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_18),
.B(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_72),
.B2(n_73),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_49),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_35),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_23),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_160)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_24),
.A2(n_28),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_24),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_25),
.A2(n_29),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_29),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_31),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.A3(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_37),
.B1(n_54),
.B2(n_55),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_37),
.B1(n_42),
.B2(n_48),
.Y(n_67)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_37),
.B(n_115),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_40),
.A2(n_41),
.B1(n_42),
.B2(n_48),
.Y(n_92)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_44),
.Y(n_99)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_65),
.C(n_68),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_56),
.B(n_59),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_53),
.B1(n_84),
.B2(n_85),
.Y(n_88)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_53),
.B(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_62),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_60),
.B(n_77),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_63),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_90),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_86),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_83),
.A2(n_86),
.B(n_131),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_83),
.B(n_98),
.Y(n_169)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_87),
.A2(n_110),
.B1(n_112),
.B2(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B(n_100),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_101),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B(n_99),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_98),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_113),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_104),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_113),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B(n_111),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_108),
.A2(n_111),
.B(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_116),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_120),
.A2(n_162),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_139),
.B(n_187),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_136),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.C(n_132),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_128),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_129),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_181),
.B(n_186),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_158),
.B(n_180),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_152),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_152),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_147),
.C(n_148),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_149),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_167),
.B(n_179),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_165),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_165),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_172),
.B(n_178),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_185),
.Y(n_186)
);


endmodule