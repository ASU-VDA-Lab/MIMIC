module fake_jpeg_15521_n_39 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_39);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_39;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

INVx2_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx4f_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_SL g19 ( 
.A1(n_16),
.A2(n_12),
.B(n_10),
.C(n_9),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_22),
.B1(n_17),
.B2(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_21),
.B(n_17),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_14),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_18),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_18),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_25),
.B(n_19),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_21),
.B1(n_22),
.B2(n_4),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_15),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_20),
.C(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.C(n_0),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_3),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_32),
.C2(n_33),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_5),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_37),
.C(n_34),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_6),
.Y(n_39)
);


endmodule