module fake_ariane_1225_n_911 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_32, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_911);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_32;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_911;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_64;
wire n_180;
wire n_730;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_34;
wire n_172;
wire n_678;
wire n_651;
wire n_423;
wire n_347;
wire n_469;
wire n_183;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_133;
wire n_610;
wire n_66;
wire n_205;
wire n_752;
wire n_341;
wire n_71;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_549;
wire n_522;
wire n_319;
wire n_49;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_50;
wire n_187;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_103;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_36;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_72;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_57;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_117;
wire n_139;
wire n_524;
wire n_85;
wire n_130;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_138;
wire n_162;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_137;
wire n_885;
wire n_122;
wire n_198;
wire n_232;
wire n_52;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_73;
wire n_327;
wire n_77;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_87;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_41;
wire n_813;
wire n_140;
wire n_725;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_154;
wire n_883;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_145;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_59;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_35;
wire n_54;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_167;
wire n_90;
wire n_38;
wire n_422;
wire n_47;
wire n_153;
wire n_784;
wire n_648;
wire n_269;
wire n_597;
wire n_816;
wire n_75;
wire n_855;
wire n_158;
wire n_69;
wire n_259;
wire n_835;
wire n_95;
wire n_808;
wire n_446;
wire n_553;
wire n_143;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_152;
wire n_557;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_115;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_62;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_561;
wire n_770;
wire n_253;
wire n_218;
wire n_821;
wire n_79;
wire n_839;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_91;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_44;
wire n_82;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_48;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_108;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_81;
wire n_352;
wire n_538;
wire n_206;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_136;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_163;
wire n_88;
wire n_869;
wire n_141;
wire n_846;
wire n_390;
wire n_498;
wire n_104;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_56;
wire n_60;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_86;
wire n_361;
wire n_458;
wire n_89;
wire n_149;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_175;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_74;
wire n_491;
wire n_810;
wire n_40;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_658;
wire n_630;
wire n_570;
wire n_53;
wire n_362;
wire n_260;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_46;
wire n_741;
wire n_747;
wire n_772;
wire n_84;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_107;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_42;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_70;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_94;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_534;
wire n_249;
wire n_355;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_444;
wire n_212;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_135;
wire n_896;
wire n_409;
wire n_171;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_61;
wire n_526;
wire n_716;
wire n_102;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_798;
wire n_769;
wire n_820;
wire n_43;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_55;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_252;
wire n_664;
wire n_629;
wire n_215;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_68;
wire n_415;
wire n_794;
wire n_763;
wire n_78;
wire n_63;
wire n_655;
wire n_99;
wire n_544;
wire n_540;
wire n_692;
wire n_216;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_83;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_110;
wire n_304;
wire n_895;
wire n_659;
wire n_67;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_92;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_757;
wire n_375;
wire n_113;
wire n_114;
wire n_33;
wire n_324;
wire n_585;
wire n_875;
wire n_785;
wire n_669;
wire n_827;
wire n_619;
wire n_437;
wire n_337;
wire n_111;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_174;
wire n_275;
wire n_100;
wire n_704;
wire n_132;
wire n_147;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_51;
wire n_496;
wire n_739;
wire n_76;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_131;
wire n_434;
wire n_263;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_144;
wire n_882;
wire n_317;
wire n_867;
wire n_101;
wire n_243;
wire n_803;
wire n_134;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_112;
wire n_45;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_470;
wire n_266;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_121;
wire n_118;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_382;
wire n_191;
wire n_797;
wire n_489;
wire n_80;
wire n_480;
wire n_211;
wire n_642;
wire n_97;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_116;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_39;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_796;
wire n_805;
wire n_127;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_11),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_1),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_1),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_2),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_3),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_5),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_27),
.Y(n_80)
);

OR2x6_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_47),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_39),
.B1(n_63),
.B2(n_62),
.Y(n_82)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_39),
.B1(n_63),
.B2(n_62),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_80),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_77),
.B1(n_35),
.B2(n_80),
.Y(n_85)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_41),
.B1(n_64),
.B2(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_73),
.A2(n_41),
.B1(n_64),
.B2(n_42),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_65),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_40),
.B1(n_42),
.B2(n_55),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_60),
.B1(n_58),
.B2(n_55),
.Y(n_95)
);

CKINVDCx6p67_ASAP7_75t_R g96 ( 
.A(n_69),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_60),
.Y(n_97)
);

OR2x6_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_58),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_54),
.B1(n_53),
.B2(n_51),
.Y(n_99)
);

AND2x4_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_33),
.B1(n_59),
.B2(n_56),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

AO22x2_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_51),
.B1(n_54),
.B2(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_69),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_74),
.B(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_69),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_100),
.B(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_66),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_66),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_69),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_66),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_67),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_77),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_70),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_86),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_77),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_90),
.A2(n_74),
.B(n_78),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_L g136 ( 
.A(n_87),
.B(n_70),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_67),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_70),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_67),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_82),
.B(n_37),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_95),
.A2(n_78),
.B(n_74),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_67),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_70),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_70),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_81),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_81),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_109),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_124),
.B(n_81),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_97),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_93),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g167 ( 
.A(n_142),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_143),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_83),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_75),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_75),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_115),
.B(n_78),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_144),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_149),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_83),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_78),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_68),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_146),
.B(n_78),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_123),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_83),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_78),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_113),
.B(n_68),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_133),
.B(n_75),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_136),
.B(n_83),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_128),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_128),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_135),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_148),
.B(n_99),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_108),
.B(n_75),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_99),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_106),
.B(n_75),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_151),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_99),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_111),
.B(n_78),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_70),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_141),
.B(n_70),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_130),
.B(n_75),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_145),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_155),
.B(n_164),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_147),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_167),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_147),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_131),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_155),
.B(n_134),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_218),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

BUFx8_ASAP7_75t_SL g236 ( 
.A(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_162),
.B(n_137),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_162),
.B(n_68),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_170),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_187),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_162),
.B(n_137),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g246 ( 
.A(n_155),
.B(n_134),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_118),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_162),
.B(n_141),
.Y(n_248)
);

NAND2x1p5_ASAP7_75t_L g249 ( 
.A(n_218),
.B(n_76),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_155),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_L g252 ( 
.A(n_169),
.B(n_75),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_209),
.B(n_141),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_155),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

AND2x4_ASAP7_75t_L g257 ( 
.A(n_155),
.B(n_68),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_187),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_118),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_193),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_193),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_170),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_181),
.B(n_114),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_193),
.Y(n_266)
);

AND2x4_ASAP7_75t_L g267 ( 
.A(n_155),
.B(n_76),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_209),
.B(n_179),
.Y(n_268)
);

OR2x6_ASAP7_75t_L g269 ( 
.A(n_155),
.B(n_72),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_165),
.B(n_114),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_170),
.Y(n_271)
);

AND2x4_ASAP7_75t_L g272 ( 
.A(n_164),
.B(n_72),
.Y(n_272)
);

AND2x4_ASAP7_75t_L g273 ( 
.A(n_164),
.B(n_72),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_190),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

NAND2x1p5_ASAP7_75t_L g277 ( 
.A(n_218),
.B(n_72),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_192),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

OR2x6_ASAP7_75t_L g280 ( 
.A(n_156),
.B(n_72),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_192),
.Y(n_281)
);

BUFx4f_ASAP7_75t_L g282 ( 
.A(n_172),
.Y(n_282)
);

OR2x6_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_156),
.Y(n_283)
);

NAND2x1p5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_244),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_231),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_236),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_192),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_192),
.Y(n_289)
);

INVx6_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g291 ( 
.A(n_275),
.Y(n_291)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_236),
.Y(n_293)
);

BUFx4f_ASAP7_75t_SL g294 ( 
.A(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_239),
.B(n_166),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

OR2x6_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_156),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_238),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_238),
.Y(n_300)
);

BUFx8_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_238),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_268),
.B(n_166),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_221),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_281),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_229),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

BUFx12f_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_282),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_278),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_238),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_221),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_226),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_239),
.A2(n_209),
.B1(n_165),
.B2(n_195),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_195),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_228),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_221),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g319 ( 
.A(n_222),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_281),
.Y(n_320)
);

BUFx12f_ASAP7_75t_L g321 ( 
.A(n_229),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_269),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_282),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_224),
.A2(n_195),
.B1(n_211),
.B2(n_194),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_223),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_222),
.B(n_164),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_282),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_226),
.B(n_166),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_238),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_227),
.B(n_166),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_275),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_227),
.B(n_165),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_238),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_240),
.Y(n_338)
);

INVx5_ASAP7_75t_SL g339 ( 
.A(n_269),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_233),
.Y(n_340)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_269),
.Y(n_341)
);

NAND2x1p5_ASAP7_75t_L g342 ( 
.A(n_244),
.B(n_218),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_223),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_238),
.Y(n_344)
);

BUFx2_ASAP7_75t_SL g345 ( 
.A(n_274),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_233),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_274),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_224),
.B(n_184),
.Y(n_348)
);

BUFx4f_ASAP7_75t_L g349 ( 
.A(n_222),
.Y(n_349)
);

CKINVDCx6p67_ASAP7_75t_R g350 ( 
.A(n_223),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_239),
.B(n_164),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_265),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_239),
.B(n_184),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_300),
.A2(n_264),
.B(n_274),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_306),
.A2(n_247),
.B1(n_259),
.B2(n_265),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_297),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_316),
.B(n_247),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_315),
.A2(n_178),
.B1(n_209),
.B2(n_264),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_325),
.A2(n_247),
.B1(n_259),
.B2(n_195),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_306),
.A2(n_259),
.B1(n_270),
.B2(n_207),
.Y(n_361)
);

BUFx6f_ASAP7_75t_SL g362 ( 
.A(n_285),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_348),
.A2(n_270),
.B1(n_245),
.B2(n_160),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_316),
.A2(n_160),
.B1(n_163),
.B2(n_184),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g366 ( 
.A1(n_308),
.A2(n_211),
.B1(n_207),
.B2(n_198),
.Y(n_366)
);

INVx4_ASAP7_75t_SL g367 ( 
.A(n_291),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_312),
.B(n_274),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_289),
.A2(n_178),
.B1(n_264),
.B2(n_241),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_285),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_353),
.A2(n_160),
.B1(n_163),
.B2(n_184),
.Y(n_372)
);

BUFx2_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_314),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_305),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_L g377 ( 
.A1(n_303),
.A2(n_163),
.B1(n_269),
.B2(n_254),
.Y(n_377)
);

INVx8_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

INVx4_ASAP7_75t_SL g379 ( 
.A(n_291),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_308),
.A2(n_211),
.B1(n_198),
.B2(n_188),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

CKINVDCx11_ASAP7_75t_R g382 ( 
.A(n_287),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_329),
.A2(n_178),
.B1(n_241),
.B2(n_271),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_346),
.Y(n_384)
);

INVx4_ASAP7_75t_SL g385 ( 
.A(n_292),
.Y(n_385)
);

BUFx12f_ASAP7_75t_L g386 ( 
.A(n_321),
.Y(n_386)
);

CKINVDCx6p67_ASAP7_75t_R g387 ( 
.A(n_293),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_321),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_332),
.A2(n_178),
.B1(n_256),
.B2(n_271),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_352),
.A2(n_211),
.B1(n_198),
.B2(n_171),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_330),
.A2(n_198),
.B1(n_182),
.B2(n_188),
.Y(n_392)
);

CKINVDCx8_ASAP7_75t_R g393 ( 
.A(n_312),
.Y(n_393)
);

INVx6_ASAP7_75t_SL g394 ( 
.A(n_327),
.Y(n_394)
);

BUFx12f_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

CKINVDCx11_ASAP7_75t_R g396 ( 
.A(n_320),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_288),
.B(n_189),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_288),
.B(n_171),
.Y(n_398)
);

INVx8_ASAP7_75t_L g399 ( 
.A(n_286),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_295),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_335),
.A2(n_178),
.B1(n_256),
.B2(n_254),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_292),
.A2(n_245),
.B1(n_274),
.B2(n_257),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_294),
.Y(n_405)
);

CKINVDCx11_ASAP7_75t_R g406 ( 
.A(n_350),
.Y(n_406)
);

INVx8_ASAP7_75t_L g407 ( 
.A(n_286),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_349),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_304),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_296),
.A2(n_204),
.B(n_237),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_351),
.A2(n_274),
.B1(n_257),
.B2(n_234),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_295),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_334),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_283),
.A2(n_189),
.B1(n_194),
.B2(n_46),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_296),
.B(n_171),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_L g416 ( 
.A1(n_351),
.A2(n_182),
.B1(n_188),
.B2(n_171),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_334),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_290),
.A2(n_274),
.B1(n_257),
.B2(n_235),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_375),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_361),
.A2(n_213),
.B1(n_182),
.B2(n_188),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_357),
.B(n_319),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_359),
.A2(n_257),
.B(n_213),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_414),
.A2(n_182),
.B1(n_203),
.B2(n_205),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_257),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_361),
.A2(n_355),
.B1(n_360),
.B2(n_366),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_412),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_400),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_355),
.A2(n_222),
.B1(n_327),
.B2(n_203),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_364),
.A2(n_349),
.B1(n_312),
.B2(n_323),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_370),
.A2(n_349),
.B1(n_312),
.B2(n_323),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_SL g433 ( 
.A1(n_402),
.A2(n_205),
.B1(n_203),
.B2(n_339),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_360),
.A2(n_222),
.B1(n_327),
.B2(n_205),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_368),
.A2(n_373),
.B1(n_388),
.B2(n_371),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_383),
.A2(n_341),
.B1(n_323),
.B2(n_290),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_319),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_366),
.A2(n_203),
.B1(n_205),
.B2(n_248),
.Y(n_442)
);

BUFx4f_ASAP7_75t_SL g443 ( 
.A(n_386),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_365),
.A2(n_283),
.B1(n_298),
.B2(n_248),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_356),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_391),
.A2(n_380),
.B1(n_392),
.B2(n_372),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_338),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_389),
.A2(n_323),
.B1(n_341),
.B2(n_290),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_377),
.A2(n_322),
.B(n_333),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_377),
.A2(n_365),
.B1(n_372),
.B2(n_341),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_338),
.Y(n_451)
);

BUFx2_ASAP7_75t_SL g452 ( 
.A(n_375),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_404),
.A2(n_323),
.B1(n_341),
.B2(n_290),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_391),
.A2(n_298),
.B1(n_283),
.B2(n_255),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_363),
.Y(n_455)
);

BUFx6f_ASAP7_75t_SL g456 ( 
.A(n_358),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_368),
.A2(n_339),
.B1(n_341),
.B2(n_251),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_368),
.A2(n_339),
.B1(n_251),
.B2(n_225),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_304),
.Y(n_459)
);

OR2x2_ASAP7_75t_L g460 ( 
.A(n_411),
.B(n_410),
.Y(n_460)
);

INVx5_ASAP7_75t_SL g461 ( 
.A(n_387),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_413),
.Y(n_463)
);

CKINVDCx6p67_ASAP7_75t_R g464 ( 
.A(n_406),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_380),
.A2(n_298),
.B1(n_283),
.B2(n_255),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_375),
.B(n_313),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_392),
.A2(n_298),
.B1(n_251),
.B2(n_255),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_416),
.B(n_267),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_395),
.A2(n_225),
.B1(n_237),
.B2(n_280),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_267),
.Y(n_470)
);

OAI22xp33_ASAP7_75t_L g471 ( 
.A1(n_408),
.A2(n_280),
.B1(n_269),
.B2(n_286),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_426),
.A2(n_232),
.B1(n_230),
.B2(n_225),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_423),
.A2(n_230),
.B1(n_232),
.B2(n_417),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_421),
.B(n_343),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_450),
.A2(n_375),
.B1(n_339),
.B2(n_362),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_446),
.A2(n_230),
.B1(n_232),
.B2(n_280),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_460),
.A2(n_362),
.B1(n_418),
.B2(n_318),
.Y(n_477)
);

OAI222xp33_ASAP7_75t_L g478 ( 
.A1(n_420),
.A2(n_393),
.B1(n_280),
.B2(n_34),
.C1(n_61),
.C2(n_44),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_433),
.A2(n_232),
.B1(n_230),
.B2(n_280),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_422),
.A2(n_405),
.B(n_322),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_468),
.A2(n_232),
.B1(n_230),
.B2(n_280),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_468),
.A2(n_280),
.B1(n_326),
.B2(n_313),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_460),
.A2(n_333),
.B1(n_328),
.B2(n_324),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_470),
.A2(n_326),
.B1(n_318),
.B2(n_208),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_470),
.A2(n_208),
.B1(n_244),
.B2(n_394),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_444),
.A2(n_324),
.B1(n_309),
.B2(n_328),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_442),
.A2(n_454),
.B1(n_465),
.B2(n_430),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_467),
.A2(n_208),
.B1(n_244),
.B2(n_394),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_309),
.B1(n_322),
.B2(n_284),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_451),
.A2(n_208),
.B1(n_244),
.B2(n_267),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_469),
.A2(n_284),
.B1(n_350),
.B2(n_274),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_435),
.A2(n_269),
.B1(n_267),
.B2(n_45),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_431),
.A2(n_267),
.B1(n_49),
.B2(n_52),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_425),
.Y(n_495)
);

AOI22xp33_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_208),
.B1(n_196),
.B2(n_217),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_438),
.B(n_369),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_439),
.A2(n_196),
.B1(n_217),
.B2(n_343),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_432),
.A2(n_448),
.B1(n_453),
.B2(n_452),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_440),
.A2(n_284),
.B1(n_234),
.B2(n_235),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_440),
.A2(n_234),
.B1(n_235),
.B2(n_246),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_471),
.A2(n_196),
.B1(n_217),
.B2(n_242),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_462),
.A2(n_242),
.B1(n_210),
.B2(n_246),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_462),
.A2(n_242),
.B1(n_210),
.B2(n_246),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_463),
.A2(n_424),
.B1(n_429),
.B2(n_445),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_463),
.A2(n_210),
.B1(n_246),
.B2(n_200),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_421),
.B(n_311),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_452),
.A2(n_190),
.B1(n_345),
.B2(n_48),
.Y(n_508)
);

AOI221xp5_ASAP7_75t_SL g509 ( 
.A1(n_437),
.A2(n_427),
.B1(n_455),
.B2(n_438),
.C(n_441),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_437),
.B(n_427),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_436),
.A2(n_179),
.B1(n_164),
.B2(n_190),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_456),
.A2(n_190),
.B1(n_345),
.B2(n_378),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_429),
.A2(n_210),
.B1(n_246),
.B2(n_200),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_461),
.A2(n_235),
.B1(n_234),
.B2(n_246),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_461),
.A2(n_235),
.B1(n_234),
.B2(n_246),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_434),
.A2(n_179),
.B1(n_164),
.B2(n_190),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_456),
.A2(n_190),
.B1(n_185),
.B2(n_161),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_447),
.B(n_240),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_441),
.A2(n_447),
.B1(n_428),
.B2(n_458),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_428),
.A2(n_210),
.B1(n_200),
.B2(n_240),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_456),
.A2(n_190),
.B1(n_399),
.B2(n_378),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_72),
.C(n_354),
.Y(n_522)
);

NAND4xp25_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_459),
.C(n_354),
.D(n_173),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_511),
.A2(n_461),
.B1(n_464),
.B2(n_457),
.Y(n_524)
);

AOI221xp5_ASAP7_75t_L g525 ( 
.A1(n_509),
.A2(n_72),
.B1(n_75),
.B2(n_273),
.C(n_272),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_461),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_L g527 ( 
.A(n_480),
.B(n_382),
.C(n_72),
.Y(n_527)
);

NAND3xp33_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_72),
.C(n_419),
.Y(n_528)
);

OA21x2_ASAP7_75t_L g529 ( 
.A1(n_480),
.A2(n_419),
.B(n_466),
.Y(n_529)
);

AOI221xp5_ASAP7_75t_L g530 ( 
.A1(n_478),
.A2(n_75),
.B1(n_273),
.B2(n_272),
.C(n_185),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g531 ( 
.A(n_522),
.B(n_154),
.C(n_161),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_495),
.B(n_466),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_511),
.A2(n_464),
.B1(n_443),
.B2(n_302),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_497),
.B(n_466),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_482),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_5),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_344),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_505),
.B(n_6),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_474),
.B(n_518),
.Y(n_539)
);

OAI221xp5_ASAP7_75t_L g540 ( 
.A1(n_488),
.A2(n_185),
.B1(n_173),
.B2(n_161),
.C(n_154),
.Y(n_540)
);

AND4x1_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_367),
.C(n_379),
.D(n_385),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_344),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_493),
.A2(n_154),
.B1(n_173),
.B2(n_385),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_477),
.B(n_153),
.C(n_174),
.Y(n_544)
);

OA21x2_ASAP7_75t_L g545 ( 
.A1(n_519),
.A2(n_153),
.B(n_157),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_517),
.A2(n_299),
.B1(n_347),
.B2(n_336),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_500),
.B(n_344),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_494),
.A2(n_190),
.B(n_214),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_496),
.B(n_6),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_485),
.B(n_7),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_499),
.B(n_299),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_514),
.A2(n_234),
.B(n_235),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_L g553 ( 
.A(n_494),
.B(n_157),
.C(n_177),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_475),
.B(n_367),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_512),
.B(n_367),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_517),
.B(n_379),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_473),
.A2(n_243),
.B1(n_262),
.B2(n_263),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_484),
.B(n_9),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_10),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_502),
.B(n_378),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g561 ( 
.A(n_486),
.B(n_180),
.C(n_177),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_516),
.B(n_159),
.C(n_158),
.Y(n_562)
);

OAI221xp5_ASAP7_75t_SL g563 ( 
.A1(n_493),
.A2(n_204),
.B1(n_197),
.B2(n_176),
.C(n_18),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g564 ( 
.A(n_483),
.B(n_180),
.C(n_177),
.Y(n_564)
);

OAI221xp5_ASAP7_75t_SL g565 ( 
.A1(n_516),
.A2(n_204),
.B1(n_197),
.B2(n_176),
.C(n_18),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_487),
.B(n_157),
.C(n_180),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_490),
.B(n_299),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_492),
.B(n_10),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_520),
.B(n_159),
.C(n_180),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_515),
.B(n_299),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_491),
.B(n_13),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_535),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_539),
.B(n_503),
.Y(n_573)
);

AO21x2_ASAP7_75t_L g574 ( 
.A1(n_568),
.A2(n_214),
.B(n_279),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_524),
.A2(n_479),
.B1(n_472),
.B2(n_476),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_537),
.B(n_504),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_532),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_523),
.B(n_521),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_532),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_534),
.B(n_481),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_536),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_529),
.B(n_299),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_537),
.B(n_506),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_529),
.B(n_302),
.Y(n_584)
);

NAND3xp33_ASAP7_75t_L g585 ( 
.A(n_528),
.B(n_508),
.C(n_489),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_529),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_529),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_526),
.B(n_545),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_545),
.A2(n_513),
.B1(n_243),
.B2(n_250),
.Y(n_589)
);

OR2x6_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_399),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_545),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_567),
.B(n_302),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_545),
.B(n_13),
.Y(n_593)
);

AOI211xp5_ASAP7_75t_L g594 ( 
.A1(n_563),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_594)
);

AOI221xp5_ASAP7_75t_L g595 ( 
.A1(n_538),
.A2(n_273),
.B1(n_272),
.B2(n_22),
.C(n_23),
.Y(n_595)
);

AOI221xp5_ASAP7_75t_L g596 ( 
.A1(n_550),
.A2(n_272),
.B1(n_273),
.B2(n_24),
.C(n_26),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_542),
.B(n_547),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_528),
.B(n_302),
.C(n_347),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_551),
.B(n_302),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_527),
.A2(n_379),
.B1(n_385),
.B2(n_177),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_551),
.B(n_337),
.Y(n_601)
);

AOI221xp5_ASAP7_75t_L g602 ( 
.A1(n_565),
.A2(n_273),
.B1(n_272),
.B2(n_24),
.C(n_26),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_542),
.Y(n_603)
);

NOR3xp33_ASAP7_75t_L g604 ( 
.A(n_558),
.B(n_331),
.C(n_153),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_544),
.A2(n_174),
.B1(n_180),
.B2(n_177),
.Y(n_605)
);

NAND3xp33_ASAP7_75t_L g606 ( 
.A(n_553),
.B(n_336),
.C(n_347),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_547),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_564),
.A2(n_279),
.B1(n_261),
.B2(n_260),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_570),
.B(n_336),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_L g611 ( 
.A(n_559),
.B(n_331),
.C(n_174),
.Y(n_611)
);

NAND3xp33_ASAP7_75t_L g612 ( 
.A(n_553),
.B(n_336),
.C(n_347),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_552),
.B(n_336),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_543),
.A2(n_174),
.B1(n_159),
.B2(n_158),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_548),
.A2(n_276),
.B1(n_260),
.B2(n_258),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_533),
.B(n_337),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_546),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_566),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_541),
.B(n_16),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

OAI211xp5_ASAP7_75t_L g621 ( 
.A1(n_543),
.A2(n_19),
.B(n_27),
.C(n_407),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_562),
.Y(n_622)
);

AOI211xp5_ASAP7_75t_L g623 ( 
.A1(n_556),
.A2(n_212),
.B(n_157),
.C(n_152),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_531),
.B(n_337),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_571),
.B(n_337),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_549),
.B(n_337),
.C(n_347),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_597),
.B(n_560),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_594),
.A2(n_554),
.B1(n_555),
.B2(n_561),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_572),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_572),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_587),
.Y(n_631)
);

NAND4xp75_ASAP7_75t_SL g632 ( 
.A(n_619),
.B(n_541),
.C(n_540),
.D(n_212),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_587),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_610),
.Y(n_634)
);

NAND4xp75_ASAP7_75t_L g635 ( 
.A(n_578),
.B(n_525),
.C(n_530),
.D(n_557),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_610),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_620),
.B(n_569),
.C(n_331),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_607),
.Y(n_638)
);

BUFx2_ASAP7_75t_SL g639 ( 
.A(n_586),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_581),
.B(n_262),
.Y(n_640)
);

NAND4xp75_ASAP7_75t_L g641 ( 
.A(n_602),
.B(n_243),
.C(n_250),
.D(n_263),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_580),
.B(n_168),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_607),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_576),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_597),
.B(n_235),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_603),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_622),
.B(n_263),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_622),
.B(n_262),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_588),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_588),
.B(n_260),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_618),
.B(n_261),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_603),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_591),
.Y(n_654)
);

NAND4xp75_ASAP7_75t_L g655 ( 
.A(n_595),
.B(n_250),
.C(n_276),
.D(n_266),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_580),
.B(n_174),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_575),
.A2(n_621),
.B1(n_585),
.B2(n_596),
.Y(n_657)
);

NAND4xp75_ASAP7_75t_SL g658 ( 
.A(n_582),
.B(n_212),
.C(n_252),
.D(n_407),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_591),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_618),
.B(n_407),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_617),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_582),
.Y(n_662)
);

XOR2x2_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_342),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_590),
.B(n_584),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_590),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_577),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_590),
.B(n_234),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_584),
.B(n_342),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_617),
.B(n_261),
.Y(n_670)
);

XNOR2x2_ASAP7_75t_L g671 ( 
.A(n_593),
.B(n_279),
.Y(n_671)
);

INVx4_ASAP7_75t_L g672 ( 
.A(n_593),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_573),
.Y(n_673)
);

NAND4xp75_ASAP7_75t_SL g674 ( 
.A(n_613),
.B(n_212),
.C(n_252),
.D(n_399),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_574),
.Y(n_676)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_600),
.B(n_157),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_583),
.B(n_159),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_672),
.A2(n_626),
.B1(n_611),
.B2(n_604),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_657),
.B(n_661),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_627),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_627),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_631),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_631),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_665),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_638),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_665),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_638),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_642),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_643),
.Y(n_690)
);

XOR2x2_ASAP7_75t_L g691 ( 
.A(n_657),
.B(n_614),
.Y(n_691)
);

OA22x2_ASAP7_75t_L g692 ( 
.A1(n_642),
.A2(n_579),
.B1(n_625),
.B2(n_599),
.Y(n_692)
);

OA22x2_ASAP7_75t_L g693 ( 
.A1(n_628),
.A2(n_601),
.B1(n_605),
.B2(n_592),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_662),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_672),
.B(n_574),
.Y(n_696)
);

BUFx12f_ASAP7_75t_L g697 ( 
.A(n_672),
.Y(n_697)
);

XOR2x2_ASAP7_75t_L g698 ( 
.A(n_656),
.B(n_598),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_647),
.B(n_624),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_633),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_647),
.B(n_606),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_634),
.B(n_592),
.Y(n_702)
);

OA22x2_ASAP7_75t_L g703 ( 
.A1(n_628),
.A2(n_609),
.B1(n_616),
.B2(n_613),
.Y(n_703)
);

XNOR2xp5_ASAP7_75t_L g704 ( 
.A(n_656),
.B(n_609),
.Y(n_704)
);

XOR2xp5_ASAP7_75t_L g705 ( 
.A(n_663),
.B(n_616),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_643),
.Y(n_706)
);

XOR2x2_ASAP7_75t_L g707 ( 
.A(n_635),
.B(n_612),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_654),
.Y(n_708)
);

XNOR2xp5_ASAP7_75t_L g709 ( 
.A(n_632),
.B(n_615),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_666),
.Y(n_710)
);

HB1xp67_ASAP7_75t_L g711 ( 
.A(n_650),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_671),
.Y(n_712)
);

XNOR2x1_ASAP7_75t_L g713 ( 
.A(n_635),
.B(n_574),
.Y(n_713)
);

XNOR2x1_ASAP7_75t_L g714 ( 
.A(n_641),
.B(n_608),
.Y(n_714)
);

XNOR2x2_ASAP7_75t_L g715 ( 
.A(n_671),
.B(n_589),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_678),
.Y(n_716)
);

XOR2x2_ASAP7_75t_L g717 ( 
.A(n_641),
.B(n_342),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_666),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_640),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_636),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

XNOR2xp5_ASAP7_75t_L g723 ( 
.A(n_663),
.B(n_159),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_686),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_685),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_685),
.B(n_662),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_680),
.Y(n_727)
);

XNOR2x1_ASAP7_75t_L g728 ( 
.A(n_691),
.B(n_655),
.Y(n_728)
);

OA22x2_ASAP7_75t_L g729 ( 
.A1(n_689),
.A2(n_639),
.B1(n_673),
.B2(n_644),
.Y(n_729)
);

AOI22x1_ASAP7_75t_L g730 ( 
.A1(n_679),
.A2(n_639),
.B1(n_634),
.B2(n_636),
.Y(n_730)
);

XOR2x2_ASAP7_75t_L g731 ( 
.A(n_691),
.B(n_655),
.Y(n_731)
);

BUFx2_ASAP7_75t_L g732 ( 
.A(n_697),
.Y(n_732)
);

AO22x1_ASAP7_75t_L g733 ( 
.A1(n_680),
.A2(n_634),
.B1(n_662),
.B2(n_650),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_SL g734 ( 
.A1(n_693),
.A2(n_664),
.B1(n_677),
.B2(n_653),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_713),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_697),
.Y(n_736)
);

XOR2x2_ASAP7_75t_L g737 ( 
.A(n_707),
.B(n_674),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_688),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_687),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_713),
.Y(n_740)
);

OA22x2_ASAP7_75t_L g741 ( 
.A1(n_705),
.A2(n_664),
.B1(n_653),
.B2(n_675),
.Y(n_741)
);

OA22x2_ASAP7_75t_L g742 ( 
.A1(n_712),
.A2(n_646),
.B1(n_676),
.B2(n_677),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_690),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_707),
.Y(n_744)
);

OA22x2_ASAP7_75t_SL g745 ( 
.A1(n_703),
.A2(n_662),
.B1(n_646),
.B2(n_667),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_706),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_679),
.A2(n_637),
.B1(n_662),
.B2(n_660),
.Y(n_747)
);

INVxp33_ASAP7_75t_SL g748 ( 
.A(n_709),
.Y(n_748)
);

XNOR2x1_ASAP7_75t_L g749 ( 
.A(n_715),
.B(n_658),
.Y(n_749)
);

OAI22x1_ASAP7_75t_L g750 ( 
.A1(n_681),
.A2(n_662),
.B1(n_667),
.B2(n_630),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_719),
.Y(n_751)
);

AOI22x1_ASAP7_75t_L g752 ( 
.A1(n_679),
.A2(n_687),
.B1(n_694),
.B2(n_721),
.Y(n_752)
);

XNOR2x1_ASAP7_75t_L g753 ( 
.A(n_715),
.B(n_668),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_682),
.B(n_670),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_722),
.Y(n_755)
);

INVx4_ASAP7_75t_L g756 ( 
.A(n_687),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_693),
.A2(n_659),
.B1(n_654),
.B2(n_652),
.Y(n_757)
);

OA22x2_ASAP7_75t_L g758 ( 
.A1(n_704),
.A2(n_676),
.B1(n_659),
.B2(n_629),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_711),
.Y(n_759)
);

OA22x2_ASAP7_75t_L g760 ( 
.A1(n_716),
.A2(n_676),
.B1(n_629),
.B2(n_630),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_702),
.B(n_668),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_728),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_724),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_738),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_743),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_746),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_732),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_751),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_759),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_755),
.Y(n_770)
);

INVxp33_ASAP7_75t_L g771 ( 
.A(n_727),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_727),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_748),
.A2(n_714),
.B1(n_698),
.B2(n_703),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_731),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_739),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_752),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_754),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_754),
.Y(n_778)
);

OAI322xp33_ASAP7_75t_L g779 ( 
.A1(n_735),
.A2(n_696),
.A3(n_692),
.B1(n_701),
.B2(n_699),
.C1(n_714),
.C2(n_718),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_725),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_756),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_756),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_761),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_729),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_753),
.B(n_720),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_729),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_760),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_760),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_742),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_742),
.Y(n_790)
);

AOI221xp5_ASAP7_75t_L g791 ( 
.A1(n_779),
.A2(n_735),
.B1(n_740),
.B2(n_744),
.C(n_748),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_774),
.A2(n_740),
.B1(n_744),
.B2(n_749),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_773),
.A2(n_730),
.B1(n_741),
.B2(n_734),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_SL g794 ( 
.A1(n_776),
.A2(n_736),
.B1(n_747),
.B2(n_737),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_765),
.Y(n_796)
);

NAND4xp75_ASAP7_75t_L g797 ( 
.A(n_789),
.B(n_757),
.C(n_745),
.D(n_701),
.Y(n_797)
);

OA22x2_ASAP7_75t_L g798 ( 
.A1(n_774),
.A2(n_747),
.B1(n_736),
.B2(n_750),
.Y(n_798)
);

NAND4xp75_ASAP7_75t_L g799 ( 
.A(n_789),
.B(n_745),
.C(n_741),
.D(n_758),
.Y(n_799)
);

AOI32xp33_ASAP7_75t_L g800 ( 
.A1(n_784),
.A2(n_758),
.A3(n_696),
.B1(n_699),
.B2(n_733),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_766),
.Y(n_801)
);

NAND4xp25_ASAP7_75t_SL g802 ( 
.A(n_785),
.B(n_702),
.C(n_645),
.D(n_726),
.Y(n_802)
);

OA22x2_ASAP7_75t_L g803 ( 
.A1(n_762),
.A2(n_726),
.B1(n_694),
.B2(n_700),
.Y(n_803)
);

OAI322xp33_ASAP7_75t_L g804 ( 
.A1(n_790),
.A2(n_692),
.A3(n_695),
.B1(n_700),
.B2(n_684),
.C1(n_683),
.C2(n_710),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_772),
.B(n_720),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_766),
.Y(n_806)
);

NAND4xp25_ASAP7_75t_L g807 ( 
.A(n_767),
.B(n_694),
.C(n_649),
.D(n_648),
.Y(n_807)
);

NOR4xp25_ASAP7_75t_L g808 ( 
.A(n_762),
.B(n_695),
.C(n_684),
.D(n_683),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_786),
.Y(n_809)
);

OA22x2_ASAP7_75t_L g810 ( 
.A1(n_787),
.A2(n_723),
.B1(n_708),
.B2(n_698),
.Y(n_810)
);

INVx1_ASAP7_75t_SL g811 ( 
.A(n_780),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_768),
.Y(n_812)
);

AOI221xp5_ASAP7_75t_L g813 ( 
.A1(n_788),
.A2(n_708),
.B1(n_669),
.B2(n_645),
.C(n_717),
.Y(n_813)
);

OA22x2_ASAP7_75t_L g814 ( 
.A1(n_777),
.A2(n_669),
.B1(n_717),
.B2(n_152),
.Y(n_814)
);

AOI221xp5_ASAP7_75t_L g815 ( 
.A1(n_771),
.A2(n_79),
.B1(n_152),
.B2(n_153),
.C(n_158),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_771),
.A2(n_202),
.B(n_152),
.C(n_153),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_778),
.A2(n_152),
.B1(n_158),
.B2(n_190),
.Y(n_817)
);

OAI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_768),
.A2(n_169),
.B1(n_202),
.B2(n_258),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_795),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_791),
.A2(n_769),
.B1(n_770),
.B2(n_763),
.Y(n_820)
);

OAI22xp5_ASAP7_75t_L g821 ( 
.A1(n_793),
.A2(n_783),
.B1(n_775),
.B2(n_764),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_792),
.A2(n_782),
.B1(n_781),
.B2(n_190),
.Y(n_822)
);

AO22x2_ASAP7_75t_L g823 ( 
.A1(n_809),
.A2(n_258),
.B1(n_276),
.B2(n_266),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_795),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_796),
.Y(n_825)
);

AOI22x1_ASAP7_75t_L g826 ( 
.A1(n_811),
.A2(n_253),
.B1(n_158),
.B2(n_277),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_SL g827 ( 
.A1(n_800),
.A2(n_216),
.B(n_191),
.C(n_266),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_801),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_806),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_799),
.A2(n_253),
.B1(n_216),
.B2(n_197),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_803),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_SL g832 ( 
.A1(n_812),
.A2(n_216),
.B(n_191),
.C(n_176),
.Y(n_832)
);

AOI221xp5_ASAP7_75t_L g833 ( 
.A1(n_808),
.A2(n_79),
.B1(n_201),
.B2(n_175),
.C(n_183),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_797),
.A2(n_253),
.B1(n_216),
.B2(n_191),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_805),
.Y(n_835)
);

AOI22x1_ASAP7_75t_L g836 ( 
.A1(n_794),
.A2(n_253),
.B1(n_277),
.B2(n_249),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_817),
.Y(n_837)
);

AOI221xp5_ASAP7_75t_L g838 ( 
.A1(n_804),
.A2(n_79),
.B1(n_201),
.B2(n_175),
.C(n_183),
.Y(n_838)
);

OA22x2_ASAP7_75t_L g839 ( 
.A1(n_798),
.A2(n_810),
.B1(n_802),
.B2(n_814),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_818),
.Y(n_840)
);

AOI221xp5_ASAP7_75t_L g841 ( 
.A1(n_813),
.A2(n_79),
.B1(n_201),
.B2(n_175),
.C(n_186),
.Y(n_841)
);

AOI31xp33_ASAP7_75t_L g842 ( 
.A1(n_815),
.A2(n_277),
.A3(n_249),
.B(n_206),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_816),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_807),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_793),
.A2(n_186),
.B(n_206),
.C(n_277),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_821),
.A2(n_190),
.B1(n_201),
.B2(n_169),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_835),
.B(n_79),
.Y(n_847)
);

AOI221xp5_ASAP7_75t_L g848 ( 
.A1(n_834),
.A2(n_79),
.B1(n_216),
.B2(n_206),
.C(n_191),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_819),
.Y(n_849)
);

AO22x2_ASAP7_75t_L g850 ( 
.A1(n_825),
.A2(n_169),
.B1(n_172),
.B2(n_253),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_822),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_824),
.Y(n_852)
);

AOI221xp5_ASAP7_75t_L g853 ( 
.A1(n_845),
.A2(n_79),
.B1(n_216),
.B2(n_191),
.C(n_199),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_820),
.Y(n_854)
);

NOR4xp25_ASAP7_75t_L g855 ( 
.A(n_828),
.B(n_216),
.C(n_199),
.D(n_191),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_839),
.A2(n_190),
.B1(n_169),
.B2(n_219),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_829),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_831),
.A2(n_190),
.B1(n_169),
.B2(n_219),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_837),
.B(n_79),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_823),
.Y(n_860)
);

NOR4xp25_ASAP7_75t_L g861 ( 
.A(n_844),
.B(n_199),
.C(n_191),
.D(n_215),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_822),
.B(n_79),
.Y(n_862)
);

NOR2xp67_ASAP7_75t_L g863 ( 
.A(n_857),
.B(n_820),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_854),
.A2(n_830),
.B1(n_838),
.B2(n_841),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_851),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_861),
.B(n_840),
.Y(n_866)
);

NOR2xp67_ASAP7_75t_L g867 ( 
.A(n_856),
.B(n_852),
.Y(n_867)
);

AO22x2_ASAP7_75t_L g868 ( 
.A1(n_849),
.A2(n_843),
.B1(n_827),
.B2(n_836),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_847),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_862),
.A2(n_833),
.B1(n_823),
.B2(n_842),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_860),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_859),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_858),
.A2(n_842),
.B1(n_832),
.B2(n_826),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_846),
.B(n_855),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_850),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_865),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_863),
.A2(n_853),
.B1(n_850),
.B2(n_848),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_868),
.Y(n_878)
);

NAND4xp25_ASAP7_75t_L g879 ( 
.A(n_867),
.B(n_169),
.C(n_215),
.D(n_190),
.Y(n_879)
);

AND4x1_ASAP7_75t_L g880 ( 
.A(n_864),
.B(n_215),
.C(n_249),
.D(n_218),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_866),
.B(n_199),
.Y(n_881)
);

NAND4xp25_ASAP7_75t_L g882 ( 
.A(n_874),
.B(n_249),
.C(n_218),
.D(n_219),
.Y(n_882)
);

NOR2x1_ASAP7_75t_L g883 ( 
.A(n_875),
.B(n_218),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_868),
.Y(n_884)
);

NAND4xp25_ASAP7_75t_L g885 ( 
.A(n_873),
.B(n_219),
.C(n_141),
.D(n_79),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_871),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_872),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_876),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_881),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_879),
.B(n_869),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_878),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_884),
.A2(n_870),
.B1(n_219),
.B2(n_79),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_886),
.Y(n_893)
);

OAI211xp5_ASAP7_75t_L g894 ( 
.A1(n_877),
.A2(n_882),
.B(n_885),
.C(n_887),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_883),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_893),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_891),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_892),
.A2(n_894),
.B1(n_888),
.B2(n_890),
.Y(n_898)
);

AO22x2_ASAP7_75t_L g899 ( 
.A1(n_888),
.A2(n_880),
.B1(n_172),
.B2(n_219),
.Y(n_899)
);

OAI22x1_ASAP7_75t_L g900 ( 
.A1(n_889),
.A2(n_172),
.B1(n_219),
.B2(n_141),
.Y(n_900)
);

AND4x2_ASAP7_75t_L g901 ( 
.A(n_895),
.B(n_219),
.C(n_141),
.D(n_79),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_896),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_897),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_901),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_898),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_SL g906 ( 
.A1(n_903),
.A2(n_900),
.B1(n_899),
.B2(n_219),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_906),
.Y(n_907)
);

AO22x2_ASAP7_75t_L g908 ( 
.A1(n_907),
.A2(n_902),
.B1(n_904),
.B2(n_905),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_908),
.Y(n_909)
);

AOI221xp5_ASAP7_75t_L g910 ( 
.A1(n_909),
.A2(n_79),
.B1(n_141),
.B2(n_219),
.C(n_897),
.Y(n_910)
);

AOI211xp5_ASAP7_75t_L g911 ( 
.A1(n_910),
.A2(n_79),
.B(n_219),
.C(n_141),
.Y(n_911)
);


endmodule