module fake_jpeg_836_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_27),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_24),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_25),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_53),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_22),
.B1(n_17),
.B2(n_20),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_34),
.B(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_26),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_0),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_33),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_18),
.B1(n_26),
.B2(n_13),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_59),
.B(n_17),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_41),
.B1(n_32),
.B2(n_30),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_16),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_20),
.C(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_65),
.B(n_66),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_71),
.B(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_69),
.Y(n_92)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_13),
.B(n_1),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_5),
.C(n_9),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_58),
.B1(n_43),
.B2(n_59),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_48),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_1),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_61),
.B(n_62),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_86),
.B(n_67),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_50),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_79),
.C(n_73),
.Y(n_97)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_4),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_60),
.B1(n_46),
.B2(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_98),
.C(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_104),
.Y(n_106)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_74),
.C(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_72),
.B(n_70),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_94),
.B(n_46),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_87),
.B1(n_85),
.B2(n_82),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_108),
.B(n_90),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_103),
.B(n_98),
.C(n_82),
.D(n_95),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_111),
.B(n_113),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_92),
.B(n_69),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_116),
.B(n_118),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_84),
.C(n_60),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_119),
.B(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_124),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_129),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_118),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_127),
.A2(n_122),
.B(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_119),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_131),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_124),
.B(n_107),
.Y(n_134)
);


endmodule