module fake_jpeg_1893_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_58),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_68),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_40),
.B1(n_37),
.B2(n_43),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_69),
.B1(n_55),
.B2(n_56),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_40),
.B1(n_50),
.B2(n_48),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_54),
.B1(n_47),
.B2(n_45),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_57),
.B(n_37),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_79),
.B1(n_51),
.B2(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_20),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_0),
.B(n_1),
.C(n_4),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_22),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_87),
.B1(n_91),
.B2(n_5),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_62),
.B1(n_1),
.B2(n_3),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_35),
.B(n_16),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_25),
.B(n_30),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_82),
.B1(n_80),
.B2(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_93),
.B(n_98),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_97),
.B(n_23),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_5),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_100),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_105),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_104),
.B1(n_10),
.B2(n_11),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_104)
);

FAx1_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_7),
.CI(n_8),
.CON(n_105),
.SN(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_24),
.C(n_29),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_13),
.C(n_18),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_123),
.B(n_114),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_10),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_114),
.A2(n_105),
.B1(n_112),
.B2(n_32),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_26),
.B1(n_27),
.B2(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_132),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_105),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_118),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_121),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_131),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_140),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_138),
.A2(n_117),
.B1(n_119),
.B2(n_130),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_142),
.B(n_133),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_135),
.B(n_136),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_125),
.C(n_126),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_145),
.Y(n_146)
);


endmodule