module fake_ibex_581_n_3895 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_602, n_355, n_474, n_594, n_407, n_102, n_490, n_568, n_52, n_448, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_267, n_245, n_589, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_3895);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_267;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3895;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_766;
wire n_3590;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_3559;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_3817;
wire n_773;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_1652;
wire n_678;
wire n_969;
wire n_1954;
wire n_1859;
wire n_2183;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_2640;
wire n_1666;
wire n_2682;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_2720;
wire n_3870;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_667;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3729;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_671;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_641;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_694;
wire n_787;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3884;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_917;
wire n_2413;
wire n_3022;
wire n_2362;
wire n_968;
wire n_2249;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_666;
wire n_2260;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_662;
wire n_3097;
wire n_2906;
wire n_3030;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_3822;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_772;
wire n_810;
wire n_1401;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_630;
wire n_1869;
wire n_3842;
wire n_2275;
wire n_1853;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3780;
wire n_3023;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_1969;
wire n_3798;
wire n_709;
wire n_1296;
wire n_3060;
wire n_971;
wire n_702;
wire n_1326;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_1506;
wire n_881;
wire n_2987;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_3630;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2625;
wire n_1742;
wire n_2350;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3800;
wire n_3887;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_3583;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_657;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_3448;
wire n_3634;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2599;
wire n_974;
wire n_1036;
wire n_2076;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_738;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_3813;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2585;
wire n_2220;
wire n_2080;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_669;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_724;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_2999;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_660;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_705;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2699;
wire n_2160;
wire n_2234;
wire n_2991;
wire n_847;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_3797;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3880;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_3087;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_3070;
wire n_2711;
wire n_2842;
wire n_3477;
wire n_650;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2612;
wire n_2193;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_633;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2716;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_668;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_774;
wire n_3137;
wire n_2459;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_1185;
wire n_1683;
wire n_3575;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_687;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_3158;
wire n_1535;
wire n_2985;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_2127;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_3632;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3608;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_673;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_785;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3818;
wire n_642;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_2959;
wire n_1625;
wire n_2610;
wire n_2380;
wire n_2420;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_636;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_659;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_648;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_3645;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_768;
wire n_3705;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_3743;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2447;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_685;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3538;
wire n_1261;
wire n_2299;
wire n_3393;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_681;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1989;
wire n_1740;
wire n_3540;
wire n_1838;
wire n_3649;
wire n_833;
wire n_3604;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_3740;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2576;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_2229;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_631;
wire n_794;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_3066;
wire n_2714;
wire n_2669;
wire n_697;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2898;
wire n_3121;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3576;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2864;
wire n_2406;
wire n_1632;
wire n_3346;
wire n_688;
wire n_3104;
wire n_3391;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_3014;
wire n_1812;
wire n_2703;
wire n_1951;
wire n_1330;
wire n_638;
wire n_2574;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_3102;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_682;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3343;
wire n_3163;
wire n_3752;
wire n_3786;
wire n_632;
wire n_1329;
wire n_2637;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_2914;
wire n_1833;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_665;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_654;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_2734;
wire n_2870;
wire n_758;
wire n_1166;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1992;
wire n_1685;
wire n_1784;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3380;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_635;
wire n_3837;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2706;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2303;
wire n_704;
wire n_2357;
wire n_2653;
wire n_2855;
wire n_2618;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_699;
wire n_2136;
wire n_3617;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_3056;
wire n_2560;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2802;
wire n_2443;
wire n_3052;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2066;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_3613;
wire n_627;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_1059;
wire n_2969;
wire n_799;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_691;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2738;
wire n_2324;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2619;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_952;
wire n_1947;
wire n_1675;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_3793;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_680;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_3635;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_683;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1849;
wire n_1674;
wire n_686;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_3482;
wire n_2282;
wire n_970;
wire n_3654;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_3677;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_649;
wire n_1854;
wire n_866;

INVx2_ASAP7_75t_L g627 ( 
.A(n_438),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_587),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_336),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_384),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_258),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_360),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_574),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_233),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_107),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_247),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_405),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_167),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_538),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_460),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_82),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_238),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_583),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_474),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_368),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_346),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_250),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_277),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_332),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_612),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_85),
.Y(n_651)
);

CKINVDCx16_ASAP7_75t_R g652 ( 
.A(n_146),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_434),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_544),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_282),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_461),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_405),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_277),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_542),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_269),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_453),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_516),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_611),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_205),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_390),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_397),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_455),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_471),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_565),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_316),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_472),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_296),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_366),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_265),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_33),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_82),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_605),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_344),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_465),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_599),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_50),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_543),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_487),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_40),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_357),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_143),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_110),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_531),
.Y(n_688)
);

INVx1_ASAP7_75t_SL g689 ( 
.A(n_290),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_499),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_429),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_618),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_107),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_123),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_491),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_579),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_262),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_591),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_325),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_339),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_488),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_614),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_409),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_539),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_426),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_590),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_227),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_311),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_554),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_215),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_354),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_560),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_385),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_240),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_276),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_323),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_210),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_86),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_398),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_541),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_511),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_261),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_409),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_14),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_69),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_330),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_6),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_520),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_423),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_533),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_23),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_27),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_593),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_254),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_449),
.Y(n_736)
);

CKINVDCx16_ASAP7_75t_R g737 ( 
.A(n_434),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_473),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_601),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_395),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_96),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_108),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_546),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_260),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_110),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_494),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_255),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_447),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_470),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_154),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_41),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_553),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_563),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_414),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_3),
.Y(n_755)
);

BUFx10_ASAP7_75t_L g756 ( 
.A(n_54),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_55),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_167),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_257),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_596),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_34),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_576),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_548),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_336),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_317),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_431),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_24),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_422),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_11),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_248),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_358),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_506),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_535),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_91),
.Y(n_774)
);

BUFx8_ASAP7_75t_SL g775 ( 
.A(n_514),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_575),
.Y(n_776)
);

CKINVDCx20_ASAP7_75t_R g777 ( 
.A(n_294),
.Y(n_777)
);

INVx1_ASAP7_75t_SL g778 ( 
.A(n_365),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_432),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_94),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_312),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_418),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_316),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_422),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_411),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_589),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_67),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_441),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_36),
.Y(n_789)
);

INVxp33_ASAP7_75t_L g790 ( 
.A(n_132),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_255),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_328),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_522),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_7),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_372),
.Y(n_795)
);

CKINVDCx16_ASAP7_75t_R g796 ( 
.A(n_220),
.Y(n_796)
);

CKINVDCx16_ASAP7_75t_R g797 ( 
.A(n_432),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_608),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_257),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_588),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_143),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_11),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_214),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_352),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_594),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_166),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_561),
.Y(n_807)
);

INVx4_ASAP7_75t_R g808 ( 
.A(n_44),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_549),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_467),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_363),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_101),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_584),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_341),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_534),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_325),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_384),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_305),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_149),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_18),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_557),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_429),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_326),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_99),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_392),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_387),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_99),
.Y(n_827)
);

BUFx10_ASAP7_75t_L g828 ( 
.A(n_420),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_199),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_477),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_617),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_62),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_288),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_622),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_509),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_572),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_613),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_463),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_625),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_624),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_357),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_370),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_479),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_502),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_49),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_540),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_192),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_515),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_585),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_597),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_537),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_125),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_210),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_450),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_265),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_559),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_430),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_163),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_389),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_567),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_507),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_555),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_359),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_228),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_104),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_407),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_343),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_447),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_112),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_231),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_151),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_245),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_475),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_510),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_476),
.Y(n_875)
);

INVxp33_ASAP7_75t_R g876 ( 
.A(n_568),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_426),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_527),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_105),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_436),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_19),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_349),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_562),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_252),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_84),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_183),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_222),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_262),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_238),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_564),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_279),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_513),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_620),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_127),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_37),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_312),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_545),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_338),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_281),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_402),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_603),
.Y(n_901)
);

INVxp67_ASAP7_75t_SL g902 ( 
.A(n_291),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_343),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_602),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_421),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_570),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_455),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_486),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_586),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_324),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_207),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_604),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_610),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_609),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_102),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_164),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_293),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_247),
.Y(n_918)
);

CKINVDCx16_ASAP7_75t_R g919 ( 
.A(n_169),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_64),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_550),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_300),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_227),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_382),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_615),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_230),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_108),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_297),
.Y(n_928)
);

BUFx10_ASAP7_75t_L g929 ( 
.A(n_306),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_421),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_106),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_235),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_370),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_517),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_285),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_442),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_58),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_412),
.Y(n_938)
);

INVxp33_ASAP7_75t_SL g939 ( 
.A(n_378),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_349),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_49),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_88),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_245),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_360),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_48),
.Y(n_945)
);

CKINVDCx14_ASAP7_75t_R g946 ( 
.A(n_418),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_623),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_441),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_61),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_218),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_472),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_361),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_321),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_371),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_296),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_461),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_87),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_26),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_577),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_20),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_135),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_462),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_263),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_205),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_592),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_621),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_182),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_188),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_595),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_453),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_307),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_600),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_484),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_356),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_606),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_113),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_214),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_52),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_165),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_571),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_232),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_268),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_211),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_243),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_104),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_393),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_149),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_607),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_109),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_35),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_242),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_341),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_204),
.Y(n_993)
);

CKINVDCx14_ASAP7_75t_R g994 ( 
.A(n_566),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_45),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_414),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_556),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_254),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_151),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_392),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_221),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_573),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_72),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_124),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_578),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_273),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_241),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_308),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_598),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_322),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_311),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_303),
.Y(n_1012)
);

BUFx10_ASAP7_75t_L g1013 ( 
.A(n_145),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_505),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_582),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_358),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_581),
.Y(n_1017)
);

CKINVDCx20_ASAP7_75t_R g1018 ( 
.A(n_498),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_334),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_310),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_148),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_278),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_134),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_309),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_0),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_404),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_188),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_204),
.Y(n_1028)
);

BUFx2_ASAP7_75t_SL g1029 ( 
.A(n_309),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_114),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_536),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_552),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_569),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_440),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_484),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_551),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_580),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_547),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_213),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_121),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_96),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_403),
.Y(n_1042)
);

BUFx10_ASAP7_75t_L g1043 ( 
.A(n_492),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_619),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_532),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_83),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_31),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_346),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_366),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_388),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_127),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_914),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_839),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_627),
.Y(n_1054)
);

BUFx3_ASAP7_75t_L g1055 ( 
.A(n_1043),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_706),
.B(n_1),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_914),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_627),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_651),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_766),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_914),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_887),
.B(n_1),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_914),
.Y(n_1063)
);

INVx5_ASAP7_75t_L g1064 ( 
.A(n_839),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_790),
.B(n_0),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_651),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_839),
.B(n_2),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_936),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_649),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_675),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_637),
.B(n_2),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_SL g1072 ( 
.A(n_775),
.B(n_626),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_637),
.B(n_3),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_764),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_649),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_764),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_671),
.B(n_4),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_671),
.B(n_4),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_685),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_685),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_993),
.B(n_6),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_995),
.B(n_7),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1004),
.B(n_8),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_675),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_736),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_790),
.B(n_652),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_675),
.Y(n_1087)
);

BUFx8_ASAP7_75t_SL g1088 ( 
.A(n_638),
.Y(n_1088)
);

CKINVDCx14_ASAP7_75t_R g1089 ( 
.A(n_946),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1045),
.B(n_8),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_675),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_1043),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_676),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_1043),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_713),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_680),
.Y(n_1096)
);

BUFx12f_ASAP7_75t_L g1097 ( 
.A(n_649),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_687),
.B(n_979),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_687),
.B(n_9),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_769),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_979),
.B(n_5),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_737),
.B(n_5),
.Y(n_1102)
);

INVx5_ASAP7_75t_L g1103 ( 
.A(n_908),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_658),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_676),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_676),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_796),
.B(n_9),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_713),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_736),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_908),
.B(n_10),
.Y(n_1110)
);

BUFx8_ASAP7_75t_L g1111 ( 
.A(n_1009),
.Y(n_1111)
);

INVxp33_ASAP7_75t_SL g1112 ( 
.A(n_658),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_749),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_749),
.B(n_10),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1009),
.B(n_12),
.Y(n_1115)
);

BUFx8_ASAP7_75t_L g1116 ( 
.A(n_767),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_769),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_797),
.B(n_12),
.Y(n_1118)
);

BUFx8_ASAP7_75t_SL g1119 ( 
.A(n_638),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_676),
.Y(n_1120)
);

INVx5_ASAP7_75t_L g1121 ( 
.A(n_742),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_905),
.B(n_13),
.Y(n_1122)
);

BUFx8_ASAP7_75t_SL g1123 ( 
.A(n_642),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_628),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_739),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_919),
.B(n_14),
.Y(n_1126)
);

INVx5_ASAP7_75t_L g1127 ( 
.A(n_742),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_663),
.B(n_13),
.Y(n_1128)
);

BUFx8_ASAP7_75t_SL g1129 ( 
.A(n_642),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_660),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_660),
.B(n_16),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_742),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_661),
.B(n_16),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_742),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_730),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_879),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_661),
.B(n_664),
.Y(n_1137)
);

AND2x6_ASAP7_75t_L g1138 ( 
.A(n_739),
.B(n_616),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_730),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_682),
.B(n_15),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_730),
.B(n_15),
.Y(n_1141)
);

INVxp33_ASAP7_75t_SL g1142 ( 
.A(n_664),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_756),
.B(n_17),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_756),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_879),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_767),
.B(n_17),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_879),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_879),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_918),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_859),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_859),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_918),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_639),
.Y(n_1153)
);

INVx5_ASAP7_75t_L g1154 ( 
.A(n_918),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_918),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_668),
.B(n_19),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_877),
.B(n_18),
.Y(n_1157)
);

INVx1_ASAP7_75t_SL g1158 ( 
.A(n_1112),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1079),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1086),
.B(n_901),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1094),
.B(n_925),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1094),
.B(n_1124),
.Y(n_1162)
);

OAI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1072),
.A2(n_670),
.B1(n_672),
.B2(n_668),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1060),
.B(n_994),
.Y(n_1164)
);

INVx8_ASAP7_75t_L g1165 ( 
.A(n_1075),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1124),
.B(n_670),
.Y(n_1166)
);

AOI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1080),
.A2(n_705),
.B1(n_734),
.B2(n_703),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1068),
.B(n_756),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_1065),
.B(n_876),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1142),
.A2(n_939),
.B1(n_654),
.B2(n_662),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1089),
.B(n_1104),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1071),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1096),
.A2(n_939),
.B1(n_654),
.B2(n_662),
.Y(n_1173)
);

OAI22xp33_ASAP7_75t_R g1174 ( 
.A1(n_1102),
.A2(n_902),
.B1(n_686),
.B2(n_689),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1130),
.B(n_828),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1137),
.A2(n_672),
.B1(n_1011),
.B2(n_1010),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_SL g1177 ( 
.A(n_1097),
.B(n_775),
.Y(n_1177)
);

AOI22x1_ASAP7_75t_SL g1178 ( 
.A1(n_1088),
.A2(n_759),
.B1(n_765),
.B2(n_744),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1094),
.B(n_690),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1153),
.B(n_1010),
.Y(n_1180)
);

OAI22xp33_ASAP7_75t_SL g1181 ( 
.A1(n_1126),
.A2(n_1012),
.B1(n_1011),
.B2(n_630),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1131),
.A2(n_1012),
.B1(n_631),
.B2(n_632),
.Y(n_1182)
);

INVx8_ASAP7_75t_L g1183 ( 
.A(n_1139),
.Y(n_1183)
);

OAI22xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1133),
.A2(n_634),
.B1(n_635),
.B2(n_629),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1055),
.B(n_659),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1144),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1098),
.Y(n_1187)
);

OAI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1056),
.A2(n_759),
.B1(n_765),
.B2(n_744),
.Y(n_1188)
);

OAI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1062),
.A2(n_1081),
.B1(n_1083),
.B2(n_1082),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1107),
.A2(n_1122),
.B1(n_1118),
.B2(n_1073),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1071),
.A2(n_677),
.B1(n_743),
.B2(n_633),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1085),
.Y(n_1192)
);

OA22x2_ASAP7_75t_L g1193 ( 
.A1(n_1069),
.A2(n_1029),
.B1(n_636),
.B2(n_712),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1109),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1073),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1092),
.B(n_828),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1077),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1113),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1153),
.Y(n_1199)
);

OAI22xp33_ASAP7_75t_R g1200 ( 
.A1(n_1119),
.A2(n_718),
.B1(n_745),
.B2(n_684),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1150),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_1077),
.A2(n_1101),
.B1(n_1078),
.B2(n_1114),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_1135),
.B(n_659),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_SL g1204 ( 
.A1(n_1123),
.A2(n_810),
.B1(n_854),
.B2(n_777),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1111),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1156),
.A2(n_810),
.B1(n_854),
.B2(n_777),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1078),
.A2(n_677),
.B1(n_743),
.B2(n_633),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1101),
.A2(n_805),
.B1(n_846),
.B2(n_798),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1114),
.Y(n_1209)
);

OAI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1090),
.A2(n_938),
.B1(n_976),
.B2(n_870),
.Y(n_1210)
);

OAI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1099),
.A2(n_938),
.B1(n_976),
.B2(n_870),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1146),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1151),
.Y(n_1213)
);

OAI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1146),
.A2(n_646),
.B1(n_647),
.B2(n_644),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1095),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1157),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1157),
.A2(n_805),
.B1(n_846),
.B2(n_798),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1098),
.A2(n_1017),
.B1(n_1018),
.B2(n_878),
.Y(n_1218)
);

INVx6_ASAP7_75t_L g1219 ( 
.A(n_1116),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1054),
.A2(n_655),
.B1(n_673),
.B2(n_653),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1108),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1141),
.A2(n_1030),
.B1(n_1025),
.B2(n_1017),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1129),
.A2(n_1030),
.B1(n_1025),
.B2(n_1018),
.Y(n_1223)
);

AO22x2_ASAP7_75t_L g1224 ( 
.A1(n_1143),
.A2(n_812),
.B1(n_819),
.B2(n_778),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1054),
.A2(n_681),
.B1(n_691),
.B2(n_679),
.Y(n_1225)
);

OAI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1058),
.A2(n_698),
.B1(n_704),
.B2(n_693),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1125),
.Y(n_1227)
);

OA22x2_ASAP7_75t_L g1228 ( 
.A1(n_1058),
.A2(n_758),
.B1(n_783),
.B2(n_724),
.Y(n_1228)
);

AND2x2_ASAP7_75t_SL g1229 ( 
.A(n_1110),
.B(n_794),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1053),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1121),
.Y(n_1231)
);

AO22x2_ASAP7_75t_L g1232 ( 
.A1(n_1059),
.A2(n_948),
.B1(n_960),
.B2(n_911),
.Y(n_1232)
);

OAI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1053),
.A2(n_878),
.B1(n_641),
.B2(n_645),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_SL g1234 ( 
.A1(n_1128),
.A2(n_709),
.B1(n_711),
.B2(n_708),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1053),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1116),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1111),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1121),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1115),
.A2(n_717),
.B1(n_719),
.B2(n_716),
.Y(n_1239)
);

AO22x2_ASAP7_75t_L g1240 ( 
.A1(n_1059),
.A2(n_1051),
.B1(n_648),
.B2(n_656),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1064),
.B(n_877),
.Y(n_1241)
);

OAI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1066),
.A2(n_723),
.B1(n_725),
.B2(n_720),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_SL g1243 ( 
.A1(n_1066),
.A2(n_728),
.B1(n_735),
.B2(n_727),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1140),
.A2(n_741),
.B1(n_747),
.B2(n_740),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1064),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1121),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1064),
.Y(n_1247)
);

OAI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1074),
.A2(n_657),
.B1(n_665),
.B2(n_640),
.Y(n_1248)
);

OAI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1074),
.A2(n_751),
.B1(n_754),
.B2(n_750),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1076),
.A2(n_667),
.B1(n_674),
.B2(n_666),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1127),
.Y(n_1251)
);

OAI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1076),
.A2(n_678),
.B1(n_700),
.B2(n_694),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1100),
.B(n_828),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1127),
.Y(n_1254)
);

AO22x2_ASAP7_75t_L g1255 ( 
.A1(n_1100),
.A2(n_714),
.B1(n_715),
.B2(n_701),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1117),
.B(n_886),
.Y(n_1256)
);

AO22x2_ASAP7_75t_L g1257 ( 
.A1(n_1117),
.A2(n_1050),
.B1(n_1049),
.B2(n_732),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1127),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1138),
.A2(n_733),
.B1(n_738),
.B2(n_726),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1067),
.Y(n_1260)
);

INVx1_ASAP7_75t_SL g1261 ( 
.A(n_1103),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1103),
.A2(n_748),
.B1(n_757),
.B2(n_755),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1103),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1136),
.B(n_886),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1136),
.B(n_886),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1136),
.B(n_929),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1148),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1070),
.B(n_974),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1148),
.A2(n_761),
.B1(n_780),
.B2(n_779),
.Y(n_1269)
);

OAI22xp33_ASAP7_75t_L g1270 ( 
.A1(n_1148),
.A2(n_785),
.B1(n_791),
.B2(n_782),
.Y(n_1270)
);

AO22x2_ASAP7_75t_L g1271 ( 
.A1(n_1138),
.A2(n_795),
.B1(n_801),
.B2(n_799),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1154),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1154),
.B(n_929),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1138),
.A2(n_768),
.B1(n_771),
.B2(n_770),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1154),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1138),
.B(n_929),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1070),
.Y(n_1277)
);

AND2x2_ASAP7_75t_SL g1278 ( 
.A(n_1070),
.B(n_794),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1084),
.B(n_922),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1084),
.B(n_1013),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1084),
.A2(n_811),
.B1(n_814),
.B2(n_803),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1087),
.B(n_832),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1087),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1087),
.A2(n_774),
.B1(n_784),
.B2(n_781),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1091),
.B(n_843),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1091),
.A2(n_853),
.B1(n_855),
.B2(n_845),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1091),
.A2(n_787),
.B1(n_789),
.B2(n_788),
.Y(n_1287)
);

AOI22x1_ASAP7_75t_SL g1288 ( 
.A1(n_1093),
.A2(n_792),
.B1(n_804),
.B2(n_802),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1093),
.A2(n_806),
.B1(n_817),
.B2(n_816),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1093),
.Y(n_1290)
);

OAI22xp33_ASAP7_75t_R g1291 ( 
.A1(n_1105),
.A2(n_868),
.B1(n_875),
.B2(n_858),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_1105),
.B(n_922),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1105),
.A2(n_818),
.B1(n_822),
.B2(n_820),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1106),
.A2(n_823),
.B1(n_825),
.B2(n_824),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1106),
.B(n_1013),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1106),
.A2(n_826),
.B1(n_829),
.B2(n_827),
.Y(n_1296)
);

AND2x4_ASAP7_75t_L g1297 ( 
.A(n_1120),
.B(n_935),
.Y(n_1297)
);

OAI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1120),
.A2(n_881),
.B1(n_882),
.B2(n_880),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1120),
.A2(n_894),
.B1(n_896),
.B2(n_884),
.Y(n_1299)
);

AOI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1132),
.A2(n_830),
.B1(n_838),
.B2(n_833),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1132),
.A2(n_907),
.B1(n_910),
.B2(n_903),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1132),
.Y(n_1302)
);

OAI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1134),
.A2(n_841),
.B1(n_847),
.B2(n_842),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1134),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1134),
.B(n_1013),
.Y(n_1305)
);

AO22x2_ASAP7_75t_L g1306 ( 
.A1(n_1145),
.A2(n_1042),
.B1(n_924),
.B2(n_928),
.Y(n_1306)
);

AO22x2_ASAP7_75t_L g1307 ( 
.A1(n_1145),
.A2(n_943),
.B1(n_950),
.B2(n_923),
.Y(n_1307)
);

AOI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1145),
.A2(n_852),
.B1(n_863),
.B2(n_857),
.Y(n_1308)
);

OAI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1147),
.A2(n_952),
.B1(n_954),
.B2(n_951),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1147),
.B(n_1041),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1147),
.A2(n_864),
.B1(n_866),
.B2(n_865),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1149),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1149),
.A2(n_957),
.B1(n_982),
.B2(n_956),
.Y(n_1313)
);

AO22x2_ASAP7_75t_L g1314 ( 
.A1(n_1149),
.A2(n_984),
.B1(n_987),
.B2(n_983),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1152),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1152),
.A2(n_867),
.B1(n_871),
.B2(n_869),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1152),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1155),
.A2(n_872),
.B1(n_885),
.B2(n_873),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1155),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1155),
.Y(n_1320)
);

OAI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1052),
.A2(n_888),
.B1(n_891),
.B2(n_889),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_1052),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1052),
.B(n_1041),
.Y(n_1323)
);

OAI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1057),
.A2(n_895),
.B1(n_899),
.B2(n_898),
.Y(n_1324)
);

XNOR2xp5_ASAP7_75t_L g1325 ( 
.A(n_1063),
.B(n_900),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1063),
.B(n_935),
.Y(n_1326)
);

INVxp33_ASAP7_75t_L g1327 ( 
.A(n_1057),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1057),
.Y(n_1328)
);

AOI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1061),
.A2(n_920),
.B1(n_926),
.B2(n_917),
.Y(n_1329)
);

OA22x2_ASAP7_75t_L g1330 ( 
.A1(n_1061),
.A2(n_953),
.B1(n_973),
.B2(n_937),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1061),
.B(n_692),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1063),
.A2(n_990),
.B1(n_991),
.B2(n_989),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_SL g1333 ( 
.A(n_1071),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1086),
.B(n_962),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_R g1335 ( 
.A1(n_1102),
.A2(n_1021),
.B1(n_1026),
.B2(n_1020),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1075),
.Y(n_1336)
);

OR2x6_ASAP7_75t_L g1337 ( 
.A(n_1075),
.B(n_1046),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1112),
.A2(n_927),
.B1(n_931),
.B2(n_930),
.Y(n_1338)
);

INVx2_ASAP7_75t_SL g1339 ( 
.A(n_1094),
.Y(n_1339)
);

AO22x2_ASAP7_75t_L g1340 ( 
.A1(n_1086),
.A2(n_1035),
.B1(n_1027),
.B2(n_916),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1086),
.A2(n_933),
.B1(n_940),
.B2(n_932),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1071),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1072),
.A2(n_1048),
.B1(n_1047),
.B2(n_944),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1060),
.B(n_962),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1086),
.A2(n_945),
.B1(n_949),
.B2(n_941),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1086),
.A2(n_961),
.B1(n_963),
.B2(n_958),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1072),
.A2(n_1040),
.B1(n_1034),
.B2(n_967),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1086),
.A2(n_968),
.B1(n_970),
.B2(n_964),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1072),
.A2(n_977),
.B1(n_978),
.B2(n_971),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1086),
.B(n_998),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1086),
.B(n_998),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1086),
.A2(n_985),
.B1(n_986),
.B2(n_981),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1075),
.Y(n_1353)
);

AO22x2_ASAP7_75t_L g1354 ( 
.A1(n_1086),
.A2(n_916),
.B1(n_942),
.B2(n_915),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1079),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1098),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1086),
.A2(n_996),
.B1(n_999),
.B2(n_992),
.Y(n_1357)
);

OR2x6_ASAP7_75t_L g1358 ( 
.A(n_1075),
.B(n_1046),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1094),
.B(n_697),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1071),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1218),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1356),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1282),
.Y(n_1363)
);

INVxp33_ASAP7_75t_L g1364 ( 
.A(n_1338),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1285),
.Y(n_1365)
);

INVxp33_ASAP7_75t_L g1366 ( 
.A(n_1168),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1202),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1306),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1164),
.B(n_1158),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1202),
.Y(n_1370)
);

AOI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1259),
.A2(n_721),
.B(n_702),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1160),
.B(n_1253),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1354),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1354),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1256),
.B(n_1001),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1187),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1173),
.B(n_1003),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1280),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1268),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1295),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1305),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1165),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_SL g1383 ( 
.A(n_1205),
.B(n_669),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1175),
.B(n_1008),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1274),
.B(n_497),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1241),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1260),
.A2(n_746),
.B(n_731),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1241),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1279),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1170),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1279),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1172),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1195),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1197),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1342),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1165),
.Y(n_1396)
);

XOR2xp5_ASAP7_75t_L g1397 ( 
.A(n_1178),
.B(n_1019),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1360),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1292),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1159),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1166),
.B(n_669),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1192),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1180),
.B(n_1014),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1292),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1334),
.B(n_1016),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1194),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1198),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1408)
);

CKINVDCx20_ASAP7_75t_R g1409 ( 
.A(n_1223),
.Y(n_1409)
);

NAND2xp33_ASAP7_75t_SL g1410 ( 
.A(n_1237),
.B(n_1014),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1297),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1201),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1268),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1213),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1355),
.Y(n_1415)
);

NOR2xp33_ASAP7_75t_L g1416 ( 
.A(n_1199),
.B(n_772),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1297),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1310),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1240),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1240),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1255),
.Y(n_1421)
);

INVxp33_ASAP7_75t_L g1422 ( 
.A(n_1325),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1255),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_1186),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1257),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1183),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1344),
.B(n_1022),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1323),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1257),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1306),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1196),
.B(n_915),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1183),
.B(n_1023),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1171),
.B(n_1028),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1340),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1326),
.Y(n_1436)
);

XNOR2xp5_ASAP7_75t_L g1437 ( 
.A(n_1169),
.B(n_20),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1176),
.B(n_942),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1278),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1307),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1204),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1230),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1199),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1307),
.Y(n_1444)
);

XOR2xp5_ASAP7_75t_L g1445 ( 
.A(n_1191),
.B(n_21),
.Y(n_1445)
);

INVx4_ASAP7_75t_SL g1446 ( 
.A(n_1219),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1314),
.Y(n_1447)
);

INVxp33_ASAP7_75t_L g1448 ( 
.A(n_1236),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1190),
.B(n_955),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1203),
.B(n_893),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1231),
.Y(n_1451)
);

INVxp33_ASAP7_75t_L g1452 ( 
.A(n_1177),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1185),
.B(n_909),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1235),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1189),
.B(n_643),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1161),
.B(n_650),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1314),
.Y(n_1457)
);

AND2x6_ASAP7_75t_L g1458 ( 
.A(n_1276),
.B(n_760),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1245),
.Y(n_1459)
);

CKINVDCx20_ASAP7_75t_R g1460 ( 
.A(n_1219),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_SL g1461 ( 
.A(n_1336),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1209),
.A2(n_705),
.B(n_703),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1212),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1353),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1247),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1216),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1215),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1333),
.B(n_683),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1221),
.Y(n_1469)
);

XOR2xp5_ASAP7_75t_L g1470 ( 
.A(n_1207),
.B(n_21),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1259),
.A2(n_809),
.B(n_734),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1208),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1227),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1217),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1261),
.B(n_1264),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1265),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1266),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1273),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1228),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1337),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1229),
.B(n_776),
.Y(n_1481)
);

XOR2xp5_ASAP7_75t_L g1482 ( 
.A(n_1222),
.B(n_22),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1330),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1167),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1193),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1339),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1190),
.B(n_955),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1337),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1332),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1238),
.Y(n_1490)
);

XOR2xp5_ASAP7_75t_L g1491 ( 
.A(n_1206),
.B(n_22),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1281),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1286),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1358),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_SL g1495 ( 
.A(n_1358),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1271),
.B(n_786),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1298),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1341),
.B(n_1346),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1299),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1271),
.A2(n_837),
.B(n_809),
.Y(n_1500)
);

XOR2xp5_ASAP7_75t_L g1501 ( 
.A(n_1188),
.B(n_23),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1301),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1214),
.B(n_688),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1348),
.B(n_974),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1309),
.Y(n_1505)
);

XOR2xp5_ASAP7_75t_L g1506 ( 
.A(n_1210),
.B(n_24),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_SL g1507 ( 
.A(n_1163),
.B(n_1343),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1288),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_1267),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1313),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1239),
.B(n_696),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1345),
.A2(n_849),
.B(n_837),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1263),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1357),
.B(n_1024),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1291),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1352),
.B(n_699),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1291),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1275),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1269),
.Y(n_1519)
);

XOR2x2_ASAP7_75t_L g1520 ( 
.A(n_1181),
.B(n_25),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1284),
.Y(n_1521)
);

INVx4_ASAP7_75t_SL g1522 ( 
.A(n_1293),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1246),
.Y(n_1523)
);

XOR2xp5_ASAP7_75t_L g1524 ( 
.A(n_1211),
.B(n_1224),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1270),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1262),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1331),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1233),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1251),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1254),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1321),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1162),
.B(n_821),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1324),
.Y(n_1533)
);

NAND2xp33_ASAP7_75t_R g1534 ( 
.A(n_1179),
.B(n_707),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1287),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1296),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1303),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1347),
.B(n_710),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1359),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1329),
.Y(n_1540)
);

NAND2xp33_ASAP7_75t_SL g1541 ( 
.A(n_1234),
.B(n_1000),
.Y(n_1541)
);

BUFx2_ASAP7_75t_R g1542 ( 
.A(n_1200),
.Y(n_1542)
);

NOR2xp67_ASAP7_75t_L g1543 ( 
.A(n_1258),
.B(n_493),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1289),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1294),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1300),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1308),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1311),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1224),
.B(n_1024),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1318),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1248),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1250),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1252),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1232),
.B(n_1000),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1316),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1272),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1349),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1220),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1225),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1226),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1242),
.Y(n_1561)
);

XNOR2xp5_ASAP7_75t_L g1562 ( 
.A(n_1232),
.B(n_25),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1174),
.B(n_1335),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1174),
.B(n_1006),
.Y(n_1564)
);

AND2x6_ASAP7_75t_L g1565 ( 
.A(n_1290),
.B(n_760),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1243),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1283),
.Y(n_1567)
);

CKINVDCx20_ASAP7_75t_R g1568 ( 
.A(n_1244),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1335),
.B(n_1006),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1249),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1182),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1200),
.B(n_1006),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1184),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1327),
.B(n_1006),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1302),
.B(n_1007),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1312),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1277),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1315),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1304),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1317),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1319),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1320),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1322),
.Y(n_1583)
);

AND2x2_ASAP7_75t_SL g1584 ( 
.A(n_1328),
.B(n_1007),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1356),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1165),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1356),
.Y(n_1587)
);

INVx4_ASAP7_75t_SL g1588 ( 
.A(n_1219),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1279),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1356),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_R g1591 ( 
.A(n_1171),
.B(n_722),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1356),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1356),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1279),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1356),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1356),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1356),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1166),
.B(n_835),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1164),
.B(n_1007),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1356),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1356),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1356),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1356),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1356),
.B(n_729),
.Y(n_1604)
);

XOR2xp5_ASAP7_75t_L g1605 ( 
.A(n_1178),
.B(n_26),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1158),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1218),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1356),
.Y(n_1608)
);

INVxp33_ASAP7_75t_L g1609 ( 
.A(n_1338),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1164),
.B(n_1007),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1356),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1356),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1356),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1356),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1164),
.B(n_1039),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1279),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1279),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1279),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1356),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1356),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1356),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1260),
.B(n_840),
.Y(n_1622)
);

XOR2x2_ASAP7_75t_L g1623 ( 
.A(n_1204),
.B(n_27),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1165),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1260),
.B(n_861),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1356),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1356),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1356),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1356),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1260),
.B(n_897),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1356),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1218),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1356),
.B(n_752),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1356),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1356),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1356),
.B(n_753),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1356),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1164),
.B(n_1039),
.Y(n_1638)
);

XOR2x2_ASAP7_75t_L g1639 ( 
.A(n_1204),
.B(n_28),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1356),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1356),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1356),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1354),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1165),
.B(n_1039),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1356),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1356),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1164),
.B(n_1039),
.Y(n_1647)
);

XOR2xp5_ASAP7_75t_L g1648 ( 
.A(n_1178),
.B(n_28),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1606),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1362),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1379),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1443),
.B(n_762),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1644),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1585),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1369),
.B(n_29),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1367),
.B(n_904),
.Y(n_1656)
);

AND2x4_ASAP7_75t_SL g1657 ( 
.A(n_1644),
.B(n_913),
.Y(n_1657)
);

INVx3_ASAP7_75t_SL g1658 ( 
.A(n_1424),
.Y(n_1658)
);

OAI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1462),
.A2(n_1031),
.B(n_966),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1372),
.B(n_29),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1443),
.B(n_763),
.Y(n_1661)
);

NOR2xp33_ASAP7_75t_L g1662 ( 
.A(n_1455),
.B(n_1032),
.Y(n_1662)
);

AND2x2_ASAP7_75t_SL g1663 ( 
.A(n_1368),
.B(n_849),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1427),
.B(n_30),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1462),
.A2(n_1598),
.B(n_1484),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1375),
.B(n_30),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1379),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1587),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1563),
.B(n_31),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1433),
.B(n_32),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1408),
.B(n_773),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1405),
.B(n_32),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1590),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_L g1674 ( 
.A1(n_1387),
.A2(n_1036),
.B(n_695),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1366),
.B(n_1377),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1368),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1426),
.B(n_33),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1592),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1521),
.B(n_793),
.Y(n_1679)
);

BUFx6f_ASAP7_75t_L g1680 ( 
.A(n_1379),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1413),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1644),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1384),
.B(n_34),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1593),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1569),
.B(n_35),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1528),
.B(n_36),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1595),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1430),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1446),
.B(n_37),
.Y(n_1689)
);

BUFx6f_ASAP7_75t_L g1690 ( 
.A(n_1413),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1528),
.B(n_38),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1446),
.B(n_1588),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_R g1693 ( 
.A(n_1460),
.B(n_800),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1400),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1430),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1596),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1515),
.B(n_38),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1597),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1392),
.B(n_807),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1461),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1517),
.B(n_39),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1402),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1393),
.B(n_813),
.Y(n_1703)
);

INVxp67_ASAP7_75t_L g1704 ( 
.A(n_1383),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1382),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1394),
.B(n_815),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1600),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1601),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1406),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1407),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1446),
.B(n_39),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1524),
.B(n_1498),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1395),
.B(n_831),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1413),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1412),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1557),
.A2(n_975),
.B1(n_980),
.B2(n_972),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1396),
.B(n_1586),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1449),
.B(n_40),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1414),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1521),
.B(n_834),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1540),
.B(n_836),
.Y(n_1721)
);

BUFx3_ASAP7_75t_L g1722 ( 
.A(n_1418),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1370),
.B(n_1588),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1487),
.B(n_41),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1551),
.B(n_1552),
.Y(n_1725)
);

INVxp67_ASAP7_75t_SL g1726 ( 
.A(n_1643),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1428),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1553),
.B(n_42),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1602),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1603),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1436),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1504),
.B(n_42),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1643),
.Y(n_1733)
);

BUFx8_ASAP7_75t_L g1734 ( 
.A(n_1495),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1588),
.B(n_1036),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1514),
.B(n_43),
.Y(n_1736)
);

INVxp67_ASAP7_75t_SL g1737 ( 
.A(n_1440),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1444),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1398),
.B(n_844),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1509),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_SL g1741 ( 
.A(n_1471),
.B(n_695),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1451),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1415),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1438),
.B(n_43),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1608),
.Y(n_1745)
);

INVx4_ASAP7_75t_L g1746 ( 
.A(n_1495),
.Y(n_1746)
);

BUFx6f_ASAP7_75t_L g1747 ( 
.A(n_1451),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1544),
.B(n_1545),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1442),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1454),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1463),
.B(n_848),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1466),
.B(n_850),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1546),
.B(n_851),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1611),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1451),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1612),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1459),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1624),
.B(n_44),
.Y(n_1758)
);

BUFx4f_ASAP7_75t_L g1759 ( 
.A(n_1464),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1465),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1448),
.B(n_1364),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1609),
.B(n_45),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1447),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1613),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1547),
.B(n_856),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1526),
.B(n_46),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1481),
.B(n_860),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1389),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1391),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1419),
.B(n_46),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1378),
.B(n_47),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1598),
.A2(n_874),
.B(n_862),
.Y(n_1772)
);

BUFx4f_ASAP7_75t_L g1773 ( 
.A(n_1434),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1548),
.B(n_883),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1614),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1399),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1431),
.B(n_1519),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1619),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1431),
.B(n_47),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1525),
.B(n_1361),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1620),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1529),
.Y(n_1782)
);

BUFx6f_ASAP7_75t_L g1783 ( 
.A(n_1529),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1481),
.B(n_890),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1404),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1411),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1529),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1607),
.B(n_48),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1621),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1417),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1632),
.B(n_50),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1626),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1471),
.B(n_695),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1589),
.Y(n_1794)
);

INVx3_ASAP7_75t_L g1795 ( 
.A(n_1594),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1616),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1494),
.B(n_51),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1627),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1617),
.Y(n_1799)
);

AND2x2_ASAP7_75t_SL g1800 ( 
.A(n_1457),
.B(n_808),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1420),
.B(n_1421),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1401),
.B(n_892),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1401),
.B(n_906),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1390),
.B(n_51),
.Y(n_1804)
);

AND2x2_ASAP7_75t_SL g1805 ( 
.A(n_1423),
.B(n_52),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1387),
.A2(n_921),
.B(n_912),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1564),
.B(n_53),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1618),
.Y(n_1808)
);

INVx4_ASAP7_75t_L g1809 ( 
.A(n_1461),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1550),
.B(n_1416),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1380),
.B(n_934),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1381),
.B(n_947),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1549),
.B(n_1558),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1518),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1416),
.B(n_959),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1383),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1490),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1363),
.B(n_965),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1628),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1559),
.B(n_53),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1512),
.A2(n_988),
.B(n_969),
.Y(n_1821)
);

NAND2x1p5_ASAP7_75t_L g1822 ( 
.A(n_1425),
.B(n_54),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1560),
.B(n_55),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1561),
.B(n_56),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1573),
.B(n_997),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1566),
.B(n_56),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1429),
.B(n_57),
.Y(n_1827)
);

BUFx3_ASAP7_75t_L g1828 ( 
.A(n_1475),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1629),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1365),
.B(n_1002),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1570),
.B(n_57),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1432),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1516),
.B(n_58),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1500),
.B(n_695),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1489),
.B(n_1005),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1482),
.B(n_1435),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1554),
.B(n_59),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1523),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1478),
.B(n_1015),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1488),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1480),
.B(n_59),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1530),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1373),
.B(n_60),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1577),
.Y(n_1845)
);

BUFx3_ASAP7_75t_L g1846 ( 
.A(n_1475),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1631),
.Y(n_1847)
);

INVxp33_ASAP7_75t_L g1848 ( 
.A(n_1507),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1578),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1511),
.B(n_60),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1501),
.B(n_61),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1506),
.B(n_62),
.Y(n_1852)
);

BUFx6f_ASAP7_75t_L g1853 ( 
.A(n_1371),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1556),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1575),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1491),
.B(n_63),
.Y(n_1856)
);

BUFx6f_ASAP7_75t_L g1857 ( 
.A(n_1584),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1467),
.Y(n_1858)
);

INVx2_ASAP7_75t_SL g1859 ( 
.A(n_1599),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1374),
.Y(n_1860)
);

INVx4_ASAP7_75t_L g1861 ( 
.A(n_1439),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1562),
.Y(n_1862)
);

BUFx6f_ASAP7_75t_L g1863 ( 
.A(n_1439),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1610),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1445),
.B(n_1470),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1492),
.B(n_1493),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1497),
.B(n_1033),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1571),
.B(n_63),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1439),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1557),
.B(n_64),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1512),
.A2(n_1038),
.B(n_1037),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1496),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1469),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1634),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1499),
.B(n_1044),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1479),
.B(n_65),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1635),
.Y(n_1877)
);

INVx4_ASAP7_75t_L g1878 ( 
.A(n_1458),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1567),
.Y(n_1879)
);

AND2x2_ASAP7_75t_SL g1880 ( 
.A(n_1496),
.B(n_65),
.Y(n_1880)
);

NAND2x1p5_ASAP7_75t_L g1881 ( 
.A(n_1513),
.B(n_66),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1473),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1485),
.B(n_66),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1502),
.B(n_695),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1572),
.B(n_67),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1505),
.B(n_695),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1386),
.Y(n_1887)
);

BUFx3_ASAP7_75t_L g1888 ( 
.A(n_1388),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1615),
.B(n_68),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1483),
.B(n_68),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1637),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1638),
.B(n_69),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1640),
.Y(n_1893)
);

BUFx12f_ASAP7_75t_L g1894 ( 
.A(n_1555),
.Y(n_1894)
);

AND2x6_ASAP7_75t_L g1895 ( 
.A(n_1531),
.B(n_695),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1641),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1647),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1376),
.B(n_70),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1591),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1510),
.B(n_70),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1579),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1642),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1583),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1468),
.B(n_71),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1645),
.B(n_71),
.Y(n_1905)
);

NOR2xp33_ASAP7_75t_L g1906 ( 
.A(n_1646),
.B(n_72),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1580),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1533),
.B(n_73),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1472),
.B(n_73),
.Y(n_1909)
);

BUFx2_ASAP7_75t_L g1910 ( 
.A(n_1508),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1535),
.B(n_1536),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_R g1912 ( 
.A(n_1410),
.B(n_74),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1422),
.B(n_74),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1581),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1622),
.Y(n_1915)
);

INVx4_ASAP7_75t_L g1916 ( 
.A(n_1458),
.Y(n_1916)
);

INVx3_ASAP7_75t_L g1917 ( 
.A(n_1486),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1403),
.B(n_75),
.Y(n_1918)
);

INVx2_ASAP7_75t_SL g1919 ( 
.A(n_1537),
.Y(n_1919)
);

INVx4_ASAP7_75t_L g1920 ( 
.A(n_1458),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1582),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1622),
.Y(n_1922)
);

BUFx6f_ASAP7_75t_L g1923 ( 
.A(n_1567),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1520),
.B(n_75),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1625),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1625),
.Y(n_1926)
);

NOR2xp67_ASAP7_75t_L g1927 ( 
.A(n_1437),
.B(n_76),
.Y(n_1927)
);

BUFx3_ASAP7_75t_L g1928 ( 
.A(n_1574),
.Y(n_1928)
);

AND2x2_ASAP7_75t_SL g1929 ( 
.A(n_1542),
.B(n_76),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1630),
.B(n_77),
.Y(n_1930)
);

AND2x2_ASAP7_75t_SL g1931 ( 
.A(n_1542),
.B(n_77),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1630),
.B(n_78),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1532),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1474),
.B(n_78),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1604),
.B(n_79),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1532),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1576),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1500),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1539),
.Y(n_1939)
);

INVx2_ASAP7_75t_L g1940 ( 
.A(n_1567),
.Y(n_1940)
);

AND2x2_ASAP7_75t_L g1941 ( 
.A(n_1633),
.B(n_79),
.Y(n_1941)
);

INVx2_ASAP7_75t_SL g1942 ( 
.A(n_1503),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1450),
.B(n_80),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_1409),
.Y(n_1944)
);

INVx4_ASAP7_75t_L g1945 ( 
.A(n_1458),
.Y(n_1945)
);

BUFx3_ASAP7_75t_L g1946 ( 
.A(n_1565),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1527),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1636),
.B(n_80),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1565),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1522),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1441),
.Y(n_1951)
);

INVxp33_ASAP7_75t_L g1952 ( 
.A(n_1453),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1456),
.B(n_81),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1522),
.Y(n_1954)
);

OAI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1543),
.A2(n_490),
.B(n_489),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1538),
.B(n_81),
.Y(n_1956)
);

AND2x6_ASAP7_75t_L g1957 ( 
.A(n_1385),
.B(n_1522),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1565),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1541),
.B(n_83),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1543),
.Y(n_1960)
);

OAI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1385),
.A2(n_496),
.B(n_495),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1565),
.Y(n_1962)
);

INVx2_ASAP7_75t_R g1963 ( 
.A(n_1534),
.Y(n_1963)
);

AND2x6_ASAP7_75t_L g1964 ( 
.A(n_1452),
.B(n_500),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1623),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1568),
.B(n_84),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1639),
.B(n_85),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1397),
.B(n_86),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1605),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1648),
.B(n_87),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1400),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1606),
.B(n_88),
.Y(n_1972)
);

AND2x6_ASAP7_75t_L g1973 ( 
.A(n_1440),
.B(n_501),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1400),
.Y(n_1974)
);

NAND2x1p5_ASAP7_75t_L g1975 ( 
.A(n_1379),
.B(n_89),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1606),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1368),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1362),
.Y(n_1978)
);

AND2x4_ASAP7_75t_L g1979 ( 
.A(n_1446),
.B(n_89),
.Y(n_1979)
);

INVx2_ASAP7_75t_SL g1980 ( 
.A(n_1606),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1362),
.Y(n_1981)
);

INVx2_ASAP7_75t_SL g1982 ( 
.A(n_1606),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1400),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1606),
.B(n_90),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1368),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1606),
.B(n_90),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1443),
.B(n_91),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1400),
.Y(n_1988)
);

CKINVDCx5p33_ASAP7_75t_R g1989 ( 
.A(n_1424),
.Y(n_1989)
);

INVxp67_ASAP7_75t_SL g1990 ( 
.A(n_1368),
.Y(n_1990)
);

INVx2_ASAP7_75t_SL g1991 ( 
.A(n_1606),
.Y(n_1991)
);

INVxp67_ASAP7_75t_SL g1992 ( 
.A(n_1368),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1606),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1400),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1993),
.B(n_92),
.Y(n_1995)
);

OR2x6_ASAP7_75t_L g1996 ( 
.A(n_1746),
.B(n_92),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1937),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1915),
.B(n_93),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1947),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1651),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1922),
.B(n_1925),
.Y(n_2001)
);

BUFx6f_ASAP7_75t_SL g2002 ( 
.A(n_1746),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1947),
.Y(n_2003)
);

BUFx2_ASAP7_75t_L g2004 ( 
.A(n_1649),
.Y(n_2004)
);

BUFx6f_ASAP7_75t_L g2005 ( 
.A(n_1651),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1649),
.B(n_93),
.Y(n_2006)
);

INVx5_ASAP7_75t_L g2007 ( 
.A(n_1651),
.Y(n_2007)
);

NAND2x1p5_ASAP7_75t_L g2008 ( 
.A(n_1692),
.B(n_94),
.Y(n_2008)
);

INVx5_ASAP7_75t_L g2009 ( 
.A(n_1651),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1926),
.Y(n_2010)
);

AND2x4_ASAP7_75t_L g2011 ( 
.A(n_1954),
.B(n_95),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1801),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1780),
.B(n_95),
.Y(n_2013)
);

OR2x2_ASAP7_75t_L g2014 ( 
.A(n_1976),
.B(n_97),
.Y(n_2014)
);

BUFx2_ASAP7_75t_L g2015 ( 
.A(n_1980),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1933),
.B(n_97),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1667),
.Y(n_2017)
);

AND2x4_ASAP7_75t_L g2018 ( 
.A(n_1950),
.B(n_98),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1833),
.B(n_98),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1801),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1936),
.B(n_100),
.Y(n_2021)
);

INVx1_ASAP7_75t_SL g2022 ( 
.A(n_1982),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1748),
.B(n_1810),
.Y(n_2023)
);

AND2x4_ASAP7_75t_L g2024 ( 
.A(n_1950),
.B(n_100),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1937),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1801),
.Y(n_2026)
);

INVx4_ASAP7_75t_L g2027 ( 
.A(n_1667),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1991),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1748),
.B(n_101),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1675),
.B(n_102),
.Y(n_2030)
);

OR2x6_ASAP7_75t_L g2031 ( 
.A(n_1809),
.B(n_103),
.Y(n_2031)
);

AND2x4_ASAP7_75t_L g2032 ( 
.A(n_1939),
.B(n_103),
.Y(n_2032)
);

BUFx6f_ASAP7_75t_L g2033 ( 
.A(n_1667),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_L g2034 ( 
.A(n_1878),
.B(n_1916),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1694),
.Y(n_2035)
);

INVx2_ASAP7_75t_L g2036 ( 
.A(n_1814),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1777),
.B(n_105),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1694),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1712),
.B(n_106),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1911),
.B(n_109),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1702),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1814),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1702),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1828),
.B(n_111),
.Y(n_2044)
);

INVx3_ASAP7_75t_L g2045 ( 
.A(n_1667),
.Y(n_2045)
);

INVx3_ASAP7_75t_L g2046 ( 
.A(n_1680),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1709),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_1734),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1828),
.B(n_111),
.Y(n_2049)
);

AND2x4_ASAP7_75t_L g2050 ( 
.A(n_1846),
.B(n_112),
.Y(n_2050)
);

INVx3_ASAP7_75t_L g2051 ( 
.A(n_1680),
.Y(n_2051)
);

BUFx8_ASAP7_75t_L g2052 ( 
.A(n_1910),
.Y(n_2052)
);

NAND2x1p5_ASAP7_75t_L g2053 ( 
.A(n_1692),
.B(n_113),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1680),
.Y(n_2054)
);

NAND2x1p5_ASAP7_75t_L g2055 ( 
.A(n_1680),
.B(n_114),
.Y(n_2055)
);

INVx3_ASAP7_75t_L g2056 ( 
.A(n_1690),
.Y(n_2056)
);

NAND2x1p5_ASAP7_75t_L g2057 ( 
.A(n_1690),
.B(n_115),
.Y(n_2057)
);

NOR2xp67_ASAP7_75t_L g2058 ( 
.A(n_1704),
.B(n_503),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1833),
.B(n_115),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1804),
.B(n_1837),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1846),
.B(n_116),
.Y(n_2061)
);

AND2x4_ASAP7_75t_L g2062 ( 
.A(n_1911),
.B(n_116),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1788),
.B(n_117),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1709),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1710),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_1734),
.Y(n_2066)
);

NAND2x1_ASAP7_75t_SL g2067 ( 
.A(n_1658),
.B(n_117),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1710),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_1658),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_L g2070 ( 
.A(n_1690),
.B(n_504),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1715),
.Y(n_2071)
);

NAND2x1p5_ASAP7_75t_L g2072 ( 
.A(n_1690),
.B(n_118),
.Y(n_2072)
);

OR2x2_ASAP7_75t_L g2073 ( 
.A(n_1841),
.B(n_118),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1715),
.Y(n_2074)
);

BUFx6f_ASAP7_75t_L g2075 ( 
.A(n_1747),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1791),
.B(n_119),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1719),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1719),
.Y(n_2078)
);

BUFx3_ASAP7_75t_L g2079 ( 
.A(n_1989),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1743),
.Y(n_2080)
);

CKINVDCx8_ASAP7_75t_R g2081 ( 
.A(n_1989),
.Y(n_2081)
);

INVx1_ASAP7_75t_SL g2082 ( 
.A(n_1693),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1911),
.B(n_1813),
.Y(n_2083)
);

NOR2x1_ASAP7_75t_L g2084 ( 
.A(n_1878),
.B(n_119),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1693),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1743),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1971),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1725),
.B(n_120),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1971),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_1809),
.B(n_120),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1909),
.B(n_121),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1974),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1934),
.B(n_122),
.Y(n_2093)
);

OR2x6_ASAP7_75t_L g2094 ( 
.A(n_1689),
.B(n_122),
.Y(n_2094)
);

BUFx8_ASAP7_75t_L g2095 ( 
.A(n_1689),
.Y(n_2095)
);

BUFx2_ASAP7_75t_L g2096 ( 
.A(n_1912),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1912),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1704),
.B(n_123),
.Y(n_2098)
);

NOR2xp33_ASAP7_75t_L g2099 ( 
.A(n_1952),
.B(n_124),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_1723),
.B(n_125),
.Y(n_2100)
);

AND2x4_ASAP7_75t_L g2101 ( 
.A(n_1723),
.B(n_126),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1974),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1919),
.B(n_126),
.Y(n_2103)
);

INVx4_ASAP7_75t_L g2104 ( 
.A(n_1657),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1832),
.B(n_128),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_1723),
.B(n_128),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1832),
.B(n_129),
.Y(n_2107)
);

INVxp67_ASAP7_75t_SL g2108 ( 
.A(n_1688),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_1700),
.Y(n_2109)
);

NOR2xp67_ASAP7_75t_SL g2110 ( 
.A(n_1700),
.B(n_129),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_1977),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_SL g2112 ( 
.A(n_1816),
.B(n_130),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1983),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1732),
.B(n_1736),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1983),
.Y(n_2115)
);

AND2x6_ASAP7_75t_L g2116 ( 
.A(n_1770),
.B(n_130),
.Y(n_2116)
);

BUFx3_ASAP7_75t_L g2117 ( 
.A(n_1740),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1747),
.Y(n_2118)
);

BUFx12f_ASAP7_75t_L g2119 ( 
.A(n_1705),
.Y(n_2119)
);

NOR2xp67_ASAP7_75t_L g2120 ( 
.A(n_1816),
.B(n_508),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1988),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_1917),
.B(n_131),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_1977),
.Y(n_2123)
);

OR2x6_ASAP7_75t_L g2124 ( 
.A(n_1711),
.B(n_1979),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_1917),
.B(n_131),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1988),
.Y(n_2126)
);

OR2x6_ASAP7_75t_L g2127 ( 
.A(n_1711),
.B(n_132),
.Y(n_2127)
);

AND2x4_ASAP7_75t_L g2128 ( 
.A(n_1726),
.B(n_133),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1994),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1994),
.Y(n_2130)
);

INVx3_ASAP7_75t_L g2131 ( 
.A(n_1681),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1747),
.Y(n_2132)
);

BUFx6f_ASAP7_75t_L g2133 ( 
.A(n_1747),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1669),
.B(n_133),
.Y(n_2134)
);

BUFx2_ASAP7_75t_L g2135 ( 
.A(n_1985),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_1862),
.B(n_134),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_1726),
.B(n_135),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_1985),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1873),
.Y(n_2139)
);

BUFx3_ASAP7_75t_L g2140 ( 
.A(n_1740),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1851),
.B(n_136),
.Y(n_2141)
);

NAND2x1p5_ASAP7_75t_L g2142 ( 
.A(n_1759),
.B(n_136),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_1852),
.B(n_137),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1738),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_1916),
.B(n_137),
.Y(n_2145)
);

BUFx12f_ASAP7_75t_L g2146 ( 
.A(n_1717),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1759),
.Y(n_2147)
);

AND2x4_ASAP7_75t_L g2148 ( 
.A(n_1920),
.B(n_138),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1660),
.B(n_1744),
.Y(n_2149)
);

BUFx2_ASAP7_75t_L g2150 ( 
.A(n_1990),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1738),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1856),
.B(n_138),
.Y(n_2152)
);

INVx4_ASAP7_75t_L g2153 ( 
.A(n_1657),
.Y(n_2153)
);

AND2x6_ASAP7_75t_L g2154 ( 
.A(n_1770),
.B(n_139),
.Y(n_2154)
);

NOR2x1_ASAP7_75t_L g2155 ( 
.A(n_1920),
.B(n_139),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_1862),
.B(n_140),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1873),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1945),
.B(n_140),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_SL g2159 ( 
.A(n_1945),
.B(n_512),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1972),
.B(n_141),
.Y(n_2160)
);

AND2x2_ASAP7_75t_L g2161 ( 
.A(n_1984),
.B(n_141),
.Y(n_2161)
);

AND2x4_ASAP7_75t_L g2162 ( 
.A(n_1733),
.B(n_142),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1721),
.B(n_142),
.Y(n_2163)
);

BUFx12f_ASAP7_75t_L g2164 ( 
.A(n_1929),
.Y(n_2164)
);

OR2x6_ASAP7_75t_L g2165 ( 
.A(n_1979),
.B(n_144),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_1986),
.B(n_144),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1721),
.B(n_1753),
.Y(n_2167)
);

INVx2_ASAP7_75t_SL g2168 ( 
.A(n_1771),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1655),
.B(n_145),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_1733),
.B(n_146),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1763),
.Y(n_2171)
);

BUFx6f_ASAP7_75t_L g2172 ( 
.A(n_1783),
.Y(n_2172)
);

BUFx12f_ASAP7_75t_L g2173 ( 
.A(n_1929),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1722),
.B(n_147),
.Y(n_2174)
);

NAND2x1p5_ASAP7_75t_L g2175 ( 
.A(n_1681),
.B(n_147),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1763),
.Y(n_2176)
);

BUFx6f_ASAP7_75t_L g2177 ( 
.A(n_1783),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_SL g2178 ( 
.A(n_1931),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1882),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1845),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1845),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_1753),
.B(n_148),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1849),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1765),
.B(n_150),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1849),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_1882),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_1924),
.B(n_1967),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_1722),
.B(n_150),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_1783),
.Y(n_2189)
);

AND2x6_ASAP7_75t_L g2190 ( 
.A(n_1770),
.B(n_152),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1765),
.B(n_152),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1860),
.Y(n_2192)
);

INVx3_ASAP7_75t_L g2193 ( 
.A(n_1863),
.Y(n_2193)
);

BUFx6f_ASAP7_75t_L g2194 ( 
.A(n_1783),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_1965),
.B(n_1865),
.Y(n_2195)
);

BUFx4f_ASAP7_75t_L g2196 ( 
.A(n_1805),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_1952),
.B(n_153),
.Y(n_2197)
);

CKINVDCx8_ASAP7_75t_R g2198 ( 
.A(n_1967),
.Y(n_2198)
);

INVx5_ASAP7_75t_L g2199 ( 
.A(n_1863),
.Y(n_2199)
);

BUFx12f_ASAP7_75t_L g2200 ( 
.A(n_1931),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1768),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_1894),
.B(n_153),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_1990),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_1761),
.B(n_154),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_1727),
.B(n_155),
.Y(n_2205)
);

OR2x6_ASAP7_75t_L g2206 ( 
.A(n_1771),
.B(n_155),
.Y(n_2206)
);

AND2x4_ASAP7_75t_L g2207 ( 
.A(n_1727),
.B(n_156),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_L g2208 ( 
.A(n_1894),
.B(n_156),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1774),
.B(n_157),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1774),
.B(n_157),
.Y(n_2210)
);

NOR2xp33_ASAP7_75t_L g2211 ( 
.A(n_1825),
.B(n_158),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_1677),
.Y(n_2212)
);

INVx2_ASAP7_75t_SL g2213 ( 
.A(n_1714),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1860),
.Y(n_2214)
);

BUFx4f_ASAP7_75t_L g2215 ( 
.A(n_1805),
.Y(n_2215)
);

BUFx6f_ASAP7_75t_L g2216 ( 
.A(n_1787),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1768),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1663),
.B(n_158),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1825),
.B(n_1872),
.Y(n_2219)
);

INVx2_ASAP7_75t_SL g2220 ( 
.A(n_1714),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1769),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_1769),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_1992),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_1872),
.B(n_159),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_L g2225 ( 
.A(n_1800),
.B(n_159),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_1731),
.B(n_160),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1737),
.Y(n_2227)
);

CKINVDCx20_ASAP7_75t_R g2228 ( 
.A(n_1899),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1666),
.B(n_160),
.Y(n_2229)
);

OR2x6_ASAP7_75t_L g2230 ( 
.A(n_1975),
.B(n_161),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1672),
.B(n_161),
.Y(n_2231)
);

BUFx6f_ASAP7_75t_L g2232 ( 
.A(n_1787),
.Y(n_2232)
);

AND2x4_ASAP7_75t_L g2233 ( 
.A(n_1731),
.B(n_162),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_1992),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1737),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1664),
.B(n_162),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_SL g2237 ( 
.A(n_1663),
.B(n_518),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_1776),
.Y(n_2238)
);

BUFx12f_ASAP7_75t_L g2239 ( 
.A(n_1899),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1776),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1749),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1749),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1966),
.B(n_163),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_1800),
.B(n_164),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1683),
.B(n_1670),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_1868),
.B(n_165),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1750),
.Y(n_2247)
);

INVxp67_ASAP7_75t_SL g2248 ( 
.A(n_1688),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_1863),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_SL g2250 ( 
.A(n_1880),
.B(n_166),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_1848),
.B(n_168),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_1850),
.B(n_168),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_1785),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_1695),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_1785),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1750),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1786),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1757),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_1942),
.B(n_169),
.Y(n_2259)
);

OAI21x1_ASAP7_75t_L g2260 ( 
.A1(n_1674),
.A2(n_521),
.B(n_519),
.Y(n_2260)
);

OR2x6_ASAP7_75t_L g2261 ( 
.A(n_1975),
.B(n_170),
.Y(n_2261)
);

CKINVDCx6p67_ASAP7_75t_R g2262 ( 
.A(n_1908),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_1888),
.B(n_170),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_1762),
.B(n_1842),
.Y(n_2264)
);

OR2x2_ASAP7_75t_L g2265 ( 
.A(n_1758),
.B(n_171),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_1695),
.Y(n_2266)
);

BUFx12f_ASAP7_75t_L g2267 ( 
.A(n_1944),
.Y(n_2267)
);

BUFx2_ASAP7_75t_L g2268 ( 
.A(n_1827),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1757),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1848),
.B(n_171),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1728),
.B(n_172),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_1888),
.B(n_172),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1779),
.B(n_173),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1650),
.B(n_173),
.Y(n_2274)
);

OR2x6_ASAP7_75t_L g2275 ( 
.A(n_1908),
.B(n_174),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1786),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_1790),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1790),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1794),
.Y(n_2279)
);

INVx4_ASAP7_75t_L g2280 ( 
.A(n_1863),
.Y(n_2280)
);

HB1xp67_ASAP7_75t_L g2281 ( 
.A(n_1827),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1760),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1686),
.B(n_174),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_1880),
.B(n_175),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1691),
.B(n_175),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_1671),
.B(n_176),
.Y(n_2286)
);

BUFx6f_ASAP7_75t_L g2287 ( 
.A(n_1787),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_1654),
.B(n_176),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1760),
.Y(n_2289)
);

BUFx6f_ASAP7_75t_L g2290 ( 
.A(n_1787),
.Y(n_2290)
);

BUFx2_ASAP7_75t_L g2291 ( 
.A(n_1827),
.Y(n_2291)
);

BUFx12f_ASAP7_75t_L g2292 ( 
.A(n_1944),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_SL g2293 ( 
.A(n_1951),
.B(n_177),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1854),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_SL g2295 ( 
.A(n_1973),
.B(n_523),
.Y(n_2295)
);

INVx3_ASAP7_75t_L g2296 ( 
.A(n_1861),
.Y(n_2296)
);

BUFx6f_ASAP7_75t_L g2297 ( 
.A(n_1879),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_SL g2298 ( 
.A(n_1951),
.B(n_177),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_SL g2299 ( 
.A(n_1973),
.B(n_524),
.Y(n_2299)
);

AND2x2_ASAP7_75t_L g2300 ( 
.A(n_1908),
.B(n_178),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1794),
.Y(n_2301)
);

OR2x2_ASAP7_75t_L g2302 ( 
.A(n_1818),
.B(n_178),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_1854),
.Y(n_2303)
);

HB1xp67_ASAP7_75t_L g2304 ( 
.A(n_1653),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_1682),
.B(n_179),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_1879),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_1879),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1796),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_1830),
.B(n_179),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1817),
.Y(n_2310)
);

INVx1_ASAP7_75t_SL g2311 ( 
.A(n_1797),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_SL g2312 ( 
.A(n_1676),
.B(n_180),
.Y(n_2312)
);

AND2x6_ASAP7_75t_L g2313 ( 
.A(n_1844),
.B(n_180),
.Y(n_2313)
);

INVxp67_ASAP7_75t_L g2314 ( 
.A(n_1890),
.Y(n_2314)
);

CKINVDCx5p33_ASAP7_75t_R g2315 ( 
.A(n_1913),
.Y(n_2315)
);

AND2x2_ASAP7_75t_L g2316 ( 
.A(n_1685),
.B(n_181),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_SL g2317 ( 
.A(n_1973),
.B(n_525),
.Y(n_2317)
);

OR2x2_ASAP7_75t_L g2318 ( 
.A(n_1969),
.B(n_181),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1817),
.Y(n_2319)
);

INVx5_ASAP7_75t_L g2320 ( 
.A(n_1973),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_1834),
.B(n_182),
.Y(n_2321)
);

INVx8_ASAP7_75t_L g2322 ( 
.A(n_1890),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1839),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_1879),
.Y(n_2324)
);

BUFx3_ASAP7_75t_L g2325 ( 
.A(n_1735),
.Y(n_2325)
);

AND2x6_ASAP7_75t_L g2326 ( 
.A(n_1844),
.B(n_183),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_1676),
.Y(n_2327)
);

CKINVDCx11_ASAP7_75t_R g2328 ( 
.A(n_1735),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_1697),
.B(n_184),
.Y(n_2329)
);

INVx5_ASAP7_75t_L g2330 ( 
.A(n_1973),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_SL g2331 ( 
.A(n_1964),
.B(n_184),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_1864),
.B(n_185),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1766),
.B(n_185),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1839),
.Y(n_2334)
);

INVx4_ASAP7_75t_L g2335 ( 
.A(n_1861),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1796),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_1811),
.B(n_186),
.Y(n_2337)
);

NOR2xp33_ASAP7_75t_SL g2338 ( 
.A(n_1964),
.B(n_186),
.Y(n_2338)
);

BUFx12f_ASAP7_75t_L g2339 ( 
.A(n_1881),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_1701),
.B(n_187),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_1869),
.Y(n_2341)
);

HB1xp67_ASAP7_75t_L g2342 ( 
.A(n_1844),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1870),
.B(n_187),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_1970),
.B(n_189),
.Y(n_2344)
);

BUFx6f_ASAP7_75t_L g2345 ( 
.A(n_1923),
.Y(n_2345)
);

AND2x4_ASAP7_75t_L g2346 ( 
.A(n_1668),
.B(n_189),
.Y(n_2346)
);

INVx4_ASAP7_75t_L g2347 ( 
.A(n_1869),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_1857),
.B(n_190),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_1843),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_1843),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_1808),
.Y(n_2351)
);

BUFx6f_ASAP7_75t_L g2352 ( 
.A(n_1923),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1679),
.B(n_190),
.Y(n_2353)
);

OR2x6_ASAP7_75t_L g2354 ( 
.A(n_1881),
.B(n_191),
.Y(n_2354)
);

INVx3_ASAP7_75t_L g2355 ( 
.A(n_1923),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1679),
.B(n_1720),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_1811),
.B(n_191),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_1923),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_1808),
.Y(n_2359)
);

AND2x4_ASAP7_75t_L g2360 ( 
.A(n_1673),
.B(n_192),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_1678),
.B(n_1684),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_1720),
.B(n_193),
.Y(n_2362)
);

NAND2x1p5_ASAP7_75t_L g2363 ( 
.A(n_1773),
.B(n_193),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1718),
.B(n_194),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1927),
.B(n_194),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_1806),
.B(n_195),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_1866),
.Y(n_2367)
);

NAND2x1p5_ASAP7_75t_L g2368 ( 
.A(n_1773),
.B(n_195),
.Y(n_2368)
);

CKINVDCx8_ASAP7_75t_R g2369 ( 
.A(n_1957),
.Y(n_2369)
);

BUFx6f_ASAP7_75t_L g2370 ( 
.A(n_1755),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1907),
.Y(n_2371)
);

INVx1_ASAP7_75t_SL g2372 ( 
.A(n_1735),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_1857),
.Y(n_2373)
);

HB1xp67_ASAP7_75t_L g2374 ( 
.A(n_1822),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_1887),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_1755),
.Y(n_2376)
);

CKINVDCx20_ASAP7_75t_R g2377 ( 
.A(n_1968),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1907),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_1858),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1724),
.B(n_196),
.Y(n_2380)
);

NOR2x1_ASAP7_75t_L g2381 ( 
.A(n_1946),
.B(n_196),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_1887),
.Y(n_2382)
);

AND2x4_ASAP7_75t_L g2383 ( 
.A(n_1687),
.B(n_197),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_1812),
.B(n_197),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_SL g2385 ( 
.A(n_1964),
.B(n_526),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_1812),
.B(n_1772),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_1696),
.B(n_198),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_1914),
.Y(n_2388)
);

BUFx4f_ASAP7_75t_L g2389 ( 
.A(n_1822),
.Y(n_2389)
);

BUFx3_ASAP7_75t_L g2390 ( 
.A(n_1928),
.Y(n_2390)
);

BUFx12f_ASAP7_75t_L g2391 ( 
.A(n_1957),
.Y(n_2391)
);

AND2x4_ASAP7_75t_L g2392 ( 
.A(n_1698),
.B(n_198),
.Y(n_2392)
);

BUFx12f_ASAP7_75t_L g2393 ( 
.A(n_1957),
.Y(n_2393)
);

BUFx6f_ASAP7_75t_L g2394 ( 
.A(n_1946),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_1656),
.B(n_199),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1914),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_1921),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_1820),
.B(n_200),
.Y(n_2398)
);

BUFx6f_ASAP7_75t_L g2399 ( 
.A(n_1742),
.Y(n_2399)
);

NAND2x1p5_ASAP7_75t_L g2400 ( 
.A(n_1858),
.B(n_200),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_1921),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1656),
.B(n_201),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1884),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_1742),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_1901),
.Y(n_2405)
);

BUFx2_ASAP7_75t_SL g2406 ( 
.A(n_1964),
.Y(n_2406)
);

AND2x6_ASAP7_75t_L g2407 ( 
.A(n_1857),
.B(n_201),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1886),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_1901),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1900),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_1840),
.B(n_202),
.Y(n_2411)
);

INVx3_ASAP7_75t_L g2412 ( 
.A(n_1928),
.Y(n_2412)
);

NAND2x1_ASAP7_75t_SL g2413 ( 
.A(n_1959),
.B(n_202),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1903),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_1903),
.Y(n_2415)
);

AND2x2_ASAP7_75t_SL g2416 ( 
.A(n_1857),
.B(n_203),
.Y(n_2416)
);

OR2x6_ASAP7_75t_L g2417 ( 
.A(n_1959),
.B(n_203),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_1707),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_1823),
.B(n_206),
.Y(n_2419)
);

NAND2x1_ASAP7_75t_SL g2420 ( 
.A(n_1716),
.B(n_206),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_1708),
.Y(n_2421)
);

BUFx5_ASAP7_75t_L g2422 ( 
.A(n_1895),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_1656),
.B(n_207),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1662),
.B(n_208),
.Y(n_2424)
);

INVx3_ASAP7_75t_L g2425 ( 
.A(n_1795),
.Y(n_2425)
);

BUFx3_ASAP7_75t_L g2426 ( 
.A(n_1824),
.Y(n_2426)
);

NAND2x1p5_ASAP7_75t_L g2427 ( 
.A(n_1859),
.B(n_208),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_1729),
.B(n_209),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1662),
.B(n_209),
.Y(n_2429)
);

AND2x4_ASAP7_75t_L g2430 ( 
.A(n_1730),
.B(n_211),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_1826),
.B(n_212),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_1745),
.B(n_212),
.Y(n_2432)
);

INVx4_ASAP7_75t_L g2433 ( 
.A(n_1964),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_1897),
.B(n_1831),
.Y(n_2434)
);

BUFx6f_ASAP7_75t_L g2435 ( 
.A(n_1782),
.Y(n_2435)
);

INVx4_ASAP7_75t_L g2436 ( 
.A(n_1782),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_1754),
.Y(n_2437)
);

AND2x2_ASAP7_75t_L g2438 ( 
.A(n_1840),
.B(n_213),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_1930),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_1756),
.Y(n_2440)
);

AND2x4_ASAP7_75t_L g2441 ( 
.A(n_1764),
.B(n_215),
.Y(n_2441)
);

HB1xp67_ASAP7_75t_L g2442 ( 
.A(n_1889),
.Y(n_2442)
);

OR2x2_ASAP7_75t_L g2443 ( 
.A(n_1775),
.B(n_216),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1906),
.B(n_216),
.Y(n_2444)
);

HB1xp67_ASAP7_75t_L g2445 ( 
.A(n_1892),
.Y(n_2445)
);

CKINVDCx5p33_ASAP7_75t_R g2446 ( 
.A(n_1963),
.Y(n_2446)
);

INVx3_ASAP7_75t_L g2447 ( 
.A(n_1795),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_1778),
.B(n_217),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_1932),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_1906),
.B(n_217),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1905),
.B(n_218),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_1781),
.Y(n_2452)
);

BUFx2_ASAP7_75t_L g2453 ( 
.A(n_1838),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1789),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_1807),
.B(n_219),
.Y(n_2455)
);

AND2x4_ASAP7_75t_L g2456 ( 
.A(n_1792),
.B(n_219),
.Y(n_2456)
);

AND2x4_ASAP7_75t_L g2457 ( 
.A(n_1798),
.B(n_220),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_SL g2458 ( 
.A(n_1652),
.B(n_221),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_1940),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1819),
.B(n_222),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_1829),
.Y(n_2461)
);

OR2x6_ASAP7_75t_L g2462 ( 
.A(n_1904),
.B(n_1898),
.Y(n_2462)
);

NAND2x1p5_ASAP7_75t_L g2463 ( 
.A(n_1799),
.B(n_223),
.Y(n_2463)
);

BUFx12f_ASAP7_75t_L g2464 ( 
.A(n_1957),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1847),
.B(n_223),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_1874),
.B(n_224),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_1877),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_1891),
.Y(n_2468)
);

OR2x2_ASAP7_75t_L g2469 ( 
.A(n_1893),
.B(n_224),
.Y(n_2469)
);

INVxp67_ASAP7_75t_SL g2470 ( 
.A(n_1885),
.Y(n_2470)
);

NAND2x1p5_ASAP7_75t_L g2471 ( 
.A(n_1799),
.B(n_225),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2361),
.Y(n_2472)
);

AND2x2_ASAP7_75t_SL g2473 ( 
.A(n_2196),
.B(n_1958),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2146),
.Y(n_2474)
);

INVx4_ASAP7_75t_L g2475 ( 
.A(n_2124),
.Y(n_2475)
);

INVx5_ASAP7_75t_L g2476 ( 
.A(n_2407),
.Y(n_2476)
);

AOI22xp33_ASAP7_75t_L g2477 ( 
.A1(n_2196),
.A2(n_1963),
.B1(n_1941),
.B2(n_1948),
.Y(n_2477)
);

BUFx8_ASAP7_75t_L g2478 ( 
.A(n_2002),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2023),
.B(n_1665),
.Y(n_2479)
);

BUFx3_ASAP7_75t_L g2480 ( 
.A(n_2048),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_2000),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2010),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2000),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2010),
.Y(n_2484)
);

BUFx6f_ASAP7_75t_L g2485 ( 
.A(n_2000),
.Y(n_2485)
);

INVx4_ASAP7_75t_L g2486 ( 
.A(n_2124),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2452),
.Y(n_2487)
);

INVx5_ASAP7_75t_L g2488 ( 
.A(n_2407),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2452),
.Y(n_2489)
);

BUFx12f_ASAP7_75t_L g2490 ( 
.A(n_2066),
.Y(n_2490)
);

BUFx3_ASAP7_75t_L g2491 ( 
.A(n_2069),
.Y(n_2491)
);

INVx1_ASAP7_75t_SL g2492 ( 
.A(n_2022),
.Y(n_2492)
);

CKINVDCx5p33_ASAP7_75t_R g2493 ( 
.A(n_2052),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2180),
.Y(n_2494)
);

BUFx12f_ASAP7_75t_L g2495 ( 
.A(n_2052),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2119),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2454),
.Y(n_2497)
);

BUFx4f_ASAP7_75t_SL g2498 ( 
.A(n_2095),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2454),
.Y(n_2499)
);

INVx3_ASAP7_75t_L g2500 ( 
.A(n_2369),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2467),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_2095),
.Y(n_2502)
);

OR2x6_ASAP7_75t_L g2503 ( 
.A(n_2322),
.B(n_1896),
.Y(n_2503)
);

INVx1_ASAP7_75t_SL g2504 ( 
.A(n_2150),
.Y(n_2504)
);

NAND2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2104),
.B(n_1958),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2367),
.B(n_1938),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_2367),
.B(n_1938),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2180),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2181),
.Y(n_2509)
);

HB1xp67_ASAP7_75t_L g2510 ( 
.A(n_2203),
.Y(n_2510)
);

NAND2x1p5_ASAP7_75t_L g2511 ( 
.A(n_2104),
.B(n_1940),
.Y(n_2511)
);

BUFx6f_ASAP7_75t_L g2512 ( 
.A(n_2005),
.Y(n_2512)
);

INVx3_ASAP7_75t_L g2513 ( 
.A(n_2373),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2181),
.Y(n_2514)
);

INVx5_ASAP7_75t_L g2515 ( 
.A(n_2407),
.Y(n_2515)
);

BUFx6f_ASAP7_75t_L g2516 ( 
.A(n_2005),
.Y(n_2516)
);

BUFx2_ASAP7_75t_L g2517 ( 
.A(n_2153),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2153),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2183),
.Y(n_2519)
);

BUFx3_ASAP7_75t_L g2520 ( 
.A(n_2081),
.Y(n_2520)
);

CKINVDCx5p33_ASAP7_75t_R g2521 ( 
.A(n_2267),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_2339),
.Y(n_2522)
);

CKINVDCx11_ASAP7_75t_R g2523 ( 
.A(n_2292),
.Y(n_2523)
);

INVx6_ASAP7_75t_L g2524 ( 
.A(n_2117),
.Y(n_2524)
);

INVx2_ASAP7_75t_L g2525 ( 
.A(n_2183),
.Y(n_2525)
);

BUFx8_ASAP7_75t_L g2526 ( 
.A(n_2002),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2467),
.Y(n_2527)
);

NOR2xp67_ASAP7_75t_SL g2528 ( 
.A(n_2320),
.B(n_1661),
.Y(n_2528)
);

INVx4_ASAP7_75t_L g2529 ( 
.A(n_2094),
.Y(n_2529)
);

CKINVDCx16_ASAP7_75t_R g2530 ( 
.A(n_1996),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2185),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2185),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_2079),
.Y(n_2533)
);

BUFx2_ASAP7_75t_L g2534 ( 
.A(n_2004),
.Y(n_2534)
);

BUFx6f_ASAP7_75t_L g2535 ( 
.A(n_2005),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2418),
.Y(n_2536)
);

INVx5_ASAP7_75t_L g2537 ( 
.A(n_2407),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2421),
.Y(n_2538)
);

INVx5_ASAP7_75t_L g2539 ( 
.A(n_2094),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2001),
.B(n_1659),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2035),
.Y(n_2541)
);

BUFx12f_ASAP7_75t_L g2542 ( 
.A(n_1996),
.Y(n_2542)
);

CKINVDCx5p33_ASAP7_75t_R g2543 ( 
.A(n_2239),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_2373),
.Y(n_2544)
);

CKINVDCx16_ASAP7_75t_R g2545 ( 
.A(n_2031),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2437),
.Y(n_2546)
);

BUFx2_ASAP7_75t_L g2547 ( 
.A(n_2015),
.Y(n_2547)
);

INVxp67_ASAP7_75t_SL g2548 ( 
.A(n_2281),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2322),
.Y(n_2549)
);

INVxp67_ASAP7_75t_SL g2550 ( 
.A(n_2342),
.Y(n_2550)
);

BUFx3_ASAP7_75t_L g2551 ( 
.A(n_2140),
.Y(n_2551)
);

BUFx3_ASAP7_75t_L g2552 ( 
.A(n_2147),
.Y(n_2552)
);

BUFx12f_ASAP7_75t_L g2553 ( 
.A(n_2031),
.Y(n_2553)
);

BUFx10_ASAP7_75t_L g2554 ( 
.A(n_2090),
.Y(n_2554)
);

BUFx2_ASAP7_75t_L g2555 ( 
.A(n_2127),
.Y(n_2555)
);

BUFx2_ASAP7_75t_SL g2556 ( 
.A(n_2044),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2335),
.Y(n_2557)
);

BUFx6f_ASAP7_75t_L g2558 ( 
.A(n_2017),
.Y(n_2558)
);

CKINVDCx11_ASAP7_75t_R g2559 ( 
.A(n_2082),
.Y(n_2559)
);

INVx3_ASAP7_75t_L g2560 ( 
.A(n_2335),
.Y(n_2560)
);

INVx6_ASAP7_75t_L g2561 ( 
.A(n_2347),
.Y(n_2561)
);

AOI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_2250),
.A2(n_1957),
.B1(n_1876),
.B2(n_1883),
.Y(n_2562)
);

INVx2_ASAP7_75t_SL g2563 ( 
.A(n_2028),
.Y(n_2563)
);

AND2x2_ASAP7_75t_L g2564 ( 
.A(n_2060),
.B(n_1902),
.Y(n_2564)
);

BUFx12f_ASAP7_75t_L g2565 ( 
.A(n_2090),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2127),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2440),
.Y(n_2567)
);

BUFx6f_ASAP7_75t_L g2568 ( 
.A(n_2017),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2461),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2468),
.Y(n_2570)
);

INVxp67_ASAP7_75t_SL g2571 ( 
.A(n_2263),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2035),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1999),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2187),
.B(n_1978),
.Y(n_2574)
);

BUFx3_ASAP7_75t_L g2575 ( 
.A(n_2109),
.Y(n_2575)
);

INVx2_ASAP7_75t_SL g2576 ( 
.A(n_2044),
.Y(n_2576)
);

INVx1_ASAP7_75t_SL g2577 ( 
.A(n_2223),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2038),
.Y(n_2578)
);

INVx1_ASAP7_75t_SL g2579 ( 
.A(n_2234),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2039),
.B(n_1981),
.Y(n_2580)
);

INVx4_ASAP7_75t_L g2581 ( 
.A(n_2165),
.Y(n_2581)
);

INVx5_ASAP7_75t_L g2582 ( 
.A(n_2165),
.Y(n_2582)
);

INVx4_ASAP7_75t_L g2583 ( 
.A(n_2275),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2123),
.Y(n_2584)
);

BUFx12f_ASAP7_75t_L g2585 ( 
.A(n_2328),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2017),
.Y(n_2586)
);

NOR2xp33_ASAP7_75t_L g2587 ( 
.A(n_2167),
.B(n_1767),
.Y(n_2587)
);

BUFx24_ASAP7_75t_L g2588 ( 
.A(n_2049),
.Y(n_2588)
);

INVx3_ASAP7_75t_L g2589 ( 
.A(n_2347),
.Y(n_2589)
);

INVx5_ASAP7_75t_L g2590 ( 
.A(n_2116),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_1999),
.Y(n_2591)
);

OR2x6_ASAP7_75t_L g2592 ( 
.A(n_2275),
.B(n_1987),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2038),
.Y(n_2593)
);

AOI22xp33_ASAP7_75t_L g2594 ( 
.A1(n_2215),
.A2(n_1935),
.B1(n_1943),
.B2(n_1918),
.Y(n_2594)
);

BUFx3_ASAP7_75t_L g2595 ( 
.A(n_2085),
.Y(n_2595)
);

INVx6_ASAP7_75t_SL g2596 ( 
.A(n_2354),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2007),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2262),
.Y(n_2598)
);

INVx8_ASAP7_75t_L g2599 ( 
.A(n_2354),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_2389),
.B(n_1961),
.Y(n_2600)
);

INVx1_ASAP7_75t_SL g2601 ( 
.A(n_2135),
.Y(n_2601)
);

INVx5_ASAP7_75t_L g2602 ( 
.A(n_2116),
.Y(n_2602)
);

BUFx2_ASAP7_75t_L g2603 ( 
.A(n_2116),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2041),
.Y(n_2604)
);

BUFx3_ASAP7_75t_L g2605 ( 
.A(n_2390),
.Y(n_2605)
);

INVx5_ASAP7_75t_SL g2606 ( 
.A(n_2230),
.Y(n_2606)
);

INVx3_ASAP7_75t_L g2607 ( 
.A(n_2007),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2041),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2007),
.Y(n_2609)
);

CKINVDCx20_ASAP7_75t_R g2610 ( 
.A(n_2228),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2047),
.Y(n_2611)
);

BUFx12f_ASAP7_75t_L g2612 ( 
.A(n_2164),
.Y(n_2612)
);

INVx1_ASAP7_75t_SL g2613 ( 
.A(n_2138),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2003),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2003),
.Y(n_2615)
);

BUFx8_ASAP7_75t_L g2616 ( 
.A(n_2178),
.Y(n_2616)
);

BUFx2_ASAP7_75t_L g2617 ( 
.A(n_2116),
.Y(n_2617)
);

AND2x6_ASAP7_75t_L g2618 ( 
.A(n_2145),
.B(n_1949),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2049),
.Y(n_2619)
);

BUFx2_ASAP7_75t_L g2620 ( 
.A(n_2154),
.Y(n_2620)
);

BUFx3_ASAP7_75t_L g2621 ( 
.A(n_2050),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2047),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2068),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2068),
.Y(n_2624)
);

CKINVDCx6p67_ASAP7_75t_R g2625 ( 
.A(n_2178),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2215),
.B(n_2206),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2443),
.Y(n_2627)
);

OAI21xp33_ASAP7_75t_L g2628 ( 
.A1(n_2356),
.A2(n_1953),
.B(n_1871),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2050),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2033),
.Y(n_2630)
);

INVxp67_ASAP7_75t_SL g2631 ( 
.A(n_2263),
.Y(n_2631)
);

INVx6_ASAP7_75t_L g2632 ( 
.A(n_2391),
.Y(n_2632)
);

BUFx3_ASAP7_75t_L g2633 ( 
.A(n_2061),
.Y(n_2633)
);

INVx3_ASAP7_75t_L g2634 ( 
.A(n_2009),
.Y(n_2634)
);

CKINVDCx16_ASAP7_75t_R g2635 ( 
.A(n_2293),
.Y(n_2635)
);

HB1xp67_ASAP7_75t_L g2636 ( 
.A(n_2266),
.Y(n_2636)
);

OR2x6_ASAP7_75t_L g2637 ( 
.A(n_2206),
.B(n_1855),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2074),
.Y(n_2638)
);

INVx3_ASAP7_75t_L g2639 ( 
.A(n_2009),
.Y(n_2639)
);

INVx5_ASAP7_75t_SL g2640 ( 
.A(n_2230),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2448),
.Y(n_2641)
);

BUFx2_ASAP7_75t_L g2642 ( 
.A(n_2154),
.Y(n_2642)
);

HB1xp67_ASAP7_75t_L g2643 ( 
.A(n_2254),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2469),
.Y(n_2644)
);

BUFx4f_ASAP7_75t_SL g2645 ( 
.A(n_2393),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2327),
.Y(n_2646)
);

INVx4_ASAP7_75t_L g2647 ( 
.A(n_2009),
.Y(n_2647)
);

INVxp67_ASAP7_75t_SL g2648 ( 
.A(n_2272),
.Y(n_2648)
);

INVx1_ASAP7_75t_SL g2649 ( 
.A(n_2272),
.Y(n_2649)
);

INVxp67_ASAP7_75t_SL g2650 ( 
.A(n_2108),
.Y(n_2650)
);

INVx3_ASAP7_75t_L g2651 ( 
.A(n_2464),
.Y(n_2651)
);

INVx1_ASAP7_75t_SL g2652 ( 
.A(n_2174),
.Y(n_2652)
);

INVx5_ASAP7_75t_L g2653 ( 
.A(n_2154),
.Y(n_2653)
);

BUFx3_ASAP7_75t_L g2654 ( 
.A(n_2061),
.Y(n_2654)
);

INVx1_ASAP7_75t_SL g2655 ( 
.A(n_2174),
.Y(n_2655)
);

BUFx12f_ASAP7_75t_L g2656 ( 
.A(n_2173),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2074),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2032),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2439),
.B(n_1821),
.Y(n_2659)
);

BUFx12f_ASAP7_75t_L g2660 ( 
.A(n_2200),
.Y(n_2660)
);

OR2x2_ASAP7_75t_L g2661 ( 
.A(n_2195),
.B(n_1836),
.Y(n_2661)
);

BUFx3_ASAP7_75t_L g2662 ( 
.A(n_2188),
.Y(n_2662)
);

INVx8_ASAP7_75t_L g2663 ( 
.A(n_2154),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2032),
.Y(n_2664)
);

INVx5_ASAP7_75t_L g2665 ( 
.A(n_2190),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2439),
.B(n_1867),
.Y(n_2666)
);

BUFx3_ASAP7_75t_L g2667 ( 
.A(n_2188),
.Y(n_2667)
);

INVx4_ASAP7_75t_L g2668 ( 
.A(n_2190),
.Y(n_2668)
);

BUFx3_ASAP7_75t_L g2669 ( 
.A(n_2205),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2033),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2274),
.Y(n_2671)
);

AOI22xp5_ASAP7_75t_L g2672 ( 
.A1(n_2190),
.A2(n_1895),
.B1(n_1956),
.B2(n_1875),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2274),
.Y(n_2673)
);

OAI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_2237),
.A2(n_1815),
.B1(n_1855),
.B2(n_1784),
.Y(n_2674)
);

BUFx6f_ASAP7_75t_L g2675 ( 
.A(n_2033),
.Y(n_2675)
);

INVx5_ASAP7_75t_L g2676 ( 
.A(n_2190),
.Y(n_2676)
);

BUFx3_ASAP7_75t_L g2677 ( 
.A(n_2205),
.Y(n_2677)
);

BUFx5_ASAP7_75t_L g2678 ( 
.A(n_2077),
.Y(n_2678)
);

INVx2_ASAP7_75t_SL g2679 ( 
.A(n_2207),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2288),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_2449),
.B(n_1895),
.Y(n_2681)
);

NOR2xp67_ASAP7_75t_L g2682 ( 
.A(n_2320),
.B(n_1962),
.Y(n_2682)
);

NAND2x1p5_ASAP7_75t_L g2683 ( 
.A(n_2320),
.B(n_1949),
.Y(n_2683)
);

INVx3_ASAP7_75t_SL g2684 ( 
.A(n_2315),
.Y(n_2684)
);

INVx6_ASAP7_75t_SL g2685 ( 
.A(n_2261),
.Y(n_2685)
);

INVx2_ASAP7_75t_SL g2686 ( 
.A(n_2207),
.Y(n_2686)
);

OR2x6_ASAP7_75t_L g2687 ( 
.A(n_2018),
.B(n_1699),
.Y(n_2687)
);

AND2x4_ASAP7_75t_L g2688 ( 
.A(n_2330),
.B(n_1703),
.Y(n_2688)
);

BUFx2_ASAP7_75t_SL g2689 ( 
.A(n_2313),
.Y(n_2689)
);

INVx1_ASAP7_75t_SL g2690 ( 
.A(n_2233),
.Y(n_2690)
);

INVx4_ASAP7_75t_L g2691 ( 
.A(n_2313),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_2417),
.A2(n_1895),
.B1(n_1793),
.B2(n_1835),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2288),
.Y(n_2693)
);

BUFx3_ASAP7_75t_L g2694 ( 
.A(n_2233),
.Y(n_2694)
);

INVx6_ASAP7_75t_L g2695 ( 
.A(n_2100),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_SL g2696 ( 
.A1(n_2313),
.A2(n_1895),
.B1(n_1955),
.B2(n_1853),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2449),
.B(n_1706),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2346),
.Y(n_2698)
);

CKINVDCx14_ASAP7_75t_R g2699 ( 
.A(n_2377),
.Y(n_2699)
);

INVx1_ASAP7_75t_SL g2700 ( 
.A(n_2111),
.Y(n_2700)
);

BUFx2_ASAP7_75t_L g2701 ( 
.A(n_2313),
.Y(n_2701)
);

INVx4_ASAP7_75t_L g2702 ( 
.A(n_2326),
.Y(n_2702)
);

AO21x2_ASAP7_75t_L g2703 ( 
.A1(n_2058),
.A2(n_1793),
.B(n_1741),
.Y(n_2703)
);

BUFx8_ASAP7_75t_L g2704 ( 
.A(n_2096),
.Y(n_2704)
);

BUFx3_ASAP7_75t_L g2705 ( 
.A(n_2100),
.Y(n_2705)
);

INVx5_ASAP7_75t_SL g2706 ( 
.A(n_2261),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2417),
.A2(n_1835),
.B1(n_1741),
.B2(n_1960),
.Y(n_2707)
);

OR2x2_ASAP7_75t_L g2708 ( 
.A(n_1995),
.B(n_1713),
.Y(n_2708)
);

INVx4_ASAP7_75t_L g2709 ( 
.A(n_2326),
.Y(n_2709)
);

CKINVDCx16_ASAP7_75t_R g2710 ( 
.A(n_2298),
.Y(n_2710)
);

BUFx3_ASAP7_75t_L g2711 ( 
.A(n_2101),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_2101),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2346),
.Y(n_2713)
);

OR2x2_ASAP7_75t_L g2714 ( 
.A(n_2344),
.B(n_1739),
.Y(n_2714)
);

BUFx2_ASAP7_75t_SL g2715 ( 
.A(n_2326),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2077),
.Y(n_2716)
);

BUFx4_ASAP7_75t_SL g2717 ( 
.A(n_2325),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2078),
.Y(n_2718)
);

INVx1_ASAP7_75t_SL g2719 ( 
.A(n_2372),
.Y(n_2719)
);

BUFx3_ASAP7_75t_L g2720 ( 
.A(n_2106),
.Y(n_2720)
);

BUFx2_ASAP7_75t_L g2721 ( 
.A(n_2326),
.Y(n_2721)
);

BUFx3_ASAP7_75t_L g2722 ( 
.A(n_2106),
.Y(n_2722)
);

INVx3_ASAP7_75t_SL g2723 ( 
.A(n_2018),
.Y(n_2723)
);

BUFx2_ASAP7_75t_SL g2724 ( 
.A(n_2024),
.Y(n_2724)
);

BUFx3_ASAP7_75t_L g2725 ( 
.A(n_2198),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2078),
.Y(n_2726)
);

AOI22xp33_ASAP7_75t_L g2727 ( 
.A1(n_2209),
.A2(n_1803),
.B1(n_1802),
.B2(n_1752),
.Y(n_2727)
);

INVx8_ASAP7_75t_L g2728 ( 
.A(n_2199),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2024),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2141),
.B(n_1751),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2389),
.Y(n_2731)
);

BUFx4_ASAP7_75t_SL g2732 ( 
.A(n_2097),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2075),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_SL g2734 ( 
.A(n_2237),
.B(n_1853),
.Y(n_2734)
);

INVx4_ASAP7_75t_L g2735 ( 
.A(n_2199),
.Y(n_2735)
);

INVx6_ASAP7_75t_L g2736 ( 
.A(n_2199),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2083),
.B(n_1853),
.Y(n_2737)
);

BUFx6f_ASAP7_75t_L g2738 ( 
.A(n_2075),
.Y(n_2738)
);

BUFx3_ASAP7_75t_L g2739 ( 
.A(n_2008),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2122),
.Y(n_2740)
);

INVx5_ASAP7_75t_SL g2741 ( 
.A(n_2416),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2360),
.Y(n_2742)
);

AOI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2219),
.A2(n_1853),
.B1(n_228),
.B2(n_225),
.Y(n_2743)
);

INVx6_ASAP7_75t_L g2744 ( 
.A(n_2062),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2360),
.Y(n_2745)
);

BUFx2_ASAP7_75t_SL g2746 ( 
.A(n_2330),
.Y(n_2746)
);

CKINVDCx20_ASAP7_75t_R g2747 ( 
.A(n_2073),
.Y(n_2747)
);

CKINVDCx20_ASAP7_75t_R g2748 ( 
.A(n_2136),
.Y(n_2748)
);

BUFx2_ASAP7_75t_SL g2749 ( 
.A(n_2330),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2410),
.B(n_226),
.Y(n_2750)
);

INVx2_ASAP7_75t_SL g2751 ( 
.A(n_2053),
.Y(n_2751)
);

INVx1_ASAP7_75t_SL g2752 ( 
.A(n_2122),
.Y(n_2752)
);

INVx5_ASAP7_75t_L g2753 ( 
.A(n_2027),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2383),
.Y(n_2754)
);

AOI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2470),
.A2(n_230),
.B1(n_226),
.B2(n_229),
.Y(n_2755)
);

BUFx3_ASAP7_75t_L g2756 ( 
.A(n_2296),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2075),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_2374),
.Y(n_2758)
);

BUFx12f_ASAP7_75t_L g2759 ( 
.A(n_2142),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_SL g2760 ( 
.A(n_2312),
.B(n_229),
.Y(n_2760)
);

NAND2x1p5_ASAP7_75t_L g2761 ( 
.A(n_2268),
.B(n_231),
.Y(n_2761)
);

INVx6_ASAP7_75t_L g2762 ( 
.A(n_2062),
.Y(n_2762)
);

BUFx3_ASAP7_75t_L g2763 ( 
.A(n_2296),
.Y(n_2763)
);

CKINVDCx5p33_ASAP7_75t_R g2764 ( 
.A(n_2156),
.Y(n_2764)
);

AND2x2_ASAP7_75t_L g2765 ( 
.A(n_2143),
.B(n_2152),
.Y(n_2765)
);

INVx4_ASAP7_75t_L g2766 ( 
.A(n_2145),
.Y(n_2766)
);

BUFx6f_ASAP7_75t_L g2767 ( 
.A(n_2118),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2118),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2383),
.Y(n_2769)
);

BUFx12f_ASAP7_75t_L g2770 ( 
.A(n_2363),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2027),
.Y(n_2771)
);

BUFx4_ASAP7_75t_SL g2772 ( 
.A(n_2087),
.Y(n_2772)
);

BUFx3_ASAP7_75t_L g2773 ( 
.A(n_2341),
.Y(n_2773)
);

INVx1_ASAP7_75t_SL g2774 ( 
.A(n_2125),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2386),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.Y(n_2775)
);

CKINVDCx6p67_ASAP7_75t_R g2776 ( 
.A(n_2162),
.Y(n_2776)
);

INVx2_ASAP7_75t_SL g2777 ( 
.A(n_2162),
.Y(n_2777)
);

BUFx2_ASAP7_75t_L g2778 ( 
.A(n_2128),
.Y(n_2778)
);

INVxp67_ASAP7_75t_SL g2779 ( 
.A(n_2248),
.Y(n_2779)
);

INVx3_ASAP7_75t_L g2780 ( 
.A(n_2148),
.Y(n_2780)
);

AOI22xp5_ASAP7_75t_L g2781 ( 
.A1(n_2291),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.Y(n_2781)
);

BUFx12f_ASAP7_75t_L g2782 ( 
.A(n_2368),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2387),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2087),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2295),
.B(n_236),
.Y(n_2785)
);

BUFx4f_ASAP7_75t_SL g2786 ( 
.A(n_2148),
.Y(n_2786)
);

BUFx4f_ASAP7_75t_SL g2787 ( 
.A(n_2158),
.Y(n_2787)
);

NAND2x1p5_ASAP7_75t_L g2788 ( 
.A(n_2158),
.B(n_237),
.Y(n_2788)
);

INVx5_ASAP7_75t_L g2789 ( 
.A(n_2370),
.Y(n_2789)
);

AND2x4_ASAP7_75t_L g2790 ( 
.A(n_2012),
.B(n_237),
.Y(n_2790)
);

BUFx3_ASAP7_75t_L g2791 ( 
.A(n_2341),
.Y(n_2791)
);

NAND2x1p5_ASAP7_75t_L g2792 ( 
.A(n_2125),
.B(n_239),
.Y(n_2792)
);

INVx1_ASAP7_75t_SL g2793 ( 
.A(n_2226),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2410),
.B(n_239),
.Y(n_2794)
);

BUFx3_ASAP7_75t_L g2795 ( 
.A(n_2170),
.Y(n_2795)
);

INVx4_ASAP7_75t_L g2796 ( 
.A(n_2370),
.Y(n_2796)
);

INVx2_ASAP7_75t_SL g2797 ( 
.A(n_2170),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2089),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2089),
.Y(n_2799)
);

INVx2_ASAP7_75t_SL g2800 ( 
.A(n_2387),
.Y(n_2800)
);

INVx2_ASAP7_75t_SL g2801 ( 
.A(n_2392),
.Y(n_2801)
);

BUFx6f_ASAP7_75t_L g2802 ( 
.A(n_2118),
.Y(n_2802)
);

AND2x4_ASAP7_75t_L g2803 ( 
.A(n_2012),
.B(n_240),
.Y(n_2803)
);

AND2x4_ASAP7_75t_L g2804 ( 
.A(n_2020),
.B(n_241),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_2102),
.Y(n_2805)
);

BUFx3_ASAP7_75t_L g2806 ( 
.A(n_2427),
.Y(n_2806)
);

INVx5_ASAP7_75t_SL g2807 ( 
.A(n_2128),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2102),
.Y(n_2808)
);

BUFx2_ASAP7_75t_SL g2809 ( 
.A(n_2392),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2403),
.B(n_242),
.Y(n_2810)
);

NAND2x1p5_ASAP7_75t_L g2811 ( 
.A(n_2137),
.B(n_243),
.Y(n_2811)
);

INVxp67_ASAP7_75t_SL g2812 ( 
.A(n_2295),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_2280),
.Y(n_2813)
);

BUFx12f_ASAP7_75t_L g2814 ( 
.A(n_2305),
.Y(n_2814)
);

INVx3_ASAP7_75t_L g2815 ( 
.A(n_2280),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2428),
.Y(n_2816)
);

BUFx12f_ASAP7_75t_L g2817 ( 
.A(n_2428),
.Y(n_2817)
);

BUFx12f_ASAP7_75t_L g2818 ( 
.A(n_2430),
.Y(n_2818)
);

NAND2x1p5_ASAP7_75t_L g2819 ( 
.A(n_2137),
.B(n_244),
.Y(n_2819)
);

INVx3_ASAP7_75t_L g2820 ( 
.A(n_2121),
.Y(n_2820)
);

BUFx3_ASAP7_75t_L g2821 ( 
.A(n_2121),
.Y(n_2821)
);

BUFx6f_ASAP7_75t_L g2822 ( 
.A(n_2132),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2430),
.Y(n_2823)
);

OAI22xp5_ASAP7_75t_L g2824 ( 
.A1(n_2453),
.A2(n_248),
.B1(n_244),
.B2(n_246),
.Y(n_2824)
);

BUFx6f_ASAP7_75t_L g2825 ( 
.A(n_2132),
.Y(n_2825)
);

INVx5_ASAP7_75t_L g2826 ( 
.A(n_2370),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2432),
.Y(n_2827)
);

BUFx4f_ASAP7_75t_SL g2828 ( 
.A(n_2412),
.Y(n_2828)
);

INVxp67_ASAP7_75t_SL g2829 ( 
.A(n_2299),
.Y(n_2829)
);

CKINVDCx20_ASAP7_75t_R g2830 ( 
.A(n_2014),
.Y(n_2830)
);

INVx3_ASAP7_75t_SL g2831 ( 
.A(n_2432),
.Y(n_2831)
);

BUFx3_ASAP7_75t_L g2832 ( 
.A(n_2129),
.Y(n_2832)
);

CKINVDCx14_ASAP7_75t_R g2833 ( 
.A(n_2202),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2129),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2130),
.Y(n_2835)
);

BUFx2_ASAP7_75t_SL g2836 ( 
.A(n_2441),
.Y(n_2836)
);

BUFx3_ASAP7_75t_L g2837 ( 
.A(n_2130),
.Y(n_2837)
);

BUFx4_ASAP7_75t_SL g2838 ( 
.A(n_2294),
.Y(n_2838)
);

INVx5_ASAP7_75t_L g2839 ( 
.A(n_2376),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2441),
.Y(n_2840)
);

INVx2_ASAP7_75t_L g2841 ( 
.A(n_2294),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2456),
.Y(n_2842)
);

CKINVDCx5p33_ASAP7_75t_R g2843 ( 
.A(n_2208),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2456),
.Y(n_2844)
);

AOI22xp33_ASAP7_75t_L g2845 ( 
.A1(n_2211),
.A2(n_250),
.B1(n_246),
.B2(n_249),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2303),
.Y(n_2846)
);

BUFx2_ASAP7_75t_L g2847 ( 
.A(n_2400),
.Y(n_2847)
);

INVx5_ASAP7_75t_L g2848 ( 
.A(n_2376),
.Y(n_2848)
);

BUFx12f_ASAP7_75t_L g2849 ( 
.A(n_2457),
.Y(n_2849)
);

BUFx2_ASAP7_75t_SL g2850 ( 
.A(n_2457),
.Y(n_2850)
);

BUFx8_ASAP7_75t_SL g2851 ( 
.A(n_2446),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2144),
.Y(n_2852)
);

INVx3_ASAP7_75t_L g2853 ( 
.A(n_2303),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2144),
.Y(n_2854)
);

AOI22xp33_ASAP7_75t_L g2855 ( 
.A1(n_2218),
.A2(n_252),
.B1(n_249),
.B2(n_251),
.Y(n_2855)
);

BUFx4f_ASAP7_75t_SL g2856 ( 
.A(n_2412),
.Y(n_2856)
);

INVx3_ASAP7_75t_L g2857 ( 
.A(n_2371),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2151),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2463),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2741),
.A2(n_2244),
.B1(n_2225),
.B2(n_2284),
.Y(n_2860)
);

AOI22xp33_ASAP7_75t_L g2861 ( 
.A1(n_2741),
.A2(n_2337),
.B1(n_2411),
.B2(n_2357),
.Y(n_2861)
);

AOI22xp33_ASAP7_75t_L g2862 ( 
.A1(n_2741),
.A2(n_2251),
.B1(n_2426),
.B2(n_2099),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_SL g2863 ( 
.A1(n_2786),
.A2(n_2338),
.B1(n_2331),
.B2(n_2299),
.Y(n_2863)
);

OAI22xp5_ASAP7_75t_L g2864 ( 
.A1(n_2786),
.A2(n_2462),
.B1(n_2300),
.B2(n_2149),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2495),
.Y(n_2865)
);

OAI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2787),
.A2(n_2462),
.B1(n_2114),
.B2(n_2314),
.Y(n_2866)
);

BUFx6f_ASAP7_75t_L g2867 ( 
.A(n_2728),
.Y(n_2867)
);

INVx6_ASAP7_75t_L g2868 ( 
.A(n_2478),
.Y(n_2868)
);

CKINVDCx20_ASAP7_75t_R g2869 ( 
.A(n_2498),
.Y(n_2869)
);

INVx6_ASAP7_75t_L g2870 ( 
.A(n_2478),
.Y(n_2870)
);

INVx2_ASAP7_75t_L g2871 ( 
.A(n_2494),
.Y(n_2871)
);

OAI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2787),
.A2(n_2442),
.B1(n_2445),
.B2(n_2245),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2508),
.Y(n_2873)
);

AOI22xp33_ASAP7_75t_SL g2874 ( 
.A1(n_2599),
.A2(n_2317),
.B1(n_2385),
.B2(n_2406),
.Y(n_2874)
);

NAND2x1p5_ASAP7_75t_L g2875 ( 
.A(n_2539),
.B(n_2110),
.Y(n_2875)
);

BUFx3_ASAP7_75t_L g2876 ( 
.A(n_2498),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2472),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2564),
.B(n_2013),
.Y(n_2878)
);

INVx2_ASAP7_75t_L g2879 ( 
.A(n_2509),
.Y(n_2879)
);

INVx1_ASAP7_75t_SL g2880 ( 
.A(n_2772),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2514),
.Y(n_2881)
);

AOI22xp33_ASAP7_75t_L g2882 ( 
.A1(n_2599),
.A2(n_2197),
.B1(n_2264),
.B2(n_2134),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2661),
.B(n_2587),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2519),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2525),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2571),
.A2(n_2168),
.B1(n_2471),
.B2(n_2011),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_SL g2887 ( 
.A1(n_2599),
.A2(n_2724),
.B1(n_2606),
.B2(n_2706),
.Y(n_2887)
);

INVx3_ASAP7_75t_SL g2888 ( 
.A(n_2493),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2536),
.Y(n_2889)
);

BUFx3_ASAP7_75t_L g2890 ( 
.A(n_2526),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2538),
.Y(n_2891)
);

INVx2_ASAP7_75t_SL g2892 ( 
.A(n_2772),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2546),
.Y(n_2893)
);

INVx8_ASAP7_75t_L g2894 ( 
.A(n_2728),
.Y(n_2894)
);

BUFx4f_ASAP7_75t_SL g2895 ( 
.A(n_2490),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2567),
.Y(n_2896)
);

OAI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_2530),
.A2(n_2317),
.B1(n_2385),
.B2(n_2159),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2531),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2526),
.Y(n_2899)
);

BUFx2_ASAP7_75t_L g2900 ( 
.A(n_2596),
.Y(n_2900)
);

BUFx12f_ASAP7_75t_L g2901 ( 
.A(n_2523),
.Y(n_2901)
);

INVx6_ASAP7_75t_L g2902 ( 
.A(n_2728),
.Y(n_2902)
);

CKINVDCx20_ASAP7_75t_R g2903 ( 
.A(n_2610),
.Y(n_2903)
);

OAI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2571),
.A2(n_2011),
.B1(n_2259),
.B2(n_2311),
.Y(n_2904)
);

AOI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2587),
.A2(n_2182),
.B1(n_2184),
.B2(n_2163),
.Y(n_2905)
);

INVxp67_ASAP7_75t_L g2906 ( 
.A(n_2534),
.Y(n_2906)
);

INVx1_ASAP7_75t_L g2907 ( 
.A(n_2569),
.Y(n_2907)
);

OAI22xp5_ASAP7_75t_L g2908 ( 
.A1(n_2631),
.A2(n_2259),
.B1(n_2316),
.B2(n_2455),
.Y(n_2908)
);

BUFx2_ASAP7_75t_L g2909 ( 
.A(n_2596),
.Y(n_2909)
);

INVx6_ASAP7_75t_L g2910 ( 
.A(n_2585),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2570),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2487),
.Y(n_2912)
);

INVx3_ASAP7_75t_SL g2913 ( 
.A(n_2521),
.Y(n_2913)
);

INVx3_ASAP7_75t_L g2914 ( 
.A(n_2663),
.Y(n_2914)
);

BUFx2_ASAP7_75t_R g2915 ( 
.A(n_2480),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2631),
.A2(n_2433),
.B1(n_2265),
.B2(n_2235),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2489),
.Y(n_2917)
);

CKINVDCx6p67_ASAP7_75t_R g2918 ( 
.A(n_2588),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2497),
.Y(n_2919)
);

BUFx2_ASAP7_75t_L g2920 ( 
.A(n_2685),
.Y(n_2920)
);

CKINVDCx5p33_ASAP7_75t_R g2921 ( 
.A(n_2838),
.Y(n_2921)
);

AND2x2_ASAP7_75t_L g2922 ( 
.A(n_2574),
.B(n_2063),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2499),
.Y(n_2923)
);

AOI22xp33_ASAP7_75t_SL g2924 ( 
.A1(n_2606),
.A2(n_2159),
.B1(n_2433),
.B2(n_2366),
.Y(n_2924)
);

CKINVDCx12_ASAP7_75t_R g2925 ( 
.A(n_2838),
.Y(n_2925)
);

NAND2x1p5_ASAP7_75t_L g2926 ( 
.A(n_2539),
.B(n_2084),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2501),
.Y(n_2927)
);

AOI22xp33_ASAP7_75t_L g2928 ( 
.A1(n_2583),
.A2(n_2210),
.B1(n_2191),
.B2(n_2243),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2527),
.Y(n_2929)
);

INVx6_ASAP7_75t_L g2930 ( 
.A(n_2616),
.Y(n_2930)
);

AND2x4_ASAP7_75t_L g2931 ( 
.A(n_2668),
.B(n_2371),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2650),
.Y(n_2932)
);

INVx6_ASAP7_75t_L g2933 ( 
.A(n_2616),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2648),
.A2(n_2227),
.B1(n_2235),
.B2(n_2076),
.Y(n_2934)
);

INVx2_ASAP7_75t_SL g2935 ( 
.A(n_2522),
.Y(n_2935)
);

AOI22xp33_ASAP7_75t_SL g2936 ( 
.A1(n_2606),
.A2(n_2019),
.B1(n_2059),
.B2(n_2091),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2650),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2779),
.Y(n_2938)
);

INVx4_ASAP7_75t_L g2939 ( 
.A(n_2663),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_SL g2940 ( 
.A1(n_2640),
.A2(n_2093),
.B1(n_2175),
.B2(n_2384),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2779),
.Y(n_2941)
);

INVx1_ASAP7_75t_L g2942 ( 
.A(n_2852),
.Y(n_2942)
);

AOI22xp33_ASAP7_75t_SL g2943 ( 
.A1(n_2640),
.A2(n_2438),
.B1(n_2246),
.B2(n_2227),
.Y(n_2943)
);

CKINVDCx20_ASAP7_75t_R g2944 ( 
.A(n_2699),
.Y(n_2944)
);

INVx1_ASAP7_75t_SL g2945 ( 
.A(n_2684),
.Y(n_2945)
);

OAI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2545),
.A2(n_2318),
.B1(n_2332),
.B2(n_2212),
.Y(n_2946)
);

INVx2_ASAP7_75t_L g2947 ( 
.A(n_2532),
.Y(n_2947)
);

INVx6_ASAP7_75t_L g2948 ( 
.A(n_2704),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2541),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2572),
.Y(n_2950)
);

BUFx6f_ASAP7_75t_SL g2951 ( 
.A(n_2554),
.Y(n_2951)
);

AOI22xp33_ASAP7_75t_L g2952 ( 
.A1(n_2583),
.A2(n_2030),
.B1(n_2362),
.B2(n_2353),
.Y(n_2952)
);

INVx2_ASAP7_75t_L g2953 ( 
.A(n_2578),
.Y(n_2953)
);

BUFx2_ASAP7_75t_L g2954 ( 
.A(n_2685),
.Y(n_2954)
);

AOI22xp33_ASAP7_75t_L g2955 ( 
.A1(n_2640),
.A2(n_2458),
.B1(n_2029),
.B2(n_2340),
.Y(n_2955)
);

BUFx3_ASAP7_75t_L g2956 ( 
.A(n_2496),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2593),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2706),
.A2(n_2329),
.B1(n_2419),
.B2(n_2398),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_SL g2959 ( 
.A1(n_2706),
.A2(n_2422),
.B1(n_2055),
.B2(n_2072),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2854),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2529),
.A2(n_2431),
.B1(n_2169),
.B2(n_2429),
.Y(n_2961)
);

AOI22xp33_ASAP7_75t_L g2962 ( 
.A1(n_2529),
.A2(n_2424),
.B1(n_2365),
.B2(n_2273),
.Y(n_2962)
);

AOI21xp33_ASAP7_75t_L g2963 ( 
.A1(n_2628),
.A2(n_2252),
.B(n_2321),
.Y(n_2963)
);

CKINVDCx14_ASAP7_75t_R g2964 ( 
.A(n_2474),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2604),
.Y(n_2965)
);

BUFx6f_ASAP7_75t_L g2966 ( 
.A(n_2481),
.Y(n_2966)
);

AOI22xp33_ASAP7_75t_L g2967 ( 
.A1(n_2581),
.A2(n_2161),
.B1(n_2166),
.B2(n_2160),
.Y(n_2967)
);

OAI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2648),
.A2(n_2364),
.B1(n_2380),
.B2(n_2378),
.Y(n_2968)
);

HB1xp67_ASAP7_75t_L g2969 ( 
.A(n_2504),
.Y(n_2969)
);

BUFx4f_ASAP7_75t_SL g2970 ( 
.A(n_2759),
.Y(n_2970)
);

OAI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2807),
.A2(n_2378),
.B1(n_2396),
.B2(n_2388),
.Y(n_2971)
);

BUFx3_ASAP7_75t_L g2972 ( 
.A(n_2575),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2805),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2608),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_2581),
.A2(n_2105),
.B1(n_2107),
.B2(n_2444),
.Y(n_2975)
);

OAI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2807),
.A2(n_2388),
.B1(n_2397),
.B2(n_2396),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2805),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2611),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2573),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2591),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2622),
.Y(n_2981)
);

CKINVDCx20_ASAP7_75t_R g2982 ( 
.A(n_2559),
.Y(n_2982)
);

CKINVDCx11_ASAP7_75t_R g2983 ( 
.A(n_2542),
.Y(n_2983)
);

AOI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_2539),
.A2(n_2450),
.B1(n_2270),
.B2(n_2006),
.Y(n_2984)
);

BUFx6f_ASAP7_75t_L g2985 ( 
.A(n_2481),
.Y(n_2985)
);

CKINVDCx11_ASAP7_75t_R g2986 ( 
.A(n_2553),
.Y(n_2986)
);

CKINVDCx20_ASAP7_75t_R g2987 ( 
.A(n_2520),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2666),
.B(n_2151),
.Y(n_2988)
);

BUFx6f_ASAP7_75t_L g2989 ( 
.A(n_2481),
.Y(n_2989)
);

BUFx10_ASAP7_75t_L g2990 ( 
.A(n_2502),
.Y(n_2990)
);

BUFx4f_ASAP7_75t_SL g2991 ( 
.A(n_2565),
.Y(n_2991)
);

INVx3_ASAP7_75t_L g2992 ( 
.A(n_2663),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2765),
.B(n_2643),
.Y(n_2993)
);

BUFx3_ASAP7_75t_L g2994 ( 
.A(n_2533),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2623),
.Y(n_2995)
);

CKINVDCx11_ASAP7_75t_R g2996 ( 
.A(n_2612),
.Y(n_2996)
);

BUFx12f_ASAP7_75t_L g2997 ( 
.A(n_2554),
.Y(n_2997)
);

BUFx2_ASAP7_75t_L g2998 ( 
.A(n_2503),
.Y(n_2998)
);

BUFx4f_ASAP7_75t_SL g2999 ( 
.A(n_2814),
.Y(n_2999)
);

CKINVDCx11_ASAP7_75t_R g3000 ( 
.A(n_2656),
.Y(n_3000)
);

INVx5_ASAP7_75t_L g3001 ( 
.A(n_2503),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2624),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2483),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2858),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2646),
.Y(n_3005)
);

AOI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2748),
.A2(n_2040),
.B1(n_2434),
.B2(n_2285),
.Y(n_3006)
);

AOI22xp33_ASAP7_75t_L g3007 ( 
.A1(n_2582),
.A2(n_2204),
.B1(n_2098),
.B2(n_2112),
.Y(n_3007)
);

BUFx3_ASAP7_75t_L g3008 ( 
.A(n_2551),
.Y(n_3008)
);

INVx6_ASAP7_75t_L g3009 ( 
.A(n_2704),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2582),
.A2(n_2809),
.B1(n_2850),
.B2(n_2836),
.Y(n_3010)
);

AOI22xp33_ASAP7_75t_L g3011 ( 
.A1(n_2582),
.A2(n_2309),
.B1(n_2302),
.B2(n_2286),
.Y(n_3011)
);

INVx1_ASAP7_75t_L g3012 ( 
.A(n_2482),
.Y(n_3012)
);

INVx1_ASAP7_75t_SL g3013 ( 
.A(n_2492),
.Y(n_3013)
);

AOI22xp33_ASAP7_75t_L g3014 ( 
.A1(n_2637),
.A2(n_2395),
.B1(n_2423),
.B2(n_2402),
.Y(n_3014)
);

AOI22xp33_ASAP7_75t_SL g3015 ( 
.A1(n_2556),
.A2(n_2422),
.B1(n_2057),
.B2(n_2176),
.Y(n_3015)
);

AOI22xp33_ASAP7_75t_L g3016 ( 
.A1(n_2637),
.A2(n_2037),
.B1(n_2021),
.B2(n_2016),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2484),
.Y(n_3017)
);

CKINVDCx14_ASAP7_75t_R g3018 ( 
.A(n_2625),
.Y(n_3018)
);

BUFx6f_ASAP7_75t_L g3019 ( 
.A(n_2483),
.Y(n_3019)
);

AOI22xp33_ASAP7_75t_L g3020 ( 
.A1(n_2637),
.A2(n_2283),
.B1(n_2343),
.B2(n_2236),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2643),
.B(n_2636),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2750),
.Y(n_3022)
);

BUFx12f_ASAP7_75t_L g3023 ( 
.A(n_2660),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2638),
.Y(n_3024)
);

INVx6_ASAP7_75t_L g3025 ( 
.A(n_2561),
.Y(n_3025)
);

INVx6_ASAP7_75t_L g3026 ( 
.A(n_2561),
.Y(n_3026)
);

AOI22xp33_ASAP7_75t_L g3027 ( 
.A1(n_2817),
.A2(n_2231),
.B1(n_2229),
.B2(n_2088),
.Y(n_3027)
);

NAND2x1p5_ASAP7_75t_L g3028 ( 
.A(n_2731),
.B(n_2084),
.Y(n_3028)
);

AOI22xp33_ASAP7_75t_L g3029 ( 
.A1(n_2818),
.A2(n_2403),
.B1(n_2408),
.B2(n_2155),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2657),
.Y(n_3030)
);

BUFx3_ASAP7_75t_L g3031 ( 
.A(n_2605),
.Y(n_3031)
);

INVx1_ASAP7_75t_SL g3032 ( 
.A(n_2492),
.Y(n_3032)
);

INVx1_ASAP7_75t_SL g3033 ( 
.A(n_2547),
.Y(n_3033)
);

AOI22xp33_ASAP7_75t_SL g3034 ( 
.A1(n_2807),
.A2(n_2422),
.B1(n_2176),
.B2(n_2192),
.Y(n_3034)
);

AOI22xp33_ASAP7_75t_SL g3035 ( 
.A1(n_2635),
.A2(n_2422),
.B1(n_2192),
.B2(n_2214),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2750),
.Y(n_3036)
);

BUFx2_ASAP7_75t_L g3037 ( 
.A(n_2503),
.Y(n_3037)
);

BUFx2_ASAP7_75t_L g3038 ( 
.A(n_2723),
.Y(n_3038)
);

BUFx2_ASAP7_75t_L g3039 ( 
.A(n_2517),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2794),
.Y(n_3040)
);

BUFx6f_ASAP7_75t_L g3041 ( 
.A(n_2483),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2794),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_SL g3043 ( 
.A1(n_2710),
.A2(n_2422),
.B1(n_2214),
.B2(n_2171),
.Y(n_3043)
);

AOI22xp33_ASAP7_75t_L g3044 ( 
.A1(n_2849),
.A2(n_2408),
.B1(n_2155),
.B2(n_2333),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2614),
.Y(n_3045)
);

CKINVDCx11_ASAP7_75t_R g3046 ( 
.A(n_2770),
.Y(n_3046)
);

BUFx10_ASAP7_75t_L g3047 ( 
.A(n_2632),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2716),
.Y(n_3048)
);

AOI22xp33_ASAP7_75t_SL g3049 ( 
.A1(n_2744),
.A2(n_2171),
.B1(n_2379),
.B2(n_2397),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2812),
.A2(n_2401),
.B(n_2070),
.Y(n_3050)
);

INVx6_ASAP7_75t_L g3051 ( 
.A(n_2524),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2718),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2555),
.A2(n_2271),
.B1(n_1998),
.B2(n_2026),
.Y(n_3053)
);

INVx1_ASAP7_75t_SL g3054 ( 
.A(n_2524),
.Y(n_3054)
);

OAI22xp33_ASAP7_75t_L g3055 ( 
.A1(n_2831),
.A2(n_2224),
.B1(n_2451),
.B2(n_2103),
.Y(n_3055)
);

CKINVDCx11_ASAP7_75t_R g3056 ( 
.A(n_2782),
.Y(n_3056)
);

INVx6_ASAP7_75t_L g3057 ( 
.A(n_2491),
.Y(n_3057)
);

AOI22xp33_ASAP7_75t_SL g3058 ( 
.A1(n_2744),
.A2(n_2379),
.B1(n_2401),
.B2(n_2304),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_SL g3059 ( 
.A1(n_2762),
.A2(n_2020),
.B1(n_2026),
.B2(n_2241),
.Y(n_3059)
);

INVx1_ASAP7_75t_SL g3060 ( 
.A(n_2732),
.Y(n_3060)
);

BUFx10_ASAP7_75t_L g3061 ( 
.A(n_2632),
.Y(n_3061)
);

BUFx10_ASAP7_75t_L g3062 ( 
.A(n_2549),
.Y(n_3062)
);

BUFx12f_ASAP7_75t_L g3063 ( 
.A(n_2543),
.Y(n_3063)
);

AOI21xp33_ASAP7_75t_L g3064 ( 
.A1(n_2628),
.A2(n_2465),
.B(n_2460),
.Y(n_3064)
);

AOI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2566),
.A2(n_2348),
.B1(n_2381),
.B2(n_2466),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_SL g3066 ( 
.A1(n_2762),
.A2(n_2242),
.B1(n_2247),
.B2(n_2241),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2615),
.Y(n_3067)
);

BUFx4f_ASAP7_75t_SL g3068 ( 
.A(n_2731),
.Y(n_3068)
);

BUFx3_ASAP7_75t_L g3069 ( 
.A(n_2552),
.Y(n_3069)
);

OAI22xp5_ASAP7_75t_L g3070 ( 
.A1(n_2776),
.A2(n_2811),
.B1(n_2819),
.B2(n_2695),
.Y(n_3070)
);

CKINVDCx20_ASAP7_75t_R g3071 ( 
.A(n_2645),
.Y(n_3071)
);

AOI22xp33_ASAP7_75t_L g3072 ( 
.A1(n_2668),
.A2(n_2381),
.B1(n_2220),
.B2(n_2213),
.Y(n_3072)
);

BUFx3_ASAP7_75t_L g3073 ( 
.A(n_2518),
.Y(n_3073)
);

INVx5_ASAP7_75t_L g3074 ( 
.A(n_2476),
.Y(n_3074)
);

INVx2_ASAP7_75t_SL g3075 ( 
.A(n_2717),
.Y(n_3075)
);

INVx1_ASAP7_75t_SL g3076 ( 
.A(n_2732),
.Y(n_3076)
);

AOI22xp33_ASAP7_75t_L g3077 ( 
.A1(n_2691),
.A2(n_2025),
.B1(n_1997),
.B2(n_2375),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2726),
.Y(n_3078)
);

INVx6_ASAP7_75t_L g3079 ( 
.A(n_2647),
.Y(n_3079)
);

INVx2_ASAP7_75t_SL g3080 ( 
.A(n_2717),
.Y(n_3080)
);

INVx6_ASAP7_75t_L g3081 ( 
.A(n_2647),
.Y(n_3081)
);

INVx1_ASAP7_75t_SL g3082 ( 
.A(n_2758),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2810),
.Y(n_3083)
);

INVx3_ASAP7_75t_L g3084 ( 
.A(n_2691),
.Y(n_3084)
);

INVx3_ASAP7_75t_L g3085 ( 
.A(n_2702),
.Y(n_3085)
);

BUFx6f_ASAP7_75t_L g3086 ( 
.A(n_2485),
.Y(n_3086)
);

OAI22xp5_ASAP7_75t_SL g3087 ( 
.A1(n_2833),
.A2(n_2067),
.B1(n_2413),
.B2(n_2420),
.Y(n_3087)
);

CKINVDCx6p67_ASAP7_75t_R g3088 ( 
.A(n_2725),
.Y(n_3088)
);

AOI22xp33_ASAP7_75t_SL g3089 ( 
.A1(n_2695),
.A2(n_2247),
.B1(n_2256),
.B2(n_2242),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2810),
.Y(n_3090)
);

BUFx6f_ASAP7_75t_SL g3091 ( 
.A(n_2739),
.Y(n_3091)
);

INVx8_ASAP7_75t_L g3092 ( 
.A(n_2557),
.Y(n_3092)
);

OAI22xp33_ASAP7_75t_L g3093 ( 
.A1(n_2687),
.A2(n_2036),
.B1(n_2042),
.B2(n_2043),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2702),
.B(n_2256),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2709),
.A2(n_2382),
.B1(n_2447),
.B2(n_2425),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2510),
.Y(n_3096)
);

OAI21xp5_ASAP7_75t_SL g3097 ( 
.A1(n_2788),
.A2(n_2034),
.B(n_2258),
.Y(n_3097)
);

CKINVDCx20_ASAP7_75t_R g3098 ( 
.A(n_2645),
.Y(n_3098)
);

AOI22xp33_ASAP7_75t_L g3099 ( 
.A1(n_2709),
.A2(n_2592),
.B1(n_2778),
.B2(n_2811),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_2851),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2510),
.Y(n_3101)
);

BUFx10_ASAP7_75t_L g3102 ( 
.A(n_2736),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2636),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2700),
.B(n_2064),
.Y(n_3104)
);

OAI21xp5_ASAP7_75t_SL g3105 ( 
.A1(n_2788),
.A2(n_2034),
.B(n_2258),
.Y(n_3105)
);

OAI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_2819),
.A2(n_2282),
.B1(n_2289),
.B2(n_2269),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2784),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2798),
.Y(n_3108)
);

AOI22xp33_ASAP7_75t_L g3109 ( 
.A1(n_2592),
.A2(n_2447),
.B1(n_2425),
.B2(n_2065),
.Y(n_3109)
);

BUFx6f_ASAP7_75t_L g3110 ( 
.A(n_2485),
.Y(n_3110)
);

CKINVDCx11_ASAP7_75t_R g3111 ( 
.A(n_2747),
.Y(n_3111)
);

CKINVDCx20_ASAP7_75t_R g3112 ( 
.A(n_2830),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2799),
.Y(n_3113)
);

AOI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_2764),
.A2(n_2282),
.B1(n_2289),
.B2(n_2269),
.Y(n_3114)
);

CKINVDCx5p33_ASAP7_75t_R g3115 ( 
.A(n_2598),
.Y(n_3115)
);

INVx4_ASAP7_75t_L g3116 ( 
.A(n_2590),
.Y(n_3116)
);

CKINVDCx6p67_ASAP7_75t_R g3117 ( 
.A(n_2806),
.Y(n_3117)
);

OAI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2687),
.A2(n_2792),
.B1(n_2649),
.B2(n_2766),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2841),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2846),
.Y(n_3120)
);

OAI22xp33_ASAP7_75t_L g3121 ( 
.A1(n_2687),
.A2(n_2071),
.B1(n_2086),
.B2(n_2080),
.Y(n_3121)
);

OR2x2_ASAP7_75t_L g3122 ( 
.A(n_2700),
.B(n_2092),
.Y(n_3122)
);

INVx4_ASAP7_75t_L g3123 ( 
.A(n_2590),
.Y(n_3123)
);

BUFx8_ASAP7_75t_SL g3124 ( 
.A(n_2651),
.Y(n_3124)
);

AND2x2_ASAP7_75t_L g3125 ( 
.A(n_2504),
.B(n_2113),
.Y(n_3125)
);

INVx6_ASAP7_75t_L g3126 ( 
.A(n_2735),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2808),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2577),
.B(n_2579),
.Y(n_3128)
);

INVx1_ASAP7_75t_SL g3129 ( 
.A(n_2584),
.Y(n_3129)
);

AOI22xp33_ASAP7_75t_SL g3130 ( 
.A1(n_2689),
.A2(n_2319),
.B1(n_2323),
.B2(n_2310),
.Y(n_3130)
);

CKINVDCx5p33_ASAP7_75t_R g3131 ( 
.A(n_2595),
.Y(n_3131)
);

INVx6_ASAP7_75t_L g3132 ( 
.A(n_2735),
.Y(n_3132)
);

OAI22xp5_ASAP7_75t_L g3133 ( 
.A1(n_2792),
.A2(n_2319),
.B1(n_2323),
.B2(n_2310),
.Y(n_3133)
);

CKINVDCx20_ASAP7_75t_R g3134 ( 
.A(n_2828),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2821),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2592),
.A2(n_2115),
.B1(n_2139),
.B2(n_2126),
.Y(n_3136)
);

INVx5_ASAP7_75t_L g3137 ( 
.A(n_2476),
.Y(n_3137)
);

BUFx4f_ASAP7_75t_SL g3138 ( 
.A(n_2651),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2727),
.A2(n_2157),
.B1(n_2186),
.B2(n_2179),
.Y(n_3139)
);

AOI22xp33_ASAP7_75t_SL g3140 ( 
.A1(n_2715),
.A2(n_2334),
.B1(n_2350),
.B2(n_2349),
.Y(n_3140)
);

OAI22xp5_ASAP7_75t_L g3141 ( 
.A1(n_2649),
.A2(n_2766),
.B1(n_2752),
.B2(n_2740),
.Y(n_3141)
);

INVx2_ASAP7_75t_SL g3142 ( 
.A(n_2736),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2832),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2835),
.Y(n_3144)
);

INVx2_ASAP7_75t_L g3145 ( 
.A(n_2837),
.Y(n_3145)
);

AOI22xp33_ASAP7_75t_L g3146 ( 
.A1(n_2727),
.A2(n_2349),
.B1(n_2350),
.B2(n_2334),
.Y(n_3146)
);

BUFx2_ASAP7_75t_L g3147 ( 
.A(n_2729),
.Y(n_3147)
);

OAI22xp33_ASAP7_75t_L g3148 ( 
.A1(n_2705),
.A2(n_2120),
.B1(n_2058),
.B2(n_2405),
.Y(n_3148)
);

BUFx2_ASAP7_75t_L g3149 ( 
.A(n_2619),
.Y(n_3149)
);

AOI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2730),
.A2(n_2201),
.B1(n_2221),
.B2(n_2217),
.Y(n_3150)
);

INVx4_ASAP7_75t_SL g3151 ( 
.A(n_2828),
.Y(n_3151)
);

OAI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_2740),
.A2(n_2414),
.B1(n_2415),
.B2(n_2409),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2820),
.Y(n_3153)
);

INVx4_ASAP7_75t_L g3154 ( 
.A(n_2590),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_2918),
.A2(n_2824),
.B1(n_2594),
.B2(n_2803),
.Y(n_3155)
);

BUFx4f_ASAP7_75t_SL g3156 ( 
.A(n_3023),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2871),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2993),
.B(n_2577),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2922),
.B(n_2579),
.Y(n_3159)
);

AOI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_2908),
.A2(n_2824),
.B1(n_3055),
.B2(n_2904),
.Y(n_3160)
);

NAND2x1p5_ASAP7_75t_L g3161 ( 
.A(n_3001),
.B(n_2602),
.Y(n_3161)
);

OAI22xp5_ASAP7_75t_L g3162 ( 
.A1(n_2863),
.A2(n_2653),
.B1(n_2665),
.B2(n_2602),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2877),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_SL g3164 ( 
.A1(n_3070),
.A2(n_2603),
.B1(n_2642),
.B2(n_2620),
.Y(n_3164)
);

OAI22xp5_ASAP7_75t_L g3165 ( 
.A1(n_2874),
.A2(n_2653),
.B1(n_2665),
.B2(n_2602),
.Y(n_3165)
);

OAI22xp5_ASAP7_75t_L g3166 ( 
.A1(n_2897),
.A2(n_2665),
.B1(n_2676),
.B2(n_2653),
.Y(n_3166)
);

BUFx3_ASAP7_75t_L g3167 ( 
.A(n_2894),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_3021),
.B(n_2584),
.Y(n_3168)
);

OAI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2924),
.A2(n_2676),
.B1(n_2829),
.B2(n_2812),
.Y(n_3169)
);

AOI22xp33_ASAP7_75t_L g3170 ( 
.A1(n_2883),
.A2(n_2594),
.B1(n_2803),
.B2(n_2790),
.Y(n_3170)
);

AOI22xp33_ASAP7_75t_L g3171 ( 
.A1(n_2936),
.A2(n_2804),
.B1(n_2790),
.B2(n_2617),
.Y(n_3171)
);

INVxp67_ASAP7_75t_L g3172 ( 
.A(n_3039),
.Y(n_3172)
);

HB1xp67_ASAP7_75t_L g3173 ( 
.A(n_3104),
.Y(n_3173)
);

AOI22xp33_ASAP7_75t_SL g3174 ( 
.A1(n_3001),
.A2(n_2721),
.B1(n_2701),
.B2(n_2676),
.Y(n_3174)
);

AOI22xp33_ASAP7_75t_L g3175 ( 
.A1(n_2861),
.A2(n_2928),
.B1(n_2952),
.B2(n_2975),
.Y(n_3175)
);

AOI22xp33_ASAP7_75t_SL g3176 ( 
.A1(n_3001),
.A2(n_2712),
.B1(n_2720),
.B2(n_2711),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2873),
.Y(n_3177)
);

INVx1_ASAP7_75t_L g3178 ( 
.A(n_3005),
.Y(n_3178)
);

AOI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2872),
.A2(n_2843),
.B1(n_2652),
.B2(n_2690),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2889),
.Y(n_3180)
);

OAI222xp33_ASAP7_75t_L g3181 ( 
.A1(n_3133),
.A2(n_2655),
.B1(n_2690),
.B2(n_2652),
.C1(n_2774),
.C2(n_2752),
.Y(n_3181)
);

CKINVDCx5p33_ASAP7_75t_R g3182 ( 
.A(n_3046),
.Y(n_3182)
);

AOI22xp33_ASAP7_75t_SL g3183 ( 
.A1(n_2998),
.A2(n_2722),
.B1(n_2667),
.B2(n_2669),
.Y(n_3183)
);

OAI22x1_ASAP7_75t_L g3184 ( 
.A1(n_2892),
.A2(n_2775),
.B1(n_2829),
.B2(n_2755),
.Y(n_3184)
);

AND2x2_ASAP7_75t_L g3185 ( 
.A(n_3128),
.B(n_2601),
.Y(n_3185)
);

BUFx6f_ASAP7_75t_L g3186 ( 
.A(n_2867),
.Y(n_3186)
);

HB1xp67_ASAP7_75t_L g3187 ( 
.A(n_2969),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2891),
.Y(n_3188)
);

INVx2_ASAP7_75t_L g3189 ( 
.A(n_2879),
.Y(n_3189)
);

CKINVDCx5p33_ASAP7_75t_R g3190 ( 
.A(n_3056),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2893),
.Y(n_3191)
);

OAI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_3114),
.A2(n_2655),
.B1(n_2774),
.B2(n_2775),
.Y(n_3192)
);

OAI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_3099),
.A2(n_2755),
.B1(n_2621),
.B2(n_2633),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2896),
.Y(n_3194)
);

AOI22xp33_ASAP7_75t_L g3195 ( 
.A1(n_2961),
.A2(n_2804),
.B1(n_2855),
.B2(n_2626),
.Y(n_3195)
);

NAND3xp33_ASAP7_75t_L g3196 ( 
.A(n_3006),
.B(n_2845),
.C(n_2855),
.Y(n_3196)
);

OAI22xp5_ASAP7_75t_L g3197 ( 
.A1(n_2943),
.A2(n_2629),
.B1(n_2654),
.B2(n_2781),
.Y(n_3197)
);

AOI222xp33_ASAP7_75t_L g3198 ( 
.A1(n_2880),
.A2(n_2666),
.B1(n_2697),
.B2(n_2641),
.C1(n_2644),
.C2(n_2627),
.Y(n_3198)
);

OAI21xp5_ASAP7_75t_SL g3199 ( 
.A1(n_2887),
.A2(n_2781),
.B(n_2761),
.Y(n_3199)
);

AOI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_2968),
.A2(n_2780),
.B1(n_2795),
.B2(n_2800),
.Y(n_3200)
);

INVx2_ASAP7_75t_L g3201 ( 
.A(n_2881),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_3087),
.A2(n_2780),
.B1(n_2801),
.B2(n_2845),
.Y(n_3202)
);

AOI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_2882),
.A2(n_2777),
.B1(n_2797),
.B2(n_2761),
.Y(n_3203)
);

AOI22xp33_ASAP7_75t_SL g3204 ( 
.A1(n_3037),
.A2(n_2677),
.B1(n_2694),
.B2(n_2662),
.Y(n_3204)
);

OAI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_2886),
.A2(n_2562),
.B1(n_2696),
.B2(n_2476),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_2967),
.A2(n_2562),
.B1(n_2696),
.B2(n_2515),
.Y(n_3206)
);

HB1xp67_ASAP7_75t_L g3207 ( 
.A(n_3122),
.Y(n_3207)
);

NAND3xp33_ASAP7_75t_L g3208 ( 
.A(n_3027),
.B(n_2477),
.C(n_2743),
.Y(n_3208)
);

AOI22xp33_ASAP7_75t_SL g3209 ( 
.A1(n_3106),
.A2(n_2515),
.B1(n_2537),
.B2(n_2488),
.Y(n_3209)
);

BUFx2_ASAP7_75t_L g3210 ( 
.A(n_3073),
.Y(n_3210)
);

AND2x2_ASAP7_75t_SL g3211 ( 
.A(n_2939),
.B(n_2475),
.Y(n_3211)
);

CKINVDCx20_ASAP7_75t_R g3212 ( 
.A(n_2970),
.Y(n_3212)
);

OAI22xp5_ASAP7_75t_L g3213 ( 
.A1(n_3146),
.A2(n_2515),
.B1(n_2537),
.B2(n_2488),
.Y(n_3213)
);

AOI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_2905),
.A2(n_2477),
.B1(n_2686),
.B2(n_2679),
.Y(n_3214)
);

AOI22xp33_ASAP7_75t_L g3215 ( 
.A1(n_2864),
.A2(n_2479),
.B1(n_2576),
.B2(n_2847),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2907),
.Y(n_3216)
);

OR2x2_ASAP7_75t_L g3217 ( 
.A(n_3129),
.B(n_2601),
.Y(n_3217)
);

OAI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_3066),
.A2(n_2537),
.B1(n_2488),
.B2(n_2507),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2911),
.Y(n_3219)
);

AOI22xp33_ASAP7_75t_SL g3220 ( 
.A1(n_3118),
.A2(n_2475),
.B1(n_2486),
.B2(n_2751),
.Y(n_3220)
);

INVx2_ASAP7_75t_L g3221 ( 
.A(n_2884),
.Y(n_3221)
);

AOI22xp33_ASAP7_75t_L g3222 ( 
.A1(n_3011),
.A2(n_2479),
.B1(n_2600),
.B2(n_2658),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2988),
.B(n_2793),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2912),
.Y(n_3224)
);

AOI22xp5_ASAP7_75t_L g3225 ( 
.A1(n_2925),
.A2(n_2793),
.B1(n_2671),
.B2(n_2673),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_L g3226 ( 
.A1(n_2962),
.A2(n_2680),
.B1(n_2693),
.B2(n_2664),
.Y(n_3226)
);

OAI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_3089),
.A2(n_2506),
.B1(n_2507),
.B2(n_2540),
.Y(n_3227)
);

OAI22xp5_ASAP7_75t_L g3228 ( 
.A1(n_2940),
.A2(n_2672),
.B1(n_2743),
.B2(n_2613),
.Y(n_3228)
);

INVx4_ASAP7_75t_L g3229 ( 
.A(n_2894),
.Y(n_3229)
);

INVx3_ASAP7_75t_L g3230 ( 
.A(n_2939),
.Y(n_3230)
);

AOI22xp33_ASAP7_75t_L g3231 ( 
.A1(n_2860),
.A2(n_2713),
.B1(n_2742),
.B2(n_2698),
.Y(n_3231)
);

CKINVDCx14_ASAP7_75t_R g3232 ( 
.A(n_2964),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2942),
.B(n_2613),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_3130),
.B(n_2678),
.Y(n_3234)
);

AOI22xp33_ASAP7_75t_SL g3235 ( 
.A1(n_2971),
.A2(n_2486),
.B1(n_2749),
.B2(n_2746),
.Y(n_3235)
);

NOR3xp33_ASAP7_75t_L g3236 ( 
.A(n_2946),
.B(n_2760),
.C(n_2859),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_2917),
.Y(n_3237)
);

OAI22xp5_ASAP7_75t_L g3238 ( 
.A1(n_2958),
.A2(n_2672),
.B1(n_2540),
.B2(n_2692),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_2919),
.Y(n_3239)
);

AOI211xp5_ASAP7_75t_L g3240 ( 
.A1(n_2866),
.A2(n_2714),
.B(n_2754),
.C(n_2745),
.Y(n_3240)
);

AOI22xp33_ASAP7_75t_L g3241 ( 
.A1(n_3022),
.A2(n_2769),
.B1(n_2816),
.B2(n_2783),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2885),
.Y(n_3242)
);

OAI22xp5_ASAP7_75t_L g3243 ( 
.A1(n_3029),
.A2(n_3136),
.B1(n_2921),
.B2(n_3044),
.Y(n_3243)
);

OAI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_2934),
.A2(n_2506),
.B1(n_2674),
.B2(n_2820),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2960),
.B(n_3004),
.Y(n_3245)
);

OAI22xp5_ASAP7_75t_L g3246 ( 
.A1(n_3140),
.A2(n_2674),
.B1(n_2853),
.B2(n_2834),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2923),
.Y(n_3247)
);

INVx1_ASAP7_75t_L g3248 ( 
.A(n_2927),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_2929),
.B(n_3045),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2932),
.Y(n_3250)
);

AOI22xp33_ASAP7_75t_L g3251 ( 
.A1(n_3036),
.A2(n_2823),
.B1(n_2840),
.B2(n_2827),
.Y(n_3251)
);

OAI21xp33_ASAP7_75t_L g3252 ( 
.A1(n_3053),
.A2(n_2563),
.B(n_2580),
.Y(n_3252)
);

OR2x6_ASAP7_75t_L g3253 ( 
.A(n_2976),
.B(n_2785),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_3040),
.A2(n_2842),
.B1(n_2844),
.B2(n_2707),
.Y(n_3254)
);

HB1xp67_ASAP7_75t_L g3255 ( 
.A(n_3125),
.Y(n_3255)
);

AOI22xp33_ASAP7_75t_L g3256 ( 
.A1(n_3042),
.A2(n_2707),
.B1(n_2697),
.B2(n_2659),
.Y(n_3256)
);

BUFx4f_ASAP7_75t_SL g3257 ( 
.A(n_2869),
.Y(n_3257)
);

AOI22xp33_ASAP7_75t_L g3258 ( 
.A1(n_3083),
.A2(n_2659),
.B1(n_2708),
.B2(n_2688),
.Y(n_3258)
);

AOI22xp33_ASAP7_75t_L g3259 ( 
.A1(n_3090),
.A2(n_2688),
.B1(n_2681),
.B2(n_2692),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_SL g3260 ( 
.A1(n_3092),
.A2(n_2618),
.B1(n_2473),
.B2(n_2678),
.Y(n_3260)
);

BUFx2_ASAP7_75t_L g3261 ( 
.A(n_2867),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_2937),
.Y(n_3262)
);

AOI22xp33_ASAP7_75t_L g3263 ( 
.A1(n_3020),
.A2(n_2681),
.B1(n_2548),
.B2(n_2550),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_L g3264 ( 
.A1(n_3016),
.A2(n_2548),
.B1(n_2550),
.B2(n_2618),
.Y(n_3264)
);

CKINVDCx11_ASAP7_75t_R g3265 ( 
.A(n_2901),
.Y(n_3265)
);

OAI22xp33_ASAP7_75t_L g3266 ( 
.A1(n_3075),
.A2(n_3080),
.B1(n_3060),
.B2(n_3076),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2938),
.Y(n_3267)
);

AOI22xp33_ASAP7_75t_L g3268 ( 
.A1(n_3014),
.A2(n_2618),
.B1(n_2856),
.B2(n_2853),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_2941),
.Y(n_3269)
);

OAI21xp33_ASAP7_75t_L g3270 ( 
.A1(n_2878),
.A2(n_2719),
.B(n_2834),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_L g3271 ( 
.A1(n_2916),
.A2(n_2618),
.B1(n_2856),
.B2(n_2857),
.Y(n_3271)
);

AOI22xp33_ASAP7_75t_SL g3272 ( 
.A1(n_3092),
.A2(n_2678),
.B1(n_2857),
.B2(n_2560),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_2979),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_2979),
.Y(n_3274)
);

INVx3_ASAP7_75t_SL g3275 ( 
.A(n_2868),
.Y(n_3275)
);

INVx3_ASAP7_75t_L g3276 ( 
.A(n_3074),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_2935),
.B(n_2756),
.Y(n_3277)
);

AOI22xp33_ASAP7_75t_SL g3278 ( 
.A1(n_3084),
.A2(n_2678),
.B1(n_2560),
.B2(n_2589),
.Y(n_3278)
);

BUFx3_ASAP7_75t_L g3279 ( 
.A(n_2999),
.Y(n_3279)
);

AND2x2_ASAP7_75t_L g3280 ( 
.A(n_3127),
.B(n_2719),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_2984),
.A2(n_2955),
.B1(n_3101),
.B2(n_3096),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_2898),
.Y(n_3282)
);

OAI21xp33_ASAP7_75t_L g3283 ( 
.A1(n_3103),
.A2(n_2773),
.B(n_2763),
.Y(n_3283)
);

OAI22xp5_ASAP7_75t_L g3284 ( 
.A1(n_3058),
.A2(n_2557),
.B1(n_2589),
.B2(n_2511),
.Y(n_3284)
);

AOI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_3007),
.A2(n_2500),
.B1(n_2678),
.B2(n_2791),
.Y(n_3285)
);

AOI22xp33_ASAP7_75t_L g3286 ( 
.A1(n_2862),
.A2(n_2500),
.B1(n_2544),
.B2(n_2513),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2947),
.Y(n_3287)
);

INVx1_ASAP7_75t_L g3288 ( 
.A(n_2980),
.Y(n_3288)
);

OAI21xp33_ASAP7_75t_L g3289 ( 
.A1(n_2963),
.A2(n_2737),
.B(n_2607),
.Y(n_3289)
);

OAI22xp5_ASAP7_75t_L g3290 ( 
.A1(n_3010),
.A2(n_2511),
.B1(n_2753),
.B2(n_2607),
.Y(n_3290)
);

AOI22xp33_ASAP7_75t_SL g3291 ( 
.A1(n_3084),
.A2(n_2544),
.B1(n_2513),
.B2(n_2597),
.Y(n_3291)
);

BUFx12f_ASAP7_75t_L g3292 ( 
.A(n_2996),
.Y(n_3292)
);

OAI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3049),
.A2(n_3059),
.B1(n_3109),
.B2(n_3043),
.Y(n_3293)
);

OAI21xp5_ASAP7_75t_SL g3294 ( 
.A1(n_3097),
.A2(n_2505),
.B(n_2597),
.Y(n_3294)
);

OAI21xp33_ASAP7_75t_L g3295 ( 
.A1(n_3013),
.A2(n_2737),
.B(n_2634),
.Y(n_3295)
);

HB1xp67_ASAP7_75t_L g3296 ( 
.A(n_3135),
.Y(n_3296)
);

NOR2xp33_ASAP7_75t_L g3297 ( 
.A(n_3112),
.B(n_2609),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_SL g3298 ( 
.A1(n_3085),
.A2(n_2914),
.B1(n_2992),
.B2(n_2902),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2980),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_3143),
.B(n_2609),
.Y(n_3300)
);

AOI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_3144),
.A2(n_2634),
.B1(n_2639),
.B2(n_2771),
.Y(n_3301)
);

INVx3_ASAP7_75t_SL g3302 ( 
.A(n_2868),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_SL g3303 ( 
.A1(n_3085),
.A2(n_2639),
.B1(n_2813),
.B2(n_2771),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3145),
.B(n_3032),
.Y(n_3304)
);

NAND3xp33_ASAP7_75t_L g3305 ( 
.A(n_3065),
.B(n_2753),
.C(n_2528),
.Y(n_3305)
);

INVx3_ASAP7_75t_SL g3306 ( 
.A(n_2870),
.Y(n_3306)
);

AOI21xp33_ASAP7_75t_L g3307 ( 
.A1(n_3093),
.A2(n_2815),
.B(n_2813),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_2949),
.Y(n_3308)
);

AOI22xp33_ASAP7_75t_SL g3309 ( 
.A1(n_2914),
.A2(n_2815),
.B1(n_2753),
.B2(n_2505),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_2867),
.B(n_251),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3067),
.Y(n_3311)
);

AOI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_2973),
.A2(n_2703),
.B1(n_2238),
.B2(n_2240),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3067),
.Y(n_3313)
);

AND2x2_ASAP7_75t_L g3314 ( 
.A(n_3082),
.B(n_253),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_L g3315 ( 
.A1(n_2973),
.A2(n_2703),
.B1(n_2253),
.B2(n_2255),
.Y(n_3315)
);

AOI21xp33_ASAP7_75t_L g3316 ( 
.A1(n_3121),
.A2(n_2131),
.B(n_2796),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_2977),
.A2(n_2257),
.B1(n_2276),
.B2(n_2222),
.Y(n_3317)
);

AOI211xp5_ASAP7_75t_L g3318 ( 
.A1(n_3105),
.A2(n_2120),
.B(n_2734),
.C(n_2682),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3012),
.B(n_2796),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_3017),
.B(n_2789),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_SL g3321 ( 
.A1(n_2992),
.A2(n_2826),
.B1(n_2839),
.B2(n_2789),
.Y(n_3321)
);

INVxp67_ASAP7_75t_L g3322 ( 
.A(n_2972),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3108),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3033),
.B(n_253),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3113),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3119),
.Y(n_3326)
);

INVx3_ASAP7_75t_L g3327 ( 
.A(n_3074),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2950),
.Y(n_3328)
);

BUFx3_ASAP7_75t_L g3329 ( 
.A(n_2956),
.Y(n_3329)
);

CKINVDCx5p33_ASAP7_75t_R g3330 ( 
.A(n_3000),
.Y(n_3330)
);

BUFx12f_ASAP7_75t_L g3331 ( 
.A(n_2865),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3120),
.Y(n_3332)
);

OAI21xp33_ASAP7_75t_L g3333 ( 
.A1(n_2906),
.A2(n_2278),
.B(n_2277),
.Y(n_3333)
);

BUFx3_ASAP7_75t_L g3334 ( 
.A(n_2876),
.Y(n_3334)
);

AND2x2_ASAP7_75t_L g3335 ( 
.A(n_2953),
.B(n_256),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_2977),
.A2(n_2279),
.B1(n_2308),
.B2(n_2301),
.Y(n_3336)
);

OAI22xp5_ASAP7_75t_L g3337 ( 
.A1(n_3035),
.A2(n_2789),
.B1(n_2839),
.B2(n_2826),
.Y(n_3337)
);

OAI22xp33_ASAP7_75t_L g3338 ( 
.A1(n_2948),
.A2(n_2826),
.B1(n_2848),
.B2(n_2839),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2957),
.Y(n_3339)
);

INVx2_ASAP7_75t_L g3340 ( 
.A(n_2965),
.Y(n_3340)
);

INVx2_ASAP7_75t_SL g3341 ( 
.A(n_2902),
.Y(n_3341)
);

CKINVDCx5p33_ASAP7_75t_R g3342 ( 
.A(n_2983),
.Y(n_3342)
);

OAI21xp5_ASAP7_75t_L g3343 ( 
.A1(n_3064),
.A2(n_2260),
.B(n_2682),
.Y(n_3343)
);

BUFx12f_ASAP7_75t_L g3344 ( 
.A(n_2986),
.Y(n_3344)
);

AOI22xp33_ASAP7_75t_L g3345 ( 
.A1(n_2951),
.A2(n_2336),
.B1(n_2359),
.B2(n_2351),
.Y(n_3345)
);

AOI22xp33_ASAP7_75t_L g3346 ( 
.A1(n_2951),
.A2(n_2131),
.B1(n_2436),
.B2(n_2848),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_2931),
.A2(n_2436),
.B1(n_2848),
.B2(n_2394),
.Y(n_3347)
);

OAI22xp5_ASAP7_75t_L g3348 ( 
.A1(n_2926),
.A2(n_2683),
.B1(n_2046),
.B2(n_2051),
.Y(n_3348)
);

AOI22xp33_ASAP7_75t_L g3349 ( 
.A1(n_2931),
.A2(n_2394),
.B1(n_2376),
.B2(n_2046),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_2903),
.B(n_256),
.Y(n_3350)
);

AO22x1_ASAP7_75t_L g3351 ( 
.A1(n_2890),
.A2(n_2485),
.B1(n_2516),
.B2(n_2512),
.Y(n_3351)
);

AOI22xp33_ASAP7_75t_SL g3352 ( 
.A1(n_3094),
.A2(n_2948),
.B1(n_3009),
.B2(n_2870),
.Y(n_3352)
);

OAI22xp5_ASAP7_75t_L g3353 ( 
.A1(n_3072),
.A2(n_2683),
.B1(n_2051),
.B2(n_2054),
.Y(n_3353)
);

AOI22xp33_ASAP7_75t_L g3354 ( 
.A1(n_3141),
.A2(n_3094),
.B1(n_2997),
.B2(n_3149),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2974),
.B(n_2193),
.Y(n_3355)
);

BUFx4f_ASAP7_75t_L g3356 ( 
.A(n_2930),
.Y(n_3356)
);

BUFx2_ASAP7_75t_L g3357 ( 
.A(n_3079),
.Y(n_3357)
);

AOI222xp33_ASAP7_75t_L g3358 ( 
.A1(n_2991),
.A2(n_260),
.B1(n_263),
.B2(n_258),
.C1(n_259),
.C2(n_261),
.Y(n_3358)
);

INVx3_ASAP7_75t_L g3359 ( 
.A(n_3074),
.Y(n_3359)
);

AOI22xp33_ASAP7_75t_L g3360 ( 
.A1(n_3147),
.A2(n_2394),
.B1(n_2054),
.B2(n_2056),
.Y(n_3360)
);

OR2x2_ASAP7_75t_L g3361 ( 
.A(n_2978),
.B(n_2981),
.Y(n_3361)
);

AOI22xp33_ASAP7_75t_L g3362 ( 
.A1(n_3038),
.A2(n_2056),
.B1(n_2045),
.B2(n_2193),
.Y(n_3362)
);

BUFx4f_ASAP7_75t_SL g3363 ( 
.A(n_3071),
.Y(n_3363)
);

AOI22xp33_ASAP7_75t_SL g3364 ( 
.A1(n_3009),
.A2(n_2512),
.B1(n_2535),
.B2(n_2516),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_2959),
.A2(n_2516),
.B1(n_2535),
.B2(n_2512),
.Y(n_3365)
);

CKINVDCx20_ASAP7_75t_R g3366 ( 
.A(n_3098),
.Y(n_3366)
);

OAI22xp5_ASAP7_75t_L g3367 ( 
.A1(n_3015),
.A2(n_2558),
.B1(n_2568),
.B2(n_2535),
.Y(n_3367)
);

CKINVDCx8_ASAP7_75t_R g3368 ( 
.A(n_3151),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_2995),
.B(n_2249),
.Y(n_3369)
);

INVx2_ASAP7_75t_SL g3370 ( 
.A(n_2899),
.Y(n_3370)
);

HB1xp67_ASAP7_75t_L g3371 ( 
.A(n_3002),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_3024),
.Y(n_3372)
);

AOI22xp5_ASAP7_75t_L g3373 ( 
.A1(n_3134),
.A2(n_2045),
.B1(n_2249),
.B2(n_2355),
.Y(n_3373)
);

AOI22xp33_ASAP7_75t_L g3374 ( 
.A1(n_2900),
.A2(n_2399),
.B1(n_2435),
.B2(n_2404),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_2909),
.A2(n_2399),
.B1(n_2435),
.B2(n_2404),
.Y(n_3375)
);

AOI22xp33_ASAP7_75t_SL g3376 ( 
.A1(n_3116),
.A2(n_2825),
.B1(n_2558),
.B2(n_2586),
.Y(n_3376)
);

INVx2_ASAP7_75t_SL g3377 ( 
.A(n_2990),
.Y(n_3377)
);

INVx1_ASAP7_75t_L g3378 ( 
.A(n_3030),
.Y(n_3378)
);

NOR2xp33_ASAP7_75t_L g3379 ( 
.A(n_2945),
.B(n_259),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_SL g3380 ( 
.A1(n_3116),
.A2(n_2558),
.B1(n_2586),
.B2(n_2568),
.Y(n_3380)
);

OAI22xp5_ASAP7_75t_L g3381 ( 
.A1(n_3139),
.A2(n_2355),
.B1(n_2586),
.B2(n_2568),
.Y(n_3381)
);

AOI22xp33_ASAP7_75t_SL g3382 ( 
.A1(n_3123),
.A2(n_3154),
.B1(n_3137),
.B2(n_2930),
.Y(n_3382)
);

INVx5_ASAP7_75t_SL g3383 ( 
.A(n_3117),
.Y(n_3383)
);

BUFx4f_ASAP7_75t_SL g3384 ( 
.A(n_3063),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_3048),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3052),
.Y(n_3386)
);

AOI22xp33_ASAP7_75t_SL g3387 ( 
.A1(n_3123),
.A2(n_2670),
.B1(n_2675),
.B2(n_2630),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3224),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3185),
.B(n_3078),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_SL g3390 ( 
.A(n_3235),
.B(n_3137),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3237),
.Y(n_3391)
);

AOI22xp33_ASAP7_75t_L g3392 ( 
.A1(n_3196),
.A2(n_2920),
.B1(n_2954),
.B2(n_3079),
.Y(n_3392)
);

AOI22xp33_ASAP7_75t_L g3393 ( 
.A1(n_3208),
.A2(n_3081),
.B1(n_3132),
.B2(n_3126),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3175),
.A2(n_3081),
.B1(n_3132),
.B2(n_3126),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3160),
.A2(n_3153),
.B1(n_3154),
.B2(n_3028),
.Y(n_3395)
);

AOI22xp33_ASAP7_75t_L g3396 ( 
.A1(n_3228),
.A2(n_3034),
.B1(n_3077),
.B2(n_2933),
.Y(n_3396)
);

OA21x2_ASAP7_75t_L g3397 ( 
.A1(n_3343),
.A2(n_3050),
.B(n_3107),
.Y(n_3397)
);

OAI21xp5_ASAP7_75t_SL g3398 ( 
.A1(n_3232),
.A2(n_3018),
.B(n_2875),
.Y(n_3398)
);

AOI22xp33_ASAP7_75t_L g3399 ( 
.A1(n_3184),
.A2(n_2933),
.B1(n_3111),
.B2(n_3152),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3207),
.B(n_3150),
.Y(n_3400)
);

AOI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_3199),
.A2(n_2944),
.B1(n_3091),
.B2(n_3138),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3159),
.B(n_2994),
.Y(n_3402)
);

OAI22xp33_ASAP7_75t_L g3403 ( 
.A1(n_3199),
.A2(n_3137),
.B1(n_3131),
.B2(n_3068),
.Y(n_3403)
);

NAND3xp33_ASAP7_75t_L g3404 ( 
.A(n_3358),
.B(n_3142),
.C(n_3095),
.Y(n_3404)
);

NOR3xp33_ASAP7_75t_L g3405 ( 
.A(n_3236),
.B(n_3054),
.C(n_3148),
.Y(n_3405)
);

AOI22xp33_ASAP7_75t_L g3406 ( 
.A1(n_3238),
.A2(n_3026),
.B1(n_3025),
.B2(n_3008),
.Y(n_3406)
);

AOI22xp5_ASAP7_75t_L g3407 ( 
.A1(n_3155),
.A2(n_3091),
.B1(n_2910),
.B2(n_3088),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3361),
.Y(n_3408)
);

AOI22xp33_ASAP7_75t_SL g3409 ( 
.A1(n_3227),
.A2(n_2982),
.B1(n_2910),
.B2(n_3025),
.Y(n_3409)
);

INVx2_ASAP7_75t_L g3410 ( 
.A(n_3371),
.Y(n_3410)
);

AOI21xp5_ASAP7_75t_SL g3411 ( 
.A1(n_3218),
.A2(n_3100),
.B(n_3031),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3158),
.B(n_3069),
.Y(n_3412)
);

OA21x2_ASAP7_75t_L g3413 ( 
.A1(n_3343),
.A2(n_2985),
.B(n_2966),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3173),
.B(n_3026),
.Y(n_3414)
);

OAI21xp5_ASAP7_75t_SL g3415 ( 
.A1(n_3352),
.A2(n_3358),
.B(n_3382),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3197),
.A2(n_3115),
.B1(n_2987),
.B2(n_3151),
.Y(n_3416)
);

OAI222xp33_ASAP7_75t_L g3417 ( 
.A1(n_3227),
.A2(n_2895),
.B1(n_2915),
.B2(n_3124),
.C1(n_2990),
.C2(n_2888),
.Y(n_3417)
);

AOI22xp33_ASAP7_75t_L g3418 ( 
.A1(n_3206),
.A2(n_3057),
.B1(n_3051),
.B2(n_3102),
.Y(n_3418)
);

AOI22xp33_ASAP7_75t_L g3419 ( 
.A1(n_3205),
.A2(n_3057),
.B1(n_3051),
.B2(n_3102),
.Y(n_3419)
);

OAI221xp5_ASAP7_75t_L g3420 ( 
.A1(n_3252),
.A2(n_2913),
.B1(n_2985),
.B2(n_2989),
.C(n_2966),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3171),
.A2(n_3110),
.B1(n_2985),
.B2(n_2989),
.Y(n_3421)
);

AOI22xp33_ASAP7_75t_L g3422 ( 
.A1(n_3195),
.A2(n_3062),
.B1(n_2989),
.B2(n_3003),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3255),
.B(n_3223),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3168),
.B(n_3304),
.Y(n_3424)
);

AOI22xp33_ASAP7_75t_L g3425 ( 
.A1(n_3198),
.A2(n_3062),
.B1(n_3003),
.B2(n_3019),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_3198),
.A2(n_3003),
.B1(n_3019),
.B2(n_2966),
.Y(n_3426)
);

AOI22xp33_ASAP7_75t_L g3427 ( 
.A1(n_3170),
.A2(n_3041),
.B1(n_3086),
.B2(n_3019),
.Y(n_3427)
);

AOI22xp33_ASAP7_75t_SL g3428 ( 
.A1(n_3246),
.A2(n_3047),
.B1(n_3061),
.B2(n_3041),
.Y(n_3428)
);

AOI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3293),
.A2(n_3086),
.B1(n_3041),
.B2(n_3110),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3246),
.A2(n_3110),
.B1(n_3086),
.B2(n_3061),
.Y(n_3430)
);

OAI21xp5_ASAP7_75t_L g3431 ( 
.A1(n_3333),
.A2(n_3047),
.B(n_264),
.Y(n_3431)
);

AOI22xp33_ASAP7_75t_L g3432 ( 
.A1(n_3244),
.A2(n_2404),
.B1(n_2435),
.B2(n_2399),
.Y(n_3432)
);

AND2x4_ASAP7_75t_L g3433 ( 
.A(n_3210),
.B(n_2630),
.Y(n_3433)
);

OAI222xp33_ASAP7_75t_L g3434 ( 
.A1(n_3244),
.A2(n_267),
.B1(n_269),
.B2(n_264),
.C1(n_266),
.C2(n_268),
.Y(n_3434)
);

AOI22xp33_ASAP7_75t_L g3435 ( 
.A1(n_3192),
.A2(n_2459),
.B1(n_2670),
.B2(n_2630),
.Y(n_3435)
);

NAND3xp33_ASAP7_75t_L g3436 ( 
.A(n_3281),
.B(n_2675),
.C(n_2670),
.Y(n_3436)
);

AOI22xp33_ASAP7_75t_L g3437 ( 
.A1(n_3193),
.A2(n_2459),
.B1(n_2733),
.B2(n_2675),
.Y(n_3437)
);

AOI22xp5_ASAP7_75t_L g3438 ( 
.A1(n_3243),
.A2(n_2733),
.B1(n_2757),
.B2(n_2738),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_SL g3439 ( 
.A1(n_3284),
.A2(n_2738),
.B1(n_2757),
.B2(n_2733),
.Y(n_3439)
);

AOI22xp33_ASAP7_75t_L g3440 ( 
.A1(n_3270),
.A2(n_3253),
.B1(n_3200),
.B2(n_3222),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3239),
.Y(n_3441)
);

AOI22xp33_ASAP7_75t_L g3442 ( 
.A1(n_3253),
.A2(n_2459),
.B1(n_2757),
.B2(n_2738),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3253),
.A2(n_2768),
.B1(n_2802),
.B2(n_2767),
.Y(n_3443)
);

OAI22xp5_ASAP7_75t_L g3444 ( 
.A1(n_3240),
.A2(n_2768),
.B1(n_2802),
.B2(n_2767),
.Y(n_3444)
);

AND2x2_ASAP7_75t_L g3445 ( 
.A(n_3296),
.B(n_266),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3163),
.B(n_267),
.Y(n_3446)
);

AOI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3215),
.A2(n_2768),
.B1(n_2802),
.B2(n_2767),
.Y(n_3447)
);

OAI222xp33_ASAP7_75t_L g3448 ( 
.A1(n_3164),
.A2(n_272),
.B1(n_274),
.B2(n_270),
.C1(n_271),
.C2(n_273),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3214),
.A2(n_3203),
.B1(n_3259),
.B2(n_3202),
.Y(n_3449)
);

INVx1_ASAP7_75t_L g3450 ( 
.A(n_3247),
.Y(n_3450)
);

OAI22xp5_ASAP7_75t_L g3451 ( 
.A1(n_3260),
.A2(n_2822),
.B1(n_2825),
.B2(n_2306),
.Y(n_3451)
);

AOI22xp33_ASAP7_75t_L g3452 ( 
.A1(n_3226),
.A2(n_2825),
.B1(n_2822),
.B2(n_2306),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_SL g3453 ( 
.A1(n_3218),
.A2(n_2822),
.B1(n_2306),
.B2(n_2307),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_L g3454 ( 
.A1(n_3264),
.A2(n_2307),
.B1(n_2324),
.B2(n_2297),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_SL g3455 ( 
.A1(n_3365),
.A2(n_2307),
.B1(n_2324),
.B2(n_2297),
.Y(n_3455)
);

AOI22xp33_ASAP7_75t_L g3456 ( 
.A1(n_3263),
.A2(n_2324),
.B1(n_2345),
.B2(n_2297),
.Y(n_3456)
);

OAI22xp5_ASAP7_75t_L g3457 ( 
.A1(n_3179),
.A2(n_2352),
.B1(n_2345),
.B2(n_2358),
.Y(n_3457)
);

INVx2_ASAP7_75t_L g3458 ( 
.A(n_3157),
.Y(n_3458)
);

AOI22xp33_ASAP7_75t_L g3459 ( 
.A1(n_3258),
.A2(n_2352),
.B1(n_2358),
.B2(n_2345),
.Y(n_3459)
);

INVx3_ASAP7_75t_L g3460 ( 
.A(n_3276),
.Y(n_3460)
);

AOI22xp33_ASAP7_75t_L g3461 ( 
.A1(n_3187),
.A2(n_2358),
.B1(n_2352),
.B2(n_2133),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3248),
.Y(n_3462)
);

AOI22xp33_ASAP7_75t_L g3463 ( 
.A1(n_3254),
.A2(n_2133),
.B1(n_2172),
.B2(n_2132),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3178),
.Y(n_3464)
);

AOI221xp5_ASAP7_75t_L g3465 ( 
.A1(n_3233),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.C(n_274),
.Y(n_3465)
);

AOI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_3231),
.A2(n_2172),
.B1(n_2177),
.B2(n_2133),
.Y(n_3466)
);

AOI22xp5_ASAP7_75t_L g3467 ( 
.A1(n_3256),
.A2(n_3268),
.B1(n_3225),
.B2(n_3266),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3177),
.Y(n_3468)
);

OAI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3294),
.A2(n_2177),
.B1(n_2189),
.B2(n_2172),
.Y(n_3469)
);

NOR3xp33_ASAP7_75t_L g3470 ( 
.A(n_3350),
.B(n_275),
.C(n_276),
.Y(n_3470)
);

OAI211xp5_ASAP7_75t_SL g3471 ( 
.A1(n_3172),
.A2(n_279),
.B(n_275),
.C(n_278),
.Y(n_3471)
);

OAI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3294),
.A2(n_2290),
.B1(n_2189),
.B2(n_2194),
.Y(n_3472)
);

AOI22xp33_ASAP7_75t_L g3473 ( 
.A1(n_3271),
.A2(n_2189),
.B1(n_2194),
.B2(n_2177),
.Y(n_3473)
);

AOI22xp33_ASAP7_75t_L g3474 ( 
.A1(n_3169),
.A2(n_2216),
.B1(n_2232),
.B2(n_2194),
.Y(n_3474)
);

AOI222xp33_ASAP7_75t_L g3475 ( 
.A1(n_3356),
.A2(n_3379),
.B1(n_3383),
.B2(n_3211),
.C1(n_3306),
.C2(n_3302),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3189),
.Y(n_3476)
);

AOI22xp33_ASAP7_75t_L g3477 ( 
.A1(n_3169),
.A2(n_2232),
.B1(n_2287),
.B2(n_2216),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3323),
.B(n_280),
.Y(n_3478)
);

AOI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3220),
.A2(n_2232),
.B1(n_2287),
.B2(n_2216),
.Y(n_3479)
);

OAI22xp5_ASAP7_75t_L g3480 ( 
.A1(n_3298),
.A2(n_2290),
.B1(n_2287),
.B2(n_282),
.Y(n_3480)
);

AOI22xp33_ASAP7_75t_L g3481 ( 
.A1(n_3310),
.A2(n_2290),
.B1(n_283),
.B2(n_280),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3180),
.Y(n_3482)
);

OAI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3230),
.A2(n_284),
.B1(n_281),
.B2(n_283),
.Y(n_3483)
);

OAI22xp5_ASAP7_75t_L g3484 ( 
.A1(n_3272),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3280),
.B(n_286),
.Y(n_3485)
);

AOI22xp33_ASAP7_75t_L g3486 ( 
.A1(n_3314),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_3486)
);

AOI22xp33_ASAP7_75t_SL g3487 ( 
.A1(n_3365),
.A2(n_290),
.B1(n_287),
.B2(n_289),
.Y(n_3487)
);

INVx2_ASAP7_75t_SL g3488 ( 
.A(n_3167),
.Y(n_3488)
);

AOI22xp33_ASAP7_75t_L g3489 ( 
.A1(n_3324),
.A2(n_293),
.B1(n_291),
.B2(n_292),
.Y(n_3489)
);

OAI22xp5_ASAP7_75t_L g3490 ( 
.A1(n_3354),
.A2(n_295),
.B1(n_292),
.B2(n_294),
.Y(n_3490)
);

AOI22xp33_ASAP7_75t_SL g3491 ( 
.A1(n_3367),
.A2(n_298),
.B1(n_295),
.B2(n_297),
.Y(n_3491)
);

BUFx2_ASAP7_75t_L g3492 ( 
.A(n_3357),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3201),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_SL g3494 ( 
.A1(n_3367),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_3494)
);

AOI222xp33_ASAP7_75t_L g3495 ( 
.A1(n_3356),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.C1(n_303),
.C2(n_304),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3325),
.B(n_301),
.Y(n_3496)
);

AOI22xp33_ASAP7_75t_L g3497 ( 
.A1(n_3289),
.A2(n_305),
.B1(n_302),
.B2(n_304),
.Y(n_3497)
);

AOI22xp33_ASAP7_75t_SL g3498 ( 
.A1(n_3166),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_3498)
);

NAND3xp33_ASAP7_75t_L g3499 ( 
.A(n_3217),
.B(n_310),
.C(n_313),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_SL g3500 ( 
.A1(n_3166),
.A2(n_315),
.B1(n_313),
.B2(n_314),
.Y(n_3500)
);

OAI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3345),
.A2(n_317),
.B1(n_314),
.B2(n_315),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_L g3502 ( 
.A1(n_3295),
.A2(n_3285),
.B1(n_3335),
.B2(n_3300),
.Y(n_3502)
);

OAI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3176),
.A2(n_3183),
.B1(n_3230),
.B2(n_3204),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_L g3504 ( 
.A(n_3326),
.B(n_318),
.Y(n_3504)
);

INVx3_ASAP7_75t_L g3505 ( 
.A(n_3276),
.Y(n_3505)
);

AOI22xp33_ASAP7_75t_SL g3506 ( 
.A1(n_3162),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_3506)
);

NAND3xp33_ASAP7_75t_L g3507 ( 
.A(n_3320),
.B(n_319),
.C(n_320),
.Y(n_3507)
);

OAI222xp33_ASAP7_75t_L g3508 ( 
.A1(n_3234),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.C1(n_324),
.C2(n_326),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_3309),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_3509)
);

NAND2xp5_ASAP7_75t_L g3510 ( 
.A(n_3332),
.B(n_327),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3188),
.B(n_329),
.Y(n_3511)
);

AO22x1_ASAP7_75t_L g3512 ( 
.A1(n_3229),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3191),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3250),
.A2(n_334),
.B1(n_331),
.B2(n_333),
.Y(n_3514)
);

AOI222xp33_ASAP7_75t_L g3515 ( 
.A1(n_3383),
.A2(n_333),
.B1(n_335),
.B2(n_337),
.C1(n_338),
.C2(n_339),
.Y(n_3515)
);

AOI22xp33_ASAP7_75t_L g3516 ( 
.A1(n_3262),
.A2(n_340),
.B1(n_335),
.B2(n_337),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3221),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3194),
.B(n_340),
.Y(n_3518)
);

AOI22xp33_ASAP7_75t_L g3519 ( 
.A1(n_3267),
.A2(n_345),
.B1(n_342),
.B2(n_344),
.Y(n_3519)
);

AOI22xp33_ASAP7_75t_L g3520 ( 
.A1(n_3269),
.A2(n_347),
.B1(n_342),
.B2(n_345),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3216),
.B(n_347),
.Y(n_3521)
);

AND2x2_ASAP7_75t_L g3522 ( 
.A(n_3219),
.B(n_348),
.Y(n_3522)
);

AOI22xp33_ASAP7_75t_L g3523 ( 
.A1(n_3283),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3305),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_3524)
);

AOI22xp33_ASAP7_75t_L g3525 ( 
.A1(n_3162),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_3525)
);

AOI22xp33_ASAP7_75t_L g3526 ( 
.A1(n_3297),
.A2(n_356),
.B1(n_353),
.B2(n_355),
.Y(n_3526)
);

AOI22xp33_ASAP7_75t_L g3527 ( 
.A1(n_3165),
.A2(n_362),
.B1(n_359),
.B2(n_361),
.Y(n_3527)
);

OAI22xp5_ASAP7_75t_L g3528 ( 
.A1(n_3278),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_3528)
);

NAND3xp33_ASAP7_75t_L g3529 ( 
.A(n_3301),
.B(n_364),
.C(n_365),
.Y(n_3529)
);

AOI22xp5_ASAP7_75t_L g3530 ( 
.A1(n_3241),
.A2(n_369),
.B1(n_367),
.B2(n_368),
.Y(n_3530)
);

AOI221xp5_ASAP7_75t_L g3531 ( 
.A1(n_3251),
.A2(n_367),
.B1(n_369),
.B2(n_371),
.C(n_372),
.Y(n_3531)
);

AOI211xp5_ASAP7_75t_L g3532 ( 
.A1(n_3338),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_3532)
);

AOI22xp33_ASAP7_75t_L g3533 ( 
.A1(n_3165),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_3533)
);

OAI222xp33_ASAP7_75t_L g3534 ( 
.A1(n_3303),
.A2(n_3291),
.B1(n_3209),
.B2(n_3368),
.C1(n_3213),
.C2(n_3229),
.Y(n_3534)
);

AOI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3286),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_3535)
);

OAI222xp33_ASAP7_75t_L g3536 ( 
.A1(n_3213),
.A2(n_376),
.B1(n_377),
.B2(n_379),
.C1(n_380),
.C2(n_381),
.Y(n_3536)
);

NAND3xp33_ASAP7_75t_L g3537 ( 
.A(n_3339),
.B(n_379),
.C(n_380),
.Y(n_3537)
);

OAI21xp33_ASAP7_75t_SL g3538 ( 
.A1(n_3377),
.A2(n_381),
.B(n_382),
.Y(n_3538)
);

AOI22xp33_ASAP7_75t_L g3539 ( 
.A1(n_3273),
.A2(n_386),
.B1(n_383),
.B2(n_385),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_SL g3540 ( 
.A(n_3409),
.B(n_3186),
.Y(n_3540)
);

NAND3xp33_ASAP7_75t_L g3541 ( 
.A(n_3409),
.B(n_3277),
.C(n_3322),
.Y(n_3541)
);

AND2x2_ASAP7_75t_L g3542 ( 
.A(n_3424),
.B(n_3274),
.Y(n_3542)
);

AND2x2_ASAP7_75t_L g3543 ( 
.A(n_3412),
.B(n_3288),
.Y(n_3543)
);

OA21x2_ASAP7_75t_L g3544 ( 
.A1(n_3534),
.A2(n_3315),
.B(n_3312),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_SL g3545 ( 
.A1(n_3503),
.A2(n_3383),
.B1(n_3359),
.B2(n_3327),
.Y(n_3545)
);

OAI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3487),
.A2(n_3181),
.B(n_3364),
.Y(n_3546)
);

AND2x2_ASAP7_75t_L g3547 ( 
.A(n_3410),
.B(n_3299),
.Y(n_3547)
);

AND2x2_ASAP7_75t_L g3548 ( 
.A(n_3402),
.B(n_3311),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3388),
.B(n_3313),
.Y(n_3549)
);

OAI21xp5_ASAP7_75t_SL g3550 ( 
.A1(n_3417),
.A2(n_3321),
.B(n_3174),
.Y(n_3550)
);

OAI22xp5_ASAP7_75t_L g3551 ( 
.A1(n_3428),
.A2(n_3336),
.B1(n_3317),
.B2(n_3319),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3408),
.B(n_3245),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3389),
.B(n_3242),
.Y(n_3553)
);

NAND3xp33_ASAP7_75t_L g3554 ( 
.A(n_3415),
.B(n_3249),
.C(n_3318),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3423),
.B(n_3282),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3391),
.B(n_3378),
.Y(n_3556)
);

AOI22xp33_ASAP7_75t_L g3557 ( 
.A1(n_3404),
.A2(n_3307),
.B1(n_3261),
.B2(n_3370),
.Y(n_3557)
);

AOI221xp5_ASAP7_75t_L g3558 ( 
.A1(n_3417),
.A2(n_3386),
.B1(n_3341),
.B2(n_3385),
.C(n_3328),
.Y(n_3558)
);

NAND2xp5_ASAP7_75t_L g3559 ( 
.A(n_3441),
.B(n_3287),
.Y(n_3559)
);

OAI21xp5_ASAP7_75t_SL g3560 ( 
.A1(n_3534),
.A2(n_3359),
.B(n_3327),
.Y(n_3560)
);

NAND3xp33_ASAP7_75t_L g3561 ( 
.A(n_3429),
.B(n_3362),
.C(n_3340),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3398),
.B(n_3275),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3492),
.B(n_3308),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3414),
.B(n_3372),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3450),
.B(n_3329),
.Y(n_3565)
);

OA21x2_ASAP7_75t_L g3566 ( 
.A1(n_3440),
.A2(n_3316),
.B(n_3355),
.Y(n_3566)
);

AOI21xp33_ASAP7_75t_SL g3567 ( 
.A1(n_3403),
.A2(n_3475),
.B(n_3401),
.Y(n_3567)
);

OA21x2_ASAP7_75t_L g3568 ( 
.A1(n_3426),
.A2(n_3369),
.B(n_3381),
.Y(n_3568)
);

NAND3xp33_ASAP7_75t_L g3569 ( 
.A(n_3428),
.B(n_3186),
.C(n_3376),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3462),
.B(n_3186),
.Y(n_3570)
);

AOI22xp33_ASAP7_75t_L g3571 ( 
.A1(n_3405),
.A2(n_3334),
.B1(n_3290),
.B2(n_3353),
.Y(n_3571)
);

AND2x2_ASAP7_75t_L g3572 ( 
.A(n_3464),
.B(n_3380),
.Y(n_3572)
);

AOI221xp5_ASAP7_75t_L g3573 ( 
.A1(n_3434),
.A2(n_3342),
.B1(n_3330),
.B2(n_3279),
.C(n_3190),
.Y(n_3573)
);

AND2x2_ASAP7_75t_L g3574 ( 
.A(n_3482),
.B(n_3387),
.Y(n_3574)
);

AOI221xp5_ASAP7_75t_L g3575 ( 
.A1(n_3434),
.A2(n_3182),
.B1(n_3337),
.B2(n_3346),
.C(n_3375),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3513),
.B(n_3351),
.Y(n_3576)
);

NAND4xp25_ASAP7_75t_L g3577 ( 
.A(n_3495),
.B(n_3347),
.C(n_3374),
.D(n_3360),
.Y(n_3577)
);

OA21x2_ASAP7_75t_L g3578 ( 
.A1(n_3436),
.A2(n_3349),
.B(n_3373),
.Y(n_3578)
);

NAND3xp33_ASAP7_75t_L g3579 ( 
.A(n_3399),
.B(n_3348),
.C(n_3265),
.Y(n_3579)
);

AOI21xp5_ASAP7_75t_SL g3580 ( 
.A1(n_3390),
.A2(n_3161),
.B(n_3156),
.Y(n_3580)
);

NAND3xp33_ASAP7_75t_L g3581 ( 
.A(n_3494),
.B(n_3366),
.C(n_3212),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_3458),
.B(n_3161),
.Y(n_3582)
);

AOI221xp5_ASAP7_75t_L g3583 ( 
.A1(n_3470),
.A2(n_383),
.B1(n_386),
.B2(n_387),
.C(n_388),
.Y(n_3583)
);

NAND3xp33_ASAP7_75t_L g3584 ( 
.A(n_3494),
.B(n_3257),
.C(n_389),
.Y(n_3584)
);

AND2x2_ASAP7_75t_L g3585 ( 
.A(n_3468),
.B(n_3476),
.Y(n_3585)
);

NAND3xp33_ASAP7_75t_L g3586 ( 
.A(n_3487),
.B(n_390),
.C(n_391),
.Y(n_3586)
);

OAI21xp33_ASAP7_75t_L g3587 ( 
.A1(n_3425),
.A2(n_391),
.B(n_393),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3493),
.B(n_394),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3517),
.B(n_394),
.Y(n_3589)
);

AND2x2_ASAP7_75t_L g3590 ( 
.A(n_3485),
.B(n_395),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3433),
.B(n_396),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_SL g3592 ( 
.A(n_3469),
.B(n_3363),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3400),
.B(n_396),
.Y(n_3593)
);

AO22x1_ASAP7_75t_L g3594 ( 
.A1(n_3431),
.A2(n_3292),
.B1(n_3344),
.B2(n_3384),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3433),
.B(n_3445),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_SL g3596 ( 
.A(n_3472),
.B(n_3331),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3502),
.B(n_397),
.Y(n_3597)
);

OAI21xp33_ASAP7_75t_L g3598 ( 
.A1(n_3430),
.A2(n_398),
.B(n_399),
.Y(n_3598)
);

NAND3xp33_ASAP7_75t_L g3599 ( 
.A(n_3392),
.B(n_399),
.C(n_400),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3511),
.B(n_400),
.Y(n_3600)
);

OAI22xp5_ASAP7_75t_SL g3601 ( 
.A1(n_3407),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_3601)
);

NOR3xp33_ASAP7_75t_L g3602 ( 
.A(n_3448),
.B(n_401),
.C(n_404),
.Y(n_3602)
);

NAND2xp5_ASAP7_75t_L g3603 ( 
.A(n_3518),
.B(n_406),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3521),
.B(n_406),
.Y(n_3604)
);

AOI221xp5_ASAP7_75t_L g3605 ( 
.A1(n_3448),
.A2(n_3536),
.B1(n_3449),
.B2(n_3508),
.C(n_3483),
.Y(n_3605)
);

OAI21xp5_ASAP7_75t_SL g3606 ( 
.A1(n_3416),
.A2(n_407),
.B(n_408),
.Y(n_3606)
);

AOI22xp33_ASAP7_75t_L g3607 ( 
.A1(n_3491),
.A2(n_408),
.B1(n_410),
.B2(n_411),
.Y(n_3607)
);

NOR2xp33_ASAP7_75t_R g3608 ( 
.A(n_3488),
.B(n_410),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3467),
.B(n_3432),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3460),
.B(n_412),
.Y(n_3610)
);

AND2x2_ASAP7_75t_L g3611 ( 
.A(n_3460),
.B(n_413),
.Y(n_3611)
);

AND2x2_ASAP7_75t_L g3612 ( 
.A(n_3505),
.B(n_413),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3522),
.B(n_415),
.Y(n_3613)
);

AOI221xp5_ASAP7_75t_L g3614 ( 
.A1(n_3536),
.A2(n_415),
.B1(n_416),
.B2(n_417),
.C(n_419),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3437),
.B(n_416),
.Y(n_3615)
);

AOI221xp5_ASAP7_75t_L g3616 ( 
.A1(n_3508),
.A2(n_417),
.B1(n_419),
.B2(n_420),
.C(n_423),
.Y(n_3616)
);

NAND3xp33_ASAP7_75t_L g3617 ( 
.A(n_3545),
.B(n_3500),
.C(n_3498),
.Y(n_3617)
);

OAI22xp33_ASAP7_75t_SL g3618 ( 
.A1(n_3540),
.A2(n_3505),
.B1(n_3420),
.B2(n_3444),
.Y(n_3618)
);

NAND3xp33_ASAP7_75t_L g3619 ( 
.A(n_3554),
.B(n_3500),
.C(n_3498),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3549),
.Y(n_3620)
);

NAND3xp33_ASAP7_75t_L g3621 ( 
.A(n_3567),
.B(n_3515),
.C(n_3499),
.Y(n_3621)
);

OR2x2_ASAP7_75t_L g3622 ( 
.A(n_3542),
.B(n_3435),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3547),
.B(n_3585),
.Y(n_3623)
);

INVx2_ASAP7_75t_SL g3624 ( 
.A(n_3565),
.Y(n_3624)
);

NOR3xp33_ASAP7_75t_L g3625 ( 
.A(n_3573),
.B(n_3512),
.C(n_3538),
.Y(n_3625)
);

OAI211xp5_ASAP7_75t_SL g3626 ( 
.A1(n_3605),
.A2(n_3411),
.B(n_3406),
.C(n_3396),
.Y(n_3626)
);

AND2x2_ASAP7_75t_L g3627 ( 
.A(n_3595),
.B(n_3555),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3553),
.B(n_3438),
.Y(n_3628)
);

NAND3xp33_ASAP7_75t_L g3629 ( 
.A(n_3560),
.B(n_3532),
.C(n_3507),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3543),
.B(n_3443),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3563),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3602),
.A2(n_3506),
.B1(n_3471),
.B2(n_3418),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3552),
.B(n_3446),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3548),
.B(n_3478),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3559),
.B(n_3397),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_3564),
.B(n_3496),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_L g3637 ( 
.A(n_3549),
.B(n_3397),
.Y(n_3637)
);

AOI221x1_ASAP7_75t_SL g3638 ( 
.A1(n_3581),
.A2(n_3510),
.B1(n_3504),
.B2(n_3490),
.C(n_3421),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3572),
.B(n_3442),
.Y(n_3639)
);

AO21x2_ASAP7_75t_L g3640 ( 
.A1(n_3576),
.A2(n_3537),
.B(n_3529),
.Y(n_3640)
);

AOI211xp5_ASAP7_75t_L g3641 ( 
.A1(n_3594),
.A2(n_3451),
.B(n_3480),
.C(n_3509),
.Y(n_3641)
);

OR2x2_ASAP7_75t_L g3642 ( 
.A(n_3556),
.B(n_3413),
.Y(n_3642)
);

NOR3xp33_ASAP7_75t_L g3643 ( 
.A(n_3606),
.B(n_3471),
.C(n_3484),
.Y(n_3643)
);

NAND3xp33_ASAP7_75t_L g3644 ( 
.A(n_3557),
.B(n_3394),
.C(n_3393),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3574),
.B(n_3422),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3576),
.Y(n_3646)
);

AOI22xp33_ASAP7_75t_L g3647 ( 
.A1(n_3609),
.A2(n_3395),
.B1(n_3419),
.B2(n_3528),
.Y(n_3647)
);

INVx2_ASAP7_75t_SL g3648 ( 
.A(n_3608),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3570),
.Y(n_3649)
);

NOR2xp33_ASAP7_75t_R g3650 ( 
.A(n_3562),
.B(n_424),
.Y(n_3650)
);

NAND4xp75_ASAP7_75t_L g3651 ( 
.A(n_3596),
.B(n_3479),
.C(n_3535),
.D(n_3465),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3582),
.B(n_3427),
.Y(n_3652)
);

AND2x2_ASAP7_75t_L g3653 ( 
.A(n_3568),
.B(n_3439),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3566),
.B(n_3413),
.Y(n_3654)
);

AOI221xp5_ASAP7_75t_L g3655 ( 
.A1(n_3593),
.A2(n_3486),
.B1(n_3489),
.B2(n_3526),
.C(n_3501),
.Y(n_3655)
);

AND2x2_ASAP7_75t_L g3656 ( 
.A(n_3568),
.B(n_3447),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3566),
.B(n_3474),
.Y(n_3657)
);

AND2x2_ASAP7_75t_L g3658 ( 
.A(n_3609),
.B(n_3477),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_L g3659 ( 
.A(n_3544),
.B(n_3466),
.Y(n_3659)
);

NOR3xp33_ASAP7_75t_L g3660 ( 
.A(n_3584),
.B(n_3531),
.C(n_3455),
.Y(n_3660)
);

OAI211xp5_ASAP7_75t_L g3661 ( 
.A1(n_3550),
.A2(n_3453),
.B(n_3524),
.C(n_3527),
.Y(n_3661)
);

AND2x4_ASAP7_75t_L g3662 ( 
.A(n_3569),
.B(n_3452),
.Y(n_3662)
);

NOR3xp33_ASAP7_75t_L g3663 ( 
.A(n_3599),
.B(n_3457),
.C(n_3530),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3588),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3591),
.B(n_3454),
.Y(n_3665)
);

NAND3xp33_ASAP7_75t_L g3666 ( 
.A(n_3558),
.B(n_3497),
.C(n_3523),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3593),
.B(n_3597),
.Y(n_3667)
);

NAND3xp33_ASAP7_75t_L g3668 ( 
.A(n_3546),
.B(n_3533),
.C(n_3525),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_SL g3669 ( 
.A(n_3546),
.B(n_3461),
.Y(n_3669)
);

INVx2_ASAP7_75t_SL g3670 ( 
.A(n_3610),
.Y(n_3670)
);

NAND2xp5_ASAP7_75t_L g3671 ( 
.A(n_3544),
.B(n_3456),
.Y(n_3671)
);

AND2x2_ASAP7_75t_L g3672 ( 
.A(n_3578),
.B(n_3463),
.Y(n_3672)
);

NOR3xp33_ASAP7_75t_L g3673 ( 
.A(n_3587),
.B(n_3481),
.C(n_3514),
.Y(n_3673)
);

AO21x2_ASAP7_75t_L g3674 ( 
.A1(n_3588),
.A2(n_3459),
.B(n_3473),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_3589),
.B(n_3516),
.Y(n_3675)
);

AND2x2_ASAP7_75t_L g3676 ( 
.A(n_3578),
.B(n_3519),
.Y(n_3676)
);

CKINVDCx8_ASAP7_75t_R g3677 ( 
.A(n_3662),
.Y(n_3677)
);

XNOR2xp5_ASAP7_75t_L g3678 ( 
.A(n_3648),
.B(n_3579),
.Y(n_3678)
);

INVx2_ASAP7_75t_SL g3679 ( 
.A(n_3624),
.Y(n_3679)
);

INVx1_ASAP7_75t_SL g3680 ( 
.A(n_3642),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3631),
.Y(n_3681)
);

OAI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3617),
.A2(n_3541),
.B1(n_3571),
.B2(n_3586),
.Y(n_3682)
);

AND2x2_ASAP7_75t_L g3683 ( 
.A(n_3627),
.B(n_3590),
.Y(n_3683)
);

BUFx3_ASAP7_75t_L g3684 ( 
.A(n_3623),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3626),
.B(n_3580),
.Y(n_3685)
);

INVx2_ASAP7_75t_L g3686 ( 
.A(n_3649),
.Y(n_3686)
);

NOR2xp33_ASAP7_75t_L g3687 ( 
.A(n_3621),
.B(n_3592),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_L g3688 ( 
.A(n_3669),
.B(n_3577),
.Y(n_3688)
);

NAND4xp75_ASAP7_75t_L g3689 ( 
.A(n_3676),
.B(n_3575),
.C(n_3611),
.D(n_3612),
.Y(n_3689)
);

AND2x2_ASAP7_75t_L g3690 ( 
.A(n_3646),
.B(n_3551),
.Y(n_3690)
);

INVxp67_ASAP7_75t_L g3691 ( 
.A(n_3645),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3658),
.B(n_3589),
.Y(n_3692)
);

NAND4xp75_ASAP7_75t_L g3693 ( 
.A(n_3653),
.B(n_3613),
.C(n_3616),
.D(n_3614),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3630),
.B(n_3551),
.Y(n_3694)
);

NAND4xp75_ASAP7_75t_SL g3695 ( 
.A(n_3657),
.B(n_3601),
.C(n_3598),
.D(n_3583),
.Y(n_3695)
);

INVx1_ASAP7_75t_L g3696 ( 
.A(n_3620),
.Y(n_3696)
);

INVxp67_ASAP7_75t_SL g3697 ( 
.A(n_3635),
.Y(n_3697)
);

XNOR2xp5_ASAP7_75t_L g3698 ( 
.A(n_3638),
.B(n_3623),
.Y(n_3698)
);

INVx3_ASAP7_75t_L g3699 ( 
.A(n_3662),
.Y(n_3699)
);

AND2x2_ASAP7_75t_L g3700 ( 
.A(n_3639),
.B(n_3561),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3664),
.Y(n_3701)
);

XNOR2xp5_ASAP7_75t_L g3702 ( 
.A(n_3638),
.B(n_3600),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3622),
.Y(n_3703)
);

NOR2x1_ASAP7_75t_R g3704 ( 
.A(n_3650),
.B(n_3613),
.Y(n_3704)
);

INVx5_ASAP7_75t_L g3705 ( 
.A(n_3672),
.Y(n_3705)
);

HB1xp67_ASAP7_75t_L g3706 ( 
.A(n_3635),
.Y(n_3706)
);

AND2x4_ASAP7_75t_L g3707 ( 
.A(n_3656),
.B(n_3615),
.Y(n_3707)
);

NAND4xp75_ASAP7_75t_L g3708 ( 
.A(n_3671),
.B(n_3604),
.C(n_3603),
.D(n_3615),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3671),
.B(n_3520),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3633),
.Y(n_3710)
);

AND4x1_ASAP7_75t_L g3711 ( 
.A(n_3641),
.B(n_3607),
.C(n_3539),
.D(n_427),
.Y(n_3711)
);

INVx1_ASAP7_75t_L g3712 ( 
.A(n_3628),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3637),
.Y(n_3713)
);

AOI22xp5_ASAP7_75t_L g3714 ( 
.A1(n_3619),
.A2(n_3668),
.B1(n_3625),
.B2(n_3629),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3637),
.Y(n_3715)
);

XNOR2xp5_ASAP7_75t_L g3716 ( 
.A(n_3644),
.B(n_424),
.Y(n_3716)
);

XOR2xp5_ASAP7_75t_L g3717 ( 
.A(n_3636),
.B(n_425),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3634),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3659),
.B(n_3652),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3670),
.Y(n_3720)
);

INVx2_ASAP7_75t_SL g3721 ( 
.A(n_3665),
.Y(n_3721)
);

NAND4xp75_ASAP7_75t_L g3722 ( 
.A(n_3659),
.B(n_425),
.C(n_427),
.D(n_428),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3674),
.B(n_428),
.Y(n_3723)
);

INVx1_ASAP7_75t_SL g3724 ( 
.A(n_3667),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3674),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3654),
.B(n_3640),
.Y(n_3726)
);

XOR2x2_ASAP7_75t_L g3727 ( 
.A(n_3651),
.B(n_430),
.Y(n_3727)
);

XOR2x2_ASAP7_75t_L g3728 ( 
.A(n_3678),
.B(n_3618),
.Y(n_3728)
);

INVx2_ASAP7_75t_SL g3729 ( 
.A(n_3679),
.Y(n_3729)
);

INVx2_ASAP7_75t_L g3730 ( 
.A(n_3684),
.Y(n_3730)
);

HB1xp67_ASAP7_75t_L g3731 ( 
.A(n_3706),
.Y(n_3731)
);

INVx1_ASAP7_75t_SL g3732 ( 
.A(n_3717),
.Y(n_3732)
);

INVxp67_ASAP7_75t_L g3733 ( 
.A(n_3687),
.Y(n_3733)
);

INVx2_ASAP7_75t_L g3734 ( 
.A(n_3686),
.Y(n_3734)
);

XNOR2xp5_ASAP7_75t_L g3735 ( 
.A(n_3727),
.B(n_3647),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3696),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3705),
.B(n_3654),
.Y(n_3737)
);

XNOR2xp5_ASAP7_75t_L g3738 ( 
.A(n_3689),
.B(n_3661),
.Y(n_3738)
);

AND2x2_ASAP7_75t_L g3739 ( 
.A(n_3705),
.B(n_3640),
.Y(n_3739)
);

AOI22xp5_ASAP7_75t_L g3740 ( 
.A1(n_3682),
.A2(n_3660),
.B1(n_3643),
.B2(n_3666),
.Y(n_3740)
);

XNOR2xp5_ASAP7_75t_L g3741 ( 
.A(n_3716),
.B(n_3632),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3701),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3703),
.Y(n_3743)
);

INVx1_ASAP7_75t_L g3744 ( 
.A(n_3713),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3715),
.Y(n_3745)
);

INVxp67_ASAP7_75t_L g3746 ( 
.A(n_3723),
.Y(n_3746)
);

INVx1_ASAP7_75t_SL g3747 ( 
.A(n_3724),
.Y(n_3747)
);

INVx1_ASAP7_75t_SL g3748 ( 
.A(n_3724),
.Y(n_3748)
);

XOR2x2_ASAP7_75t_L g3749 ( 
.A(n_3714),
.B(n_3688),
.Y(n_3749)
);

INVx2_ASAP7_75t_L g3750 ( 
.A(n_3680),
.Y(n_3750)
);

OR2x2_ASAP7_75t_L g3751 ( 
.A(n_3697),
.B(n_3680),
.Y(n_3751)
);

XOR2x2_ASAP7_75t_L g3752 ( 
.A(n_3714),
.B(n_3673),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3712),
.Y(n_3753)
);

OR2x2_ASAP7_75t_L g3754 ( 
.A(n_3719),
.B(n_3675),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3710),
.Y(n_3755)
);

INVx2_ASAP7_75t_L g3756 ( 
.A(n_3681),
.Y(n_3756)
);

XOR2x2_ASAP7_75t_L g3757 ( 
.A(n_3702),
.B(n_3663),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3753),
.Y(n_3758)
);

INVx1_ASAP7_75t_L g3759 ( 
.A(n_3744),
.Y(n_3759)
);

OA22x2_ASAP7_75t_L g3760 ( 
.A1(n_3740),
.A2(n_3698),
.B1(n_3699),
.B2(n_3682),
.Y(n_3760)
);

INVx3_ASAP7_75t_L g3761 ( 
.A(n_3730),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3731),
.Y(n_3762)
);

OAI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3730),
.A2(n_3677),
.B1(n_3699),
.B2(n_3705),
.Y(n_3763)
);

OAI22x1_ASAP7_75t_L g3764 ( 
.A1(n_3738),
.A2(n_3725),
.B1(n_3685),
.B2(n_3726),
.Y(n_3764)
);

OAI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_3733),
.A2(n_3691),
.B1(n_3694),
.B2(n_3707),
.Y(n_3765)
);

AOI22xp5_ASAP7_75t_L g3766 ( 
.A1(n_3749),
.A2(n_3707),
.B1(n_3690),
.B2(n_3700),
.Y(n_3766)
);

OA22x2_ASAP7_75t_L g3767 ( 
.A1(n_3733),
.A2(n_3721),
.B1(n_3683),
.B2(n_3718),
.Y(n_3767)
);

INVxp67_ASAP7_75t_L g3768 ( 
.A(n_3732),
.Y(n_3768)
);

OA22x2_ASAP7_75t_L g3769 ( 
.A1(n_3746),
.A2(n_3709),
.B1(n_3720),
.B2(n_3692),
.Y(n_3769)
);

AO22x2_ASAP7_75t_L g3770 ( 
.A1(n_3739),
.A2(n_3695),
.B1(n_3708),
.B2(n_3693),
.Y(n_3770)
);

AO22x1_ASAP7_75t_L g3771 ( 
.A1(n_3746),
.A2(n_3704),
.B1(n_3675),
.B2(n_3711),
.Y(n_3771)
);

INVx1_ASAP7_75t_L g3772 ( 
.A(n_3731),
.Y(n_3772)
);

OAI22xp33_ASAP7_75t_SL g3773 ( 
.A1(n_3751),
.A2(n_3729),
.B1(n_3754),
.B2(n_3748),
.Y(n_3773)
);

INVx1_ASAP7_75t_SL g3774 ( 
.A(n_3747),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3750),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3750),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3755),
.Y(n_3777)
);

CKINVDCx5p33_ASAP7_75t_R g3778 ( 
.A(n_3749),
.Y(n_3778)
);

OA22x2_ASAP7_75t_L g3779 ( 
.A1(n_3735),
.A2(n_3704),
.B1(n_3711),
.B2(n_3722),
.Y(n_3779)
);

INVx2_ASAP7_75t_SL g3780 ( 
.A(n_3756),
.Y(n_3780)
);

INVx2_ASAP7_75t_SL g3781 ( 
.A(n_3756),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3736),
.Y(n_3782)
);

XOR2x2_ASAP7_75t_L g3783 ( 
.A(n_3728),
.B(n_3655),
.Y(n_3783)
);

INVx2_ASAP7_75t_SL g3784 ( 
.A(n_3737),
.Y(n_3784)
);

OA22x2_ASAP7_75t_SL g3785 ( 
.A1(n_3752),
.A2(n_431),
.B1(n_433),
.B2(n_435),
.Y(n_3785)
);

XOR2x2_ASAP7_75t_L g3786 ( 
.A(n_3757),
.B(n_433),
.Y(n_3786)
);

BUFx12f_ASAP7_75t_L g3787 ( 
.A(n_3757),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3742),
.Y(n_3788)
);

INVxp67_ASAP7_75t_L g3789 ( 
.A(n_3741),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3743),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3734),
.Y(n_3791)
);

INVx1_ASAP7_75t_L g3792 ( 
.A(n_3762),
.Y(n_3792)
);

BUFx2_ASAP7_75t_L g3793 ( 
.A(n_3761),
.Y(n_3793)
);

BUFx2_ASAP7_75t_L g3794 ( 
.A(n_3768),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3772),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3774),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_3775),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3776),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3759),
.Y(n_3799)
);

AOI322xp5_ASAP7_75t_L g3800 ( 
.A1(n_3787),
.A2(n_3745),
.A3(n_3734),
.B1(n_437),
.B2(n_438),
.C1(n_439),
.C2(n_440),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3759),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3758),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3791),
.Y(n_3803)
);

INVx2_ASAP7_75t_SL g3804 ( 
.A(n_3784),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3777),
.Y(n_3805)
);

NOR2x1_ASAP7_75t_SL g3806 ( 
.A(n_3763),
.B(n_3745),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3782),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3788),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3790),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3766),
.B(n_435),
.Y(n_3810)
);

BUFx2_ASAP7_75t_L g3811 ( 
.A(n_3767),
.Y(n_3811)
);

INVxp67_ASAP7_75t_L g3812 ( 
.A(n_3789),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3780),
.Y(n_3813)
);

XOR2x2_ASAP7_75t_L g3814 ( 
.A(n_3783),
.B(n_436),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3781),
.Y(n_3815)
);

INVx1_ASAP7_75t_L g3816 ( 
.A(n_3773),
.Y(n_3816)
);

AOI22xp5_ASAP7_75t_L g3817 ( 
.A1(n_3811),
.A2(n_3760),
.B1(n_3770),
.B2(n_3771),
.Y(n_3817)
);

BUFx4f_ASAP7_75t_SL g3818 ( 
.A(n_3796),
.Y(n_3818)
);

AOI31xp33_ASAP7_75t_L g3819 ( 
.A1(n_3812),
.A2(n_3778),
.A3(n_3786),
.B(n_3770),
.Y(n_3819)
);

AOI22xp5_ASAP7_75t_L g3820 ( 
.A1(n_3804),
.A2(n_3771),
.B1(n_3779),
.B2(n_3764),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3794),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_SL g3822 ( 
.A(n_3812),
.B(n_3785),
.Y(n_3822)
);

AND4x1_ASAP7_75t_L g3823 ( 
.A(n_3816),
.B(n_3769),
.C(n_3765),
.D(n_442),
.Y(n_3823)
);

AOI221xp5_ASAP7_75t_L g3824 ( 
.A1(n_3810),
.A2(n_437),
.B1(n_439),
.B2(n_443),
.C(n_444),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3792),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3795),
.Y(n_3826)
);

OAI322xp33_ASAP7_75t_L g3827 ( 
.A1(n_3810),
.A2(n_443),
.A3(n_444),
.B1(n_445),
.B2(n_446),
.C1(n_448),
.C2(n_449),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3815),
.Y(n_3828)
);

INVx1_ASAP7_75t_L g3829 ( 
.A(n_3799),
.Y(n_3829)
);

AOI22xp5_ASAP7_75t_L g3830 ( 
.A1(n_3814),
.A2(n_445),
.B1(n_446),
.B2(n_448),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3801),
.Y(n_3831)
);

OA22x2_ASAP7_75t_L g3832 ( 
.A1(n_3813),
.A2(n_450),
.B1(n_451),
.B2(n_452),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3813),
.Y(n_3833)
);

NAND2x1_ASAP7_75t_SL g3834 ( 
.A(n_3797),
.B(n_451),
.Y(n_3834)
);

AOI22xp5_ASAP7_75t_L g3835 ( 
.A1(n_3814),
.A2(n_452),
.B1(n_454),
.B2(n_456),
.Y(n_3835)
);

AOI22xp33_ASAP7_75t_L g3836 ( 
.A1(n_3821),
.A2(n_3793),
.B1(n_3797),
.B2(n_3798),
.Y(n_3836)
);

INVxp67_ASAP7_75t_L g3837 ( 
.A(n_3822),
.Y(n_3837)
);

AOI22xp5_ASAP7_75t_L g3838 ( 
.A1(n_3817),
.A2(n_3809),
.B1(n_3808),
.B2(n_3807),
.Y(n_3838)
);

A2O1A1Ixp33_ASAP7_75t_L g3839 ( 
.A1(n_3819),
.A2(n_3800),
.B(n_3805),
.C(n_3802),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3833),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3818),
.Y(n_3841)
);

AOI221xp5_ASAP7_75t_L g3842 ( 
.A1(n_3828),
.A2(n_3798),
.B1(n_3803),
.B2(n_3806),
.C(n_458),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3832),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3825),
.Y(n_3844)
);

AOI31xp33_ASAP7_75t_L g3845 ( 
.A1(n_3820),
.A2(n_3835),
.A3(n_3830),
.B(n_3824),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3826),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3829),
.Y(n_3847)
);

O2A1O1Ixp33_ASAP7_75t_SL g3848 ( 
.A1(n_3823),
.A2(n_3803),
.B(n_456),
.C(n_457),
.Y(n_3848)
);

OAI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3831),
.A2(n_454),
.B1(n_457),
.B2(n_458),
.Y(n_3849)
);

OAI22xp5_ASAP7_75t_L g3850 ( 
.A1(n_3823),
.A2(n_3834),
.B1(n_3827),
.B2(n_462),
.Y(n_3850)
);

OAI211xp5_ASAP7_75t_L g3851 ( 
.A1(n_3817),
.A2(n_459),
.B(n_460),
.C(n_463),
.Y(n_3851)
);

OAI31xp33_ASAP7_75t_L g3852 ( 
.A1(n_3822),
.A2(n_459),
.A3(n_464),
.B(n_465),
.Y(n_3852)
);

AOI22xp5_ASAP7_75t_L g3853 ( 
.A1(n_3837),
.A2(n_464),
.B1(n_466),
.B2(n_467),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3843),
.B(n_466),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_SL g3855 ( 
.A(n_3841),
.B(n_468),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3840),
.Y(n_3856)
);

AOI221xp5_ASAP7_75t_L g3857 ( 
.A1(n_3839),
.A2(n_468),
.B1(n_469),
.B2(n_470),
.C(n_471),
.Y(n_3857)
);

NOR2x1_ASAP7_75t_L g3858 ( 
.A(n_3851),
.B(n_469),
.Y(n_3858)
);

INVxp67_ASAP7_75t_L g3859 ( 
.A(n_3850),
.Y(n_3859)
);

NOR2x1_ASAP7_75t_L g3860 ( 
.A(n_3845),
.B(n_473),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3849),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3836),
.B(n_474),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_SL g3863 ( 
.A(n_3852),
.B(n_475),
.Y(n_3863)
);

AOI221xp5_ASAP7_75t_SL g3864 ( 
.A1(n_3842),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.C(n_479),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3854),
.Y(n_3865)
);

NAND2xp5_ASAP7_75t_L g3866 ( 
.A(n_3859),
.B(n_3838),
.Y(n_3866)
);

AOI22xp5_ASAP7_75t_L g3867 ( 
.A1(n_3857),
.A2(n_3848),
.B1(n_3846),
.B2(n_3844),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3862),
.Y(n_3868)
);

HB1xp67_ASAP7_75t_L g3869 ( 
.A(n_3856),
.Y(n_3869)
);

BUFx2_ASAP7_75t_L g3870 ( 
.A(n_3858),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3853),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3861),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3863),
.Y(n_3873)
);

NOR4xp25_ASAP7_75t_L g3874 ( 
.A(n_3872),
.B(n_3847),
.C(n_3860),
.D(n_3864),
.Y(n_3874)
);

AOI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3871),
.A2(n_3855),
.B1(n_480),
.B2(n_481),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3869),
.Y(n_3876)
);

AOI22xp5_ASAP7_75t_L g3877 ( 
.A1(n_3873),
.A2(n_478),
.B1(n_480),
.B2(n_481),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3870),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3878),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3875),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3876),
.Y(n_3881)
);

INVx1_ASAP7_75t_SL g3882 ( 
.A(n_3877),
.Y(n_3882)
);

BUFx2_ASAP7_75t_L g3883 ( 
.A(n_3874),
.Y(n_3883)
);

INVx1_ASAP7_75t_L g3884 ( 
.A(n_3879),
.Y(n_3884)
);

AO22x1_ASAP7_75t_L g3885 ( 
.A1(n_3883),
.A2(n_3868),
.B1(n_3866),
.B2(n_3865),
.Y(n_3885)
);

INVxp67_ASAP7_75t_L g3886 ( 
.A(n_3881),
.Y(n_3886)
);

OAI22xp5_ASAP7_75t_L g3887 ( 
.A1(n_3882),
.A2(n_3867),
.B1(n_3866),
.B2(n_3880),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3884),
.Y(n_3888)
);

INVx1_ASAP7_75t_L g3889 ( 
.A(n_3887),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3889),
.A2(n_3882),
.B1(n_3886),
.B2(n_3885),
.Y(n_3890)
);

INVx1_ASAP7_75t_L g3891 ( 
.A(n_3890),
.Y(n_3891)
);

OAI22xp33_ASAP7_75t_L g3892 ( 
.A1(n_3891),
.A2(n_3888),
.B1(n_483),
.B2(n_485),
.Y(n_3892)
);

INVx1_ASAP7_75t_L g3893 ( 
.A(n_3892),
.Y(n_3893)
);

AOI221xp5_ASAP7_75t_L g3894 ( 
.A1(n_3893),
.A2(n_482),
.B1(n_483),
.B2(n_485),
.C(n_528),
.Y(n_3894)
);

AOI211xp5_ASAP7_75t_L g3895 ( 
.A1(n_3894),
.A2(n_482),
.B(n_529),
.C(n_530),
.Y(n_3895)
);


endmodule