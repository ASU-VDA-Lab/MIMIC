module fake_ariane_743_n_667 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_143, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_667);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_667;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_663;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_309;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_661;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_212;
wire n_444;
wire n_355;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_484;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

INVx2_ASAP7_75t_SL g145 ( 
.A(n_29),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_43),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_2),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_20),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_61),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_70),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_79),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_59),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_13),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_112),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_42),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_65),
.Y(n_161)
);

BUFx10_ASAP7_75t_L g162 ( 
.A(n_46),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_33),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_6),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_25),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_106),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_23),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_84),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_95),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_100),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_82),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_3),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_10),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_108),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_27),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_40),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_75),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_109),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_56),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_2),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_32),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_17),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_9),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_58),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_99),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_80),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_8),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_137),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_45),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_10),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_98),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_73),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_30),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_15),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_139),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_150),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_151),
.B(n_0),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_157),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_162),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_173),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_184),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_187),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_175),
.B(n_0),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_166),
.B(n_1),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_152),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_181),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_197),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_191),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_3),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_198),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_146),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_204),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_186),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_154),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_203),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_155),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_158),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_218),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_218),
.Y(n_264)
);

AND2x6_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_240),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_232),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_167),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_252),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_167),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

BUFx8_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_228),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_199),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_199),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_242),
.Y(n_292)
);

NAND2xp33_ASAP7_75t_SL g293 ( 
.A(n_238),
.B(n_145),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_258),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_231),
.A2(n_214),
.B(n_206),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_249),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_241),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_261),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_243),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_244),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_247),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_248),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

BUFx8_ASAP7_75t_L g310 ( 
.A(n_215),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_224),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_242),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_222),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_310),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_264),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_270),
.B(n_277),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_264),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_287),
.Y(n_321)
);

NAND2x1p5_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_205),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_289),
.A2(n_205),
.B1(n_163),
.B2(n_209),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_305),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_266),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_267),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_285),
.B(n_211),
.Y(n_334)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_225),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_294),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_269),
.Y(n_338)
);

NOR2x1p5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_159),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_264),
.Y(n_340)
);

AOI21x1_ASAP7_75t_L g341 ( 
.A1(n_270),
.A2(n_210),
.B(n_169),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_284),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_265),
.B(n_213),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_285),
.B(n_171),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_271),
.B(n_160),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_271),
.B(n_172),
.Y(n_346)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_279),
.B(n_193),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_272),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_294),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_L g350 ( 
.A1(n_289),
.A2(n_208),
.B(n_202),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_201),
.B1(n_156),
.B2(n_189),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_286),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_274),
.B(n_161),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_268),
.B(n_168),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_274),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_170),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_R g359 ( 
.A(n_293),
.B(n_178),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_285),
.B(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_313),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_286),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_282),
.Y(n_364)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_302),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_262),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_262),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_278),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_300),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_292),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_277),
.B(n_156),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_281),
.Y(n_374)
);

BUFx4f_ASAP7_75t_L g375 ( 
.A(n_302),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_281),
.Y(n_376)
);

OR2x6_ASAP7_75t_L g377 ( 
.A(n_307),
.B(n_201),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_298),
.B(n_194),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_288),
.B(n_4),
.Y(n_379)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_265),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_291),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_R g382 ( 
.A(n_293),
.B(n_14),
.Y(n_382)
);

AO22x2_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_308),
.B1(n_314),
.B2(n_357),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_337),
.B(n_311),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_316),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_370),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_381),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_329),
.Y(n_388)
);

AO22x2_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_308),
.B1(n_307),
.B2(n_299),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_329),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_321),
.B(n_287),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_372),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_372),
.Y(n_395)
);

AO22x2_ASAP7_75t_L g396 ( 
.A1(n_323),
.A2(n_311),
.B1(n_312),
.B2(n_291),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_361),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

BUFx8_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_323),
.B(n_301),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_287),
.B1(n_303),
.B2(n_265),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g402 ( 
.A(n_371),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

NAND2x1p5_ASAP7_75t_L g404 ( 
.A(n_328),
.B(n_309),
.Y(n_404)
);

AO22x2_ASAP7_75t_L g405 ( 
.A1(n_370),
.A2(n_346),
.B1(n_347),
.B2(n_368),
.Y(n_405)
);

NAND2x1p5_ASAP7_75t_L g406 ( 
.A(n_349),
.B(n_290),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_367),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_333),
.Y(n_408)
);

NAND2x1p5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_295),
.Y(n_409)
);

AO22x2_ASAP7_75t_L g410 ( 
.A1(n_346),
.A2(n_292),
.B1(n_296),
.B2(n_310),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_321),
.B(n_265),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_338),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_348),
.Y(n_413)
);

AO22x2_ASAP7_75t_L g414 ( 
.A1(n_347),
.A2(n_304),
.B1(n_306),
.B2(n_276),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_356),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_362),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_364),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_306),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

OAI221xp5_ASAP7_75t_L g423 ( 
.A1(n_325),
.A2(n_276),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_423)
);

AO22x2_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_276),
.B1(n_265),
.B2(n_297),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_324),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_326),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_374),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_375),
.B(n_297),
.Y(n_430)
);

AO22x2_ASAP7_75t_L g431 ( 
.A1(n_325),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_317),
.Y(n_432)
);

AO22x2_ASAP7_75t_L g433 ( 
.A1(n_379),
.A2(n_11),
.B1(n_12),
.B2(n_156),
.Y(n_433)
);

AO22x2_ASAP7_75t_L g434 ( 
.A1(n_337),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_369),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_369),
.Y(n_436)
);

OAI221xp5_ASAP7_75t_L g437 ( 
.A1(n_322),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.C(n_22),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_352),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_327),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_352),
.B(n_31),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_359),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_334),
.B(n_142),
.Y(n_442)
);

AND2x4_ASAP7_75t_L g443 ( 
.A(n_365),
.B(n_34),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_318),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_319),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_322),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_318),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_365),
.B(n_141),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_334),
.B(n_35),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g450 ( 
.A(n_395),
.B(n_339),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_419),
.B(n_420),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_418),
.B(n_320),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_394),
.B(n_320),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_400),
.B(n_330),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_403),
.B(n_330),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_403),
.B(n_335),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_384),
.B(n_335),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_441),
.B(n_382),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_360),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_385),
.B(n_382),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_386),
.B(n_377),
.Y(n_461)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_439),
.B(n_359),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_377),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_397),
.B(n_355),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_SL g465 ( 
.A(n_393),
.B(n_351),
.Y(n_465)
);

NAND2xp33_ASAP7_75t_SL g466 ( 
.A(n_398),
.B(n_351),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_360),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_SL g468 ( 
.A(n_408),
.B(n_332),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_401),
.B(n_343),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_440),
.B(n_343),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_SL g471 ( 
.A(n_412),
.B(n_413),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_440),
.B(n_350),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_443),
.B(n_344),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_443),
.B(n_344),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_409),
.B(n_399),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_399),
.B(n_380),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_406),
.B(n_380),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_415),
.B(n_416),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_417),
.B(n_380),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_405),
.B(n_340),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_391),
.B(n_380),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_421),
.B(n_341),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_404),
.B(n_442),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_449),
.B(n_373),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_388),
.B(n_373),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_36),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_390),
.B(n_37),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_396),
.B(n_38),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_SL g489 ( 
.A(n_435),
.B(n_39),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_436),
.B(n_44),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_448),
.B(n_47),
.Y(n_491)
);

NAND2xp33_ASAP7_75t_SL g492 ( 
.A(n_425),
.B(n_48),
.Y(n_492)
);

NAND2xp33_ASAP7_75t_SL g493 ( 
.A(n_430),
.B(n_49),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_478),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_459),
.A2(n_433),
.B1(n_434),
.B2(n_431),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_467),
.B(n_387),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_471),
.A2(n_423),
.B(n_428),
.C(n_426),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_464),
.B(n_405),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_484),
.A2(n_411),
.B(n_429),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_437),
.B(n_438),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_474),
.B(n_422),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_457),
.A2(n_407),
.B(n_392),
.Y(n_503)
);

AOI211x1_ASAP7_75t_L g504 ( 
.A1(n_451),
.A2(n_433),
.B(n_431),
.C(n_434),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_482),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_470),
.B(n_427),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_445),
.B(n_432),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_424),
.B(n_383),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_481),
.A2(n_483),
.B(n_490),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_482),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_461),
.Y(n_511)
);

INVx8_ASAP7_75t_L g512 ( 
.A(n_463),
.Y(n_512)
);

O2A1O1Ixp33_ASAP7_75t_SL g513 ( 
.A1(n_454),
.A2(n_424),
.B(n_414),
.C(n_410),
.Y(n_513)
);

OAI21x1_ASAP7_75t_SL g514 ( 
.A1(n_486),
.A2(n_383),
.B(n_389),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_463),
.B(n_389),
.Y(n_515)
);

AOI21x1_ASAP7_75t_L g516 ( 
.A1(n_469),
.A2(n_414),
.B(n_410),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_402),
.Y(n_517)
);

A2O1A1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_492),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_472),
.A2(n_53),
.B(n_54),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_476),
.B(n_455),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_487),
.A2(n_55),
.B(n_57),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_456),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_517),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_512),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

CKINVDCx8_ASAP7_75t_R g527 ( 
.A(n_512),
.Y(n_527)
);

OA21x2_ASAP7_75t_L g528 ( 
.A1(n_522),
.A2(n_479),
.B(n_477),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_506),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_509),
.A2(n_453),
.B(n_452),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_494),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_500),
.A2(n_493),
.B(n_489),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_521),
.A2(n_468),
.B(n_466),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_512),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g536 ( 
.A1(n_497),
.A2(n_460),
.B1(n_450),
.B2(n_462),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_458),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_501),
.A2(n_465),
.B(n_63),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_507),
.A2(n_60),
.B(n_64),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_503),
.A2(n_66),
.B(n_67),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_498),
.A2(n_68),
.B(n_69),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_495),
.A2(n_72),
.B1(n_74),
.B2(n_76),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_508),
.A2(n_77),
.B(n_83),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_497),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_495),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_545)
);

AOI221xp5_ASAP7_75t_SL g546 ( 
.A1(n_523),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.C(n_96),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_502),
.A2(n_97),
.B(n_101),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

AO31x2_ASAP7_75t_L g549 ( 
.A1(n_505),
.A2(n_102),
.A3(n_103),
.B(n_104),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_496),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_531),
.B(n_516),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_550),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_504),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_530),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_526),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_530),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_524),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_528),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_529),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_529),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_548),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_528),
.Y(n_565)
);

CKINVDCx11_ASAP7_75t_R g566 ( 
.A(n_527),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_537),
.B(n_515),
.Y(n_567)
);

AO31x2_ASAP7_75t_L g568 ( 
.A1(n_538),
.A2(n_518),
.A3(n_510),
.B(n_514),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_528),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_535),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_534),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_525),
.B(n_520),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_549),
.Y(n_573)
);

AOI21x1_ASAP7_75t_L g574 ( 
.A1(n_534),
.A2(n_513),
.B(n_519),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_533),
.A2(n_105),
.B(n_107),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_549),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_541),
.A2(n_140),
.B(n_113),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

NAND2x1p5_ASAP7_75t_L g579 ( 
.A(n_535),
.B(n_110),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_536),
.B(n_117),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_543),
.Y(n_581)
);

NAND2x1p5_ASAP7_75t_L g582 ( 
.A(n_543),
.B(n_119),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_566),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_R g584 ( 
.A(n_566),
.B(n_545),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_572),
.B(n_545),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_555),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_558),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_R g588 ( 
.A(n_557),
.B(n_547),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_560),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_R g590 ( 
.A(n_561),
.B(n_539),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_567),
.B(n_542),
.Y(n_591)
);

CKINVDCx11_ASAP7_75t_R g592 ( 
.A(n_564),
.Y(n_592)
);

NOR2x1_ASAP7_75t_L g593 ( 
.A(n_580),
.B(n_544),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_553),
.B(n_542),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_552),
.B(n_570),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_562),
.B(n_122),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_551),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_551),
.Y(n_598)
);

NAND2xp33_ASAP7_75t_R g599 ( 
.A(n_565),
.B(n_539),
.Y(n_599)
);

CKINVDCx8_ASAP7_75t_R g600 ( 
.A(n_570),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_559),
.B(n_540),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_559),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_R g603 ( 
.A(n_577),
.B(n_124),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_581),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_554),
.B(n_546),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_595),
.B(n_569),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_597),
.B(n_569),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_556),
.Y(n_608)
);

AOI22xp33_ASAP7_75t_L g609 ( 
.A1(n_585),
.A2(n_563),
.B1(n_578),
.B2(n_576),
.Y(n_609)
);

BUFx2_ASAP7_75t_SL g610 ( 
.A(n_600),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_586),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_602),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_584),
.A2(n_563),
.B1(n_573),
.B2(n_582),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_601),
.B(n_554),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_601),
.B(n_556),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_554),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_590),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g619 ( 
.A(n_589),
.B(n_556),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_593),
.B(n_574),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_612),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_611),
.Y(n_622)
);

INVx5_ASAP7_75t_SL g623 ( 
.A(n_615),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_614),
.B(n_571),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_606),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_618),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_616),
.Y(n_627)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_613),
.A2(n_594),
.B1(n_591),
.B2(n_596),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_607),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_626),
.B(n_615),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_623),
.B(n_614),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_622),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_623),
.B(n_615),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_624),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_621),
.B(n_608),
.Y(n_635)
);

OAI31xp33_ASAP7_75t_SL g636 ( 
.A1(n_630),
.A2(n_620),
.A3(n_628),
.B(n_624),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_630),
.B(n_583),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_632),
.A2(n_603),
.B1(n_620),
.B2(n_592),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_629),
.B(n_627),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_635),
.B(n_608),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_637),
.B(n_634),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_639),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_636),
.B(n_634),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_640),
.B(n_619),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_638),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_644),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_645),
.B(n_610),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_642),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_646),
.B(n_643),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_648),
.B(n_641),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_649),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_650),
.C(n_647),
.Y(n_652)
);

AOI221xp5_ASAP7_75t_L g653 ( 
.A1(n_652),
.A2(n_605),
.B1(n_609),
.B2(n_582),
.C(n_617),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_579),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_654),
.B(n_631),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g656 ( 
.A(n_655),
.B(n_579),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_656),
.Y(n_657)
);

OAI22x1_ASAP7_75t_L g658 ( 
.A1(n_657),
.A2(n_633),
.B1(n_575),
.B2(n_617),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_658),
.A2(n_604),
.B1(n_619),
.B2(n_571),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_659),
.B(n_125),
.Y(n_660)
);

AOI22xp33_ASAP7_75t_L g661 ( 
.A1(n_659),
.A2(n_571),
.B1(n_588),
.B2(n_533),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_660),
.A2(n_599),
.B1(n_568),
.B2(n_129),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_661),
.A2(n_126),
.B(n_127),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_663),
.Y(n_664)
);

INVxp33_ASAP7_75t_L g665 ( 
.A(n_662),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_664),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.C(n_138),
.Y(n_666)
);

OAI31xp33_ASAP7_75t_L g667 ( 
.A1(n_666),
.A2(n_568),
.A3(n_665),
.B(n_657),
.Y(n_667)
);


endmodule