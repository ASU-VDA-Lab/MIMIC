module fake_jpeg_13742_n_94 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_31),
.Y(n_39)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_12),
.B(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_15),
.Y(n_35)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_30),
.Y(n_34)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_14),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_17),
.B1(n_30),
.B2(n_22),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_24),
.A2(n_22),
.B1(n_21),
.B2(n_20),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_13),
.B1(n_16),
.B2(n_11),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_25),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_25),
.B1(n_31),
.B2(n_28),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

A2O1A1O1Ixp25_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_25),
.B(n_23),
.C(n_14),
.D(n_16),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_33),
.B(n_40),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_30),
.C(n_23),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_34),
.C(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_52),
.B1(n_29),
.B2(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_50),
.B1(n_52),
.B2(n_46),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_41),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_51),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_65),
.Y(n_75)
);

AO21x1_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_57),
.B(n_58),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_71),
.C(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_45),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_13),
.C(n_11),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_74),
.B1(n_29),
.B2(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_73),
.B(n_78),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_60),
.B1(n_61),
.B2(n_27),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_71),
.C(n_60),
.Y(n_79)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_10),
.B1(n_9),
.B2(n_7),
.C(n_8),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_74),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_76),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_89),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_83),
.C(n_7),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_8),
.B(n_9),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_2),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_91),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_2),
.Y(n_94)
);


endmodule