module fake_ibex_827_n_16 (n_1, n_4, n_3, n_6, n_5, n_2, n_0, n_16);

input n_1;
input n_4;
input n_3;
input n_6;
input n_5;
input n_2;
input n_0;

output n_16;


SDFHx2_ASAP7_75t_R g7 ( 
.CLK(n_1),
.D(n_5),
.SE(n_2),
.SI(n_0),
.QN(n_7)
);


endmodule