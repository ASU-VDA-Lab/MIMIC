module real_jpeg_4728_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_400;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_1),
.A2(n_147),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_1),
.A2(n_158),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_1),
.A2(n_118),
.B1(n_125),
.B2(n_158),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_1),
.A2(n_158),
.B1(n_361),
.B2(n_362),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_3),
.A2(n_238),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_3),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_3),
.A2(n_261),
.B1(n_269),
.B2(n_276),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_3),
.A2(n_276),
.B1(n_350),
.B2(n_352),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_3),
.A2(n_276),
.B1(n_430),
.B2(n_432),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_4),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_4),
.A2(n_93),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_4),
.A2(n_93),
.B1(n_262),
.B2(n_271),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_4),
.A2(n_58),
.B1(n_93),
.B2(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_5),
.A2(n_34),
.B1(n_35),
.B2(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_34),
.B1(n_50),
.B2(n_53),
.Y(n_173)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_7),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_7),
.Y(n_303)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_7),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_8),
.A2(n_46),
.B1(n_160),
.B2(n_165),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_8),
.A2(n_46),
.B1(n_269),
.B2(n_390),
.Y(n_389)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_9),
.Y(n_109)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_11),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g384 ( 
.A(n_11),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_11),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_12),
.A2(n_112),
.B1(n_113),
.B2(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_12),
.A2(n_54),
.B1(n_112),
.B2(n_245),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_112),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_12),
.A2(n_112),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_13),
.A2(n_113),
.B1(n_114),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_13),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_13),
.A2(n_203),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_13),
.A2(n_203),
.B1(n_238),
.B2(n_315),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_13),
.A2(n_203),
.B1(n_404),
.B2(n_406),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_14),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_14),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_14),
.A2(n_40),
.B1(n_80),
.B2(n_179),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_14),
.A2(n_80),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_16),
.A2(n_238),
.B1(n_239),
.B2(n_242),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_16),
.B(n_251),
.C(n_254),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_16),
.B(n_149),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_16),
.B(n_183),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_16),
.B(n_87),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_16),
.B(n_321),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_228),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_226),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_205),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_20),
.B(n_205),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_130),
.C(n_175),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_21),
.A2(n_22),
.B1(n_130),
.B2(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_88),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_23),
.A2(n_24),
.B(n_90),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_44),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_24),
.A2(n_89),
.B1(n_90),
.B2(n_129),
.Y(n_88)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_24),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_24),
.A2(n_44),
.B1(n_129),
.B2(n_418),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_33),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_25),
.A2(n_33),
.B1(n_178),
.B2(n_181),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_25),
.A2(n_260),
.B(n_266),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_25),
.A2(n_242),
.B(n_266),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_25),
.A2(n_334),
.B1(n_387),
.B2(n_388),
.Y(n_386)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_26),
.B(n_268),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_26),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_26),
.A2(n_333),
.B1(n_360),
.B2(n_365),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_26),
.A2(n_389),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_31),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g270 ( 
.A(n_38),
.Y(n_270)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_38),
.Y(n_391)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_39),
.Y(n_261)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_42),
.Y(n_257)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_42),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_44),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_56),
.B1(n_79),
.B2(n_87),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_45),
.A2(n_56),
.B1(n_87),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g149 ( 
.A1(n_50),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_51),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_51),
.Y(n_238)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_51),
.Y(n_247)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_52),
.Y(n_277)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_56),
.A2(n_79),
.B1(n_87),
.B2(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_56),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_56),
.B(n_244),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_70),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_63),
.B2(n_67),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_69),
.Y(n_151)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_69),
.Y(n_409)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_70),
.A2(n_275),
.B(n_278),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_78),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_72),
.Y(n_253)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_75),
.Y(n_288)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_77),
.Y(n_364)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_84),
.Y(n_241)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_87),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_87),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_110),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_99),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_92),
.Y(n_210)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_122),
.B1(n_125),
.B2(n_127),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_99),
.B(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_100),
.B(n_242),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_100),
.A2(n_201),
.B1(n_202),
.B2(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_108),
.Y(n_100)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_102),
.Y(n_405)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_103),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_104),
.Y(n_377)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_105),
.Y(n_148)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g336 ( 
.A(n_107),
.Y(n_336)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_110),
.A2(n_211),
.B(n_429),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_118),
.Y(n_433)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_119),
.Y(n_431)
);

INVx2_ASAP7_75t_SL g201 ( 
.A(n_120),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_120),
.A2(n_398),
.B(n_400),
.Y(n_397)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g376 ( 
.A1(n_125),
.A2(n_377),
.A3(n_378),
.B1(n_379),
.B2(n_381),
.Y(n_376)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_127),
.Y(n_378)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_128),
.Y(n_380)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_130),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_170),
.B(n_174),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_171),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_149),
.B1(n_154),
.B2(n_159),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_133),
.A2(n_318),
.B(n_324),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_133),
.B(n_356),
.Y(n_355)
);

AOI22x1_ASAP7_75t_L g434 ( 
.A1(n_133),
.A2(n_149),
.B1(n_356),
.B2(n_435),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_133),
.A2(n_324),
.B(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_134),
.A2(n_155),
.B1(n_194),
.B2(n_199),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_134),
.A2(n_199),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_134),
.A2(n_199),
.B1(n_349),
.B2(n_403),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_149),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_141),
.B1(n_142),
.B2(n_146),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_140),
.Y(n_145)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_146),
.B(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_147),
.A2(n_242),
.B(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_148),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_149),
.Y(n_199)
);

AOI32xp33_ASAP7_75t_L g335 ( 
.A1(n_152),
.A2(n_238),
.A3(n_320),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_153),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_157),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_169),
.Y(n_323)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_169),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_174),
.B(n_206),
.CI(n_207),
.CON(n_205),
.SN(n_205)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_175),
.B(n_437),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_193),
.C(n_200),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_176),
.B(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_177),
.B(n_184),
.Y(n_445)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_178),
.Y(n_424)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_185),
.Y(n_422)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_193),
.B(n_200),
.Y(n_416)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_194),
.Y(n_435)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_198),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_199),
.B(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_199),
.A2(n_349),
.B(n_355),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B(n_204),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_201),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_209)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_204),
.Y(n_400)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_205),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_225),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_224),
.Y(n_213)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_237),
.B(n_243),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_215),
.A2(n_216),
.B1(n_275),
.B2(n_314),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_215),
.A2(n_243),
.B(n_314),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_215),
.A2(n_216),
.B1(n_408),
.B2(n_422),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_216),
.A2(n_278),
.B(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI311xp33_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_412),
.A3(n_453),
.B1(n_471),
.C1(n_472),
.Y(n_229)
);

AOI21x1_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_370),
.B(n_411),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_340),
.B(n_369),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_308),
.B(n_339),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_281),
.B(n_307),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_258),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_235),
.B(n_258),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_248),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_236),
.A2(n_248),
.B1(n_249),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_236),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_242),
.B(n_382),
.Y(n_381)
);

OAI21xp33_ASAP7_75t_SL g398 ( 
.A1(n_242),
.A2(n_381),
.B(n_399),
.Y(n_398)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_246),
.Y(n_315)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_257),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_272),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_273),
.C(n_280),
.Y(n_309)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_260),
.Y(n_301)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_271),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_279),
.B2(n_280),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g337 ( 
.A(n_277),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_298),
.B(n_306),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_291),
.B(n_297),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_296),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B(n_295),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_332),
.B(n_334),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_299),
.B(n_304),
.Y(n_306)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_302),
.Y(n_334)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_310),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_330),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_316),
.B2(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_316),
.C(n_330),
.Y(n_341)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_335),
.Y(n_346)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_342),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_347),
.B2(n_368),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_346),
.C(n_368),
.Y(n_371)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_357),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_358),
.C(n_359),
.Y(n_392)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_350),
.Y(n_406)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_360),
.Y(n_387)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_371),
.B(n_372),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_395),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_373)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_385),
.B2(n_386),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_385),
.Y(n_449)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_392),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_392),
.B(n_393),
.C(n_395),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_397),
.B1(n_401),
.B2(n_410),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_402),
.C(n_407),
.Y(n_462)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_401),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_407),
.Y(n_401)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_403),
.Y(n_451)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_439),
.Y(n_412)
);

A2O1A1Ixp33_ASAP7_75t_SL g472 ( 
.A1(n_413),
.A2(n_439),
.B(n_473),
.C(n_476),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_436),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_436),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_417),
.C(n_419),
.Y(n_414)
);

FAx1_ASAP7_75t_SL g452 ( 
.A(n_415),
.B(n_417),
.CI(n_419),
.CON(n_452),
.SN(n_452)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_427),
.C(n_434),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_423),
.Y(n_461)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_427),
.A2(n_428),
.B1(n_434),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_434),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_452),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_452),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_445),
.C(n_446),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_441),
.A2(n_442),
.B1(n_445),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_445),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.C(n_450),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_447),
.A2(n_448),
.B1(n_450),
.B2(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_450),
.Y(n_459)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_452),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_466),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_455),
.A2(n_474),
.B(n_475),
.Y(n_473)
);

NOR2x1_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_463),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_463),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_460),
.C(n_462),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_469),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_460),
.A2(n_461),
.B1(n_462),
.B2(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_468),
.Y(n_474)
);


endmodule