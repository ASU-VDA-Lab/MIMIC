module fake_jpeg_9960_n_261 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_261);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_261;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_23),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_43),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_33),
.B1(n_37),
.B2(n_35),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_37),
.B1(n_15),
.B2(n_26),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_22),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_26),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_15),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_48),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_56),
.Y(n_86)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_71),
.B1(n_73),
.B2(n_51),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_19),
.B1(n_18),
.B2(n_26),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_21),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_63),
.Y(n_78)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_68),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_30),
.C(n_29),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_46),
.C(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_41),
.B(n_25),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_39),
.B1(n_52),
.B2(n_53),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_84),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_44),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_21),
.B(n_13),
.C(n_19),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_63),
.A2(n_53),
.B1(n_45),
.B2(n_49),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_53),
.B1(n_71),
.B2(n_73),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_90),
.A2(n_72),
.B1(n_45),
.B2(n_59),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_43),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_100),
.B1(n_110),
.B2(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_101),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_55),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_98),
.A2(n_62),
.B(n_19),
.Y(n_133)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_107),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_75),
.A2(n_51),
.B1(n_70),
.B2(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_113),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_90),
.A2(n_81),
.B(n_85),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_109),
.B(n_91),
.Y(n_121)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_57),
.B(n_70),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_114),
.Y(n_118)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_109),
.B(n_103),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_133),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_108),
.A2(n_81),
.B1(n_83),
.B2(n_74),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_100),
.B1(n_97),
.B2(n_110),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_78),
.C(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_122),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_47),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_101),
.A3(n_95),
.B1(n_113),
.B2(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_51),
.B1(n_92),
.B2(n_50),
.Y(n_127)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_64),
.A3(n_62),
.B1(n_77),
.B2(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_103),
.A2(n_80),
.B1(n_92),
.B2(n_77),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_76),
.B1(n_86),
.B2(n_29),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_136),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_80),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_137),
.A2(n_118),
.B1(n_127),
.B2(n_18),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_104),
.C(n_112),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_153),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_100),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_127),
.B1(n_133),
.B2(n_116),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_152),
.B1(n_145),
.B2(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_17),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_150),
.B(n_155),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_86),
.B1(n_23),
.B2(n_18),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_151),
.A2(n_122),
.B1(n_124),
.B2(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_27),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_157),
.B(n_159),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_136),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_180),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_115),
.B(n_121),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_165),
.B(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_162),
.B(n_164),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_126),
.B(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_168),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_119),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_171),
.B(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_138),
.B(n_125),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_142),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_179),
.B(n_149),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_145),
.B1(n_152),
.B2(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_144),
.B1(n_154),
.B2(n_23),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_148),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_181),
.B(n_183),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_170),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_168),
.Y(n_201)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_69),
.Y(n_212)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_170),
.B(n_154),
.C(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_197),
.C(n_162),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_194),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_117),
.B1(n_13),
.B2(n_21),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_176),
.B1(n_173),
.B2(n_27),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_69),
.C(n_30),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_165),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_182),
.Y(n_213)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_200),
.B(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_212),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_203),
.C(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_178),
.C(n_166),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_186),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_69),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_184),
.B1(n_191),
.B2(n_194),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_220),
.B1(n_13),
.B2(n_8),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_207),
.B1(n_203),
.B2(n_210),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_195),
.Y(n_226)
);

NOR3xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_189),
.C(n_197),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_9),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_223),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_185),
.C(n_187),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_198),
.C(n_17),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_232),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_234),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_235),
.C(n_221),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_215),
.B(n_0),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_60),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_60),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_219),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_32),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_236),
.A2(n_214),
.B(n_216),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_230),
.B(n_229),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_244),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_218),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_245),
.B(n_249),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_250),
.B(n_238),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_239),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_243),
.A2(n_235),
.B(n_230),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_238),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_251),
.A2(n_252),
.B(n_253),
.Y(n_254)
);

AOI322xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_255),
.A3(n_6),
.B1(n_12),
.B2(n_11),
.C1(n_10),
.C2(n_8),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_253),
.A2(n_248),
.B(n_227),
.Y(n_255)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_6),
.B(n_12),
.C(n_11),
.D(n_10),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g258 ( 
.A1(n_257),
.A2(n_10),
.A3(n_8),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_1),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_0),
.C(n_1),
.Y(n_259)
);

AOI221xp5_ASAP7_75t_L g260 ( 
.A1(n_259),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.C(n_50),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_50),
.Y(n_261)
);


endmodule