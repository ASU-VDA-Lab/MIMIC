module fake_jpeg_31885_n_454 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_454);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_454;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_4),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_15),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_49),
.B(n_41),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_19),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_53),
.B(n_72),
.Y(n_104)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_64),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_91),
.Y(n_127)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_37),
.B(n_15),
.Y(n_84)
);

OR2x2_ASAP7_75t_SL g146 ( 
.A(n_84),
.B(n_25),
.Y(n_146)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_17),
.B(n_0),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_65),
.A2(n_39),
.B1(n_46),
.B2(n_27),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_96),
.A2(n_53),
.B1(n_68),
.B2(n_71),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_41),
.B1(n_44),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_108),
.A2(n_145),
.B1(n_77),
.B2(n_76),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_111),
.B(n_38),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_113),
.A2(n_44),
.B1(n_30),
.B2(n_28),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_49),
.B(n_27),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_139),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_146),
.Y(n_165)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_72),
.B(n_17),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_60),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_52),
.A2(n_25),
.B1(n_42),
.B2(n_38),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_32),
.B(n_18),
.C(n_20),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_150),
.B(n_154),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_121),
.A2(n_57),
.B1(n_80),
.B2(n_29),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_178),
.B1(n_195),
.B2(n_124),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_152),
.B(n_177),
.Y(n_199)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_100),
.Y(n_153)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_156),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_157),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_61),
.B1(n_59),
.B2(n_62),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_158),
.A2(n_188),
.B1(n_192),
.B2(n_117),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_63),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_159),
.A2(n_191),
.B1(n_97),
.B2(n_140),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_18),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_161),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_51),
.Y(n_161)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_162),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_125),
.B(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_171),
.Y(n_210)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_164),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_42),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_167),
.B(n_173),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_26),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_168),
.B(n_169),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_26),
.Y(n_169)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_113),
.B(n_16),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_134),
.Y(n_174)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_30),
.B1(n_28),
.B2(n_44),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_179),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_105),
.Y(n_180)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_182),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_120),
.B(n_136),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_183),
.B(n_184),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_44),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_113),
.B(n_90),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_193),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_148),
.B(n_132),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_72),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_196),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_131),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_99),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_102),
.A2(n_44),
.B1(n_30),
.B2(n_5),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_116),
.B(n_142),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_114),
.A2(n_30),
.B1(n_3),
.B2(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_109),
.B(n_1),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_197),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_198),
.A2(n_158),
.B1(n_192),
.B2(n_190),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_138),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_225),
.C(n_229),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_202),
.A2(n_157),
.B1(n_194),
.B2(n_175),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_214),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_155),
.B(n_114),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_218),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_130),
.B1(n_119),
.B2(n_117),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_220),
.A2(n_223),
.B1(n_181),
.B2(n_194),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_161),
.A2(n_112),
.B1(n_97),
.B2(n_140),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_222),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_185),
.A2(n_130),
.B1(n_119),
.B2(n_95),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_152),
.B(n_112),
.C(n_95),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_165),
.B(n_147),
.C(n_3),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_171),
.B(n_1),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_196),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_149),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_237),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_161),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_236),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_160),
.B(n_3),
.Y(n_237)
);

INVx11_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_239),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_240),
.B(n_247),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_161),
.B(n_193),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_241),
.A2(n_242),
.B(n_254),
.Y(n_286)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_222),
.A2(n_191),
.B1(n_150),
.B2(n_173),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_165),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_225),
.C(n_222),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_199),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_163),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_248),
.B(n_256),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_182),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_252),
.B(n_266),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_191),
.B(n_193),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_255),
.A2(n_264),
.B1(n_202),
.B2(n_220),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_191),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_213),
.A2(n_186),
.B(n_189),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_257),
.A2(n_265),
.B(n_268),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_274),
.B1(n_224),
.B2(n_157),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_201),
.B(n_159),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_176),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_263),
.B(n_267),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_153),
.B1(n_172),
.B2(n_164),
.Y(n_264)
);

AOI22x1_ASAP7_75t_SL g265 ( 
.A1(n_222),
.A2(n_159),
.B1(n_166),
.B2(n_197),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_205),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_174),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_207),
.A2(n_166),
.B(n_156),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_200),
.Y(n_271)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_271),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_179),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_216),
.B(n_170),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_208),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_277),
.A2(n_255),
.B1(n_264),
.B2(n_268),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_217),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_278),
.B(n_279),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_209),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_296),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_284),
.A2(n_274),
.B1(n_250),
.B2(n_258),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_234),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_287),
.B(n_293),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_251),
.A2(n_223),
.B1(n_224),
.B2(n_234),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_301),
.B1(n_277),
.B2(n_306),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_208),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_289),
.B(n_300),
.C(n_304),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_256),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_226),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_259),
.B(n_227),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_275),
.B(n_232),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_232),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_231),
.C(n_212),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_251),
.A2(n_231),
.B1(n_212),
.B2(n_204),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_162),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_248),
.B(n_204),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_245),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_311),
.B(n_290),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_319),
.B1(n_321),
.B2(n_334),
.Y(n_348)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_276),
.Y(n_315)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_257),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_322),
.C(n_304),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_295),
.A2(n_265),
.B(n_241),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_318),
.A2(n_281),
.B(n_308),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_282),
.A2(n_250),
.B1(n_242),
.B2(n_254),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_246),
.Y(n_322)
);

AOI21xp33_ASAP7_75t_SL g323 ( 
.A1(n_307),
.A2(n_242),
.B(n_273),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_325),
.Y(n_340)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_276),
.Y(n_324)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_324),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_296),
.B(n_289),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_327),
.B(n_200),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_288),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_328),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_329),
.A2(n_284),
.B1(n_295),
.B2(n_300),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_302),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_331),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_273),
.B1(n_263),
.B2(n_267),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_294),
.B1(n_299),
.B2(n_280),
.Y(n_343)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_280),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_292),
.A2(n_240),
.B1(n_270),
.B2(n_262),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_292),
.A2(n_260),
.B1(n_261),
.B2(n_269),
.Y(n_335)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_302),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_336),
.B(n_337),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_294),
.B(n_271),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_338),
.A2(n_362),
.B1(n_315),
.B2(n_239),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_351),
.Y(n_364)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_309),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_363),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_329),
.A2(n_281),
.B1(n_299),
.B2(n_286),
.Y(n_345)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

XOR2x2_ASAP7_75t_L g349 ( 
.A(n_317),
.B(n_286),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_350),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_353),
.B(n_355),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_320),
.B(n_177),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_316),
.A2(n_283),
.B1(n_291),
.B2(n_261),
.Y(n_356)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_356),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_203),
.C(n_283),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_327),
.C(n_326),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_322),
.B(n_203),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_215),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_330),
.A2(n_328),
.B1(n_313),
.B2(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_361),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_337),
.A2(n_321),
.B1(n_318),
.B2(n_311),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_312),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_357),
.B(n_334),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_366),
.B(n_351),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_367),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_348),
.A2(n_328),
.B1(n_336),
.B2(n_312),
.Y(n_370)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_375),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_355),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_326),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_376),
.B(n_377),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_335),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_348),
.A2(n_319),
.B1(n_324),
.B2(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_379),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_381),
.A2(n_383),
.B1(n_360),
.B2(n_342),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_269),
.Y(n_382)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_215),
.B1(n_7),
.B2(n_9),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_339),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_354),
.Y(n_386)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_354),
.Y(n_387)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_371),
.A2(n_360),
.B1(n_344),
.B2(n_349),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_389),
.B(n_398),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_399),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_373),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_396),
.Y(n_411)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_373),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_381),
.A2(n_365),
.B1(n_383),
.B2(n_344),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_401),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g402 ( 
.A1(n_377),
.A2(n_342),
.B(n_352),
.Y(n_402)
);

OAI21x1_ASAP7_75t_SL g406 ( 
.A1(n_402),
.A2(n_372),
.B(n_364),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_374),
.C(n_376),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_408),
.C(n_414),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_412),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_384),
.C(n_364),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_380),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_409),
.B(n_413),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_395),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_380),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_393),
.B(n_375),
.C(n_369),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_369),
.C(n_350),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_387),
.C(n_396),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_410),
.A2(n_388),
.B1(n_390),
.B2(n_394),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_423),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_416),
.B(n_408),
.C(n_414),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_419),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_399),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_403),
.A2(n_415),
.B(n_411),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_421),
.A2(n_352),
.B(n_346),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_404),
.B(n_400),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_424),
.B(n_425),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_405),
.B(n_402),
.C(n_346),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_407),
.B(n_402),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_428),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_386),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_430),
.B(n_437),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g431 ( 
.A(n_426),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_428),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_398),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_433),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_427),
.A2(n_341),
.B(n_11),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_435),
.A2(n_6),
.B(n_11),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_419),
.A2(n_6),
.B1(n_11),
.B2(n_12),
.Y(n_437)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_439),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g445 ( 
.A1(n_440),
.A2(n_435),
.B(n_432),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_429),
.B(n_424),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_442),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_434),
.B(n_422),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_420),
.Y(n_449)
);

OAI321xp33_ASAP7_75t_L g447 ( 
.A1(n_438),
.A2(n_436),
.A3(n_437),
.B1(n_434),
.B2(n_418),
.C(n_422),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_447),
.B(n_443),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_448),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_450),
.A2(n_446),
.B(n_444),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_451),
.B(n_449),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_452),
.A2(n_13),
.B1(n_450),
.B2(n_446),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_13),
.Y(n_454)
);


endmodule