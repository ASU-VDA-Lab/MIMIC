module real_jpeg_21903_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_323, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_323;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_0),
.A2(n_51),
.B1(n_60),
.B2(n_61),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_69),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_1),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_69),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_2),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_2),
.B(n_34),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_2),
.A2(n_57),
.B(n_60),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_117),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_2),
.A2(n_97),
.B1(n_98),
.B2(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_2),
.B(n_42),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_2),
.A2(n_36),
.B(n_207),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_3),
.A2(n_60),
.B1(n_61),
.B2(n_114),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_44),
.B1(n_45),
.B2(n_114),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_253)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_5),
.Y(n_98)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_5),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_6),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_82),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_82),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_82),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_7),
.A2(n_39),
.B1(n_60),
.B2(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_7),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_8),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_10),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_108),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_108),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_108),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_12),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_119),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_119),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_13),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_13),
.A2(n_60),
.B1(n_61),
.B2(n_112),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_112),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_14),
.A2(n_36),
.A3(n_45),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_SL g45 ( 
.A(n_17),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_87),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_22),
.B(n_72),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_27),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_32),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_29),
.B(n_117),
.CON(n_116),
.SN(n_116)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_31),
.A2(n_34),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_31),
.A2(n_34),
.B1(n_81),
.B2(n_298),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_32),
.B(n_36),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_33),
.A2(n_35),
.B1(n_116),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_43),
.B(n_46),
.C(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_46),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_35),
.B(n_117),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_50),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_47),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_42),
.A2(n_47),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_42),
.A2(n_47),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_43),
.A2(n_48),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_43),
.A2(n_48),
.B1(n_113),
.B2(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_43),
.A2(n_48),
.B1(n_146),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_43),
.A2(n_48),
.B1(n_127),
.B2(n_255),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_43),
.A2(n_48),
.B1(n_86),
.B2(n_291),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_45),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_44),
.B(n_46),
.Y(n_202)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_45),
.A2(n_58),
.B(n_117),
.C(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.C(n_65),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_63),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_54),
.A2(n_78),
.B1(n_84),
.B2(n_307),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_59),
.B(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_55),
.A2(n_59),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_59),
.B1(n_102),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_55),
.A2(n_59),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_55),
.A2(n_59),
.B1(n_172),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_55),
.A2(n_59),
.B1(n_192),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_55),
.A2(n_59),
.B1(n_107),
.B2(n_210),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_55),
.A2(n_59),
.B1(n_103),
.B2(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_55),
.A2(n_59),
.B1(n_246),
.B2(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_55),
.A2(n_59),
.B1(n_62),
.B2(n_279),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

CKINVDCx9p33_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_59),
.B(n_117),
.Y(n_177)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_61),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_66),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_67),
.A2(n_68),
.B1(n_70),
.B2(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_67),
.A2(n_70),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_67),
.A2(n_70),
.B1(n_125),
.B2(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_67),
.A2(n_70),
.B1(n_253),
.B2(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_79),
.C(n_83),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_309),
.Y(n_313)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_79),
.C(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_79),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_79),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_83),
.B(n_313),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_84),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI321xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_302),
.A3(n_314),
.B1(n_320),
.B2(n_321),
.C(n_323),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_283),
.B(n_301),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_259),
.B(n_282),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_152),
.B(n_235),
.C(n_258),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_137),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_93),
.B(n_137),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_120),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_104),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_95),
.B(n_104),
.C(n_120),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_96),
.B(n_101),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_97),
.A2(n_99),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_97),
.A2(n_98),
.B1(n_133),
.B2(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_97),
.A2(n_134),
.B1(n_162),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_97),
.A2(n_98),
.B1(n_164),
.B2(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_97),
.A2(n_134),
.B1(n_151),
.B2(n_194),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_97),
.A2(n_100),
.B1(n_134),
.B2(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_97),
.A2(n_134),
.B(n_244),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_98),
.B(n_117),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_115),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_115),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_118),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_128),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_122),
.B(n_128),
.C(n_129),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_126),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_132),
.Y(n_141)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_159)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_142),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_138),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_144),
.B(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_148),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_234),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_229),
.B(n_233),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_215),
.B(n_228),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_196),
.B(n_214),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_184),
.B(n_195),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_173),
.B(n_183),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_165),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_178),
.B(n_182),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_177),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_186),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_198),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_204),
.B1(n_212),
.B2(n_213),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_199),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_201),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_217),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_225),
.C(n_226),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_224),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_225),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_230),
.B(n_231),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_236),
.B(n_237),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_257),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_238),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_247),
.B2(n_248),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_248),
.C(n_257),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_245),
.Y(n_265)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_251),
.C(n_256),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_256),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_254),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_260),
.B(n_261),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_281),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_274),
.B2(n_275),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_275),
.C(n_281),
.Y(n_284)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_267),
.C(n_271),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_269),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_273),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_277),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_278),
.Y(n_294)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_277),
.A2(n_294),
.B(n_297),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_285),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_299),
.B2(n_300),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_293),
.C(n_300),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_304),
.C(n_310),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_292),
.A2(n_304),
.B1(n_305),
.B2(n_319),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_292),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_312),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_306),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_310),
.A2(n_311),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);


endmodule