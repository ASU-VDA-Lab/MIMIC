module fake_netlist_5_1653_n_786 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_786);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_786;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_629;
wire n_590;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_607;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_163;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_273;
wire n_161;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_728;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_SL g154 ( 
.A(n_85),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_2),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_6),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_79),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_46),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_150),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_59),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_52),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_39),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_102),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_127),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_36),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_94),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_67),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_28),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_6),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_15),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_12),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_74),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_73),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_17),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_117),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_38),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_141),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_143),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_34),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_98),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_50),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_44),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_136),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_13),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_130),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_90),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_65),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_27),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_149),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_47),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_75),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_97),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_119),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_71),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_0),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_164),
.B(n_18),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g214 ( 
.A(n_164),
.B(n_19),
.Y(n_214)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_208),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_156),
.B(n_174),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

BUFx8_ASAP7_75t_SL g226 ( 
.A(n_185),
.Y(n_226)
);

BUFx8_ASAP7_75t_SL g227 ( 
.A(n_189),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_158),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_20),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_176),
.B(n_3),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_176),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_179),
.B(n_4),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_179),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

OAI22x1_ASAP7_75t_R g240 ( 
.A1(n_193),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_201),
.Y(n_241)
);

OAI22x1_ASAP7_75t_L g242 ( 
.A1(n_192),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_177),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_207),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_154),
.B(n_21),
.Y(n_247)
);

NAND2x1p5_ASAP7_75t_L g248 ( 
.A(n_191),
.B(n_22),
.Y(n_248)
);

OAI21x1_ASAP7_75t_L g249 ( 
.A1(n_180),
.A2(n_9),
.B(n_10),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_180),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_180),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

CKINVDCx6p67_ASAP7_75t_R g254 ( 
.A(n_209),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_226),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_229),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_227),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_223),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_222),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_225),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_225),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_217),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_215),
.Y(n_265)
);

NOR2xp67_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_157),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

BUFx2_ASAP7_75t_SL g268 ( 
.A(n_213),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_217),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_215),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_217),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_219),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_219),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_219),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_210),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_215),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_234),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_211),
.B(n_199),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_228),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_234),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_228),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_251),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_232),
.B(n_159),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_238),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_251),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_243),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_243),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_231),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_233),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_257),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_213),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_239),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_267),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_276),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_260),
.B(n_214),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_285),
.B(n_214),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_237),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_282),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_268),
.B(n_266),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_214),
.Y(n_311)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_236),
.C(n_235),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_230),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_269),
.B(n_248),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_230),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_261),
.B(n_230),
.C(n_221),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_239),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_288),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_270),
.B(n_239),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_287),
.B(n_272),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_274),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_243),
.Y(n_324)
);

AND2x6_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_247),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_277),
.B(n_243),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_262),
.B(n_160),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

BUFx6f_ASAP7_75t_SL g331 ( 
.A(n_254),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_246),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_263),
.B(n_245),
.C(n_212),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_297),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_248),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_246),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_290),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_290),
.B(n_246),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g339 ( 
.A(n_293),
.B(n_218),
.C(n_246),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_291),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_241),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_271),
.A2(n_242),
.B1(n_161),
.B2(n_196),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_279),
.B(n_202),
.C(n_166),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_R g348 ( 
.A(n_255),
.B(n_163),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_291),
.B(n_167),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_250),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_258),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_289),
.B(n_241),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_289),
.B(n_241),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_283),
.B(n_170),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_283),
.B(n_171),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_289),
.B(n_172),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_289),
.B(n_182),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_254),
.B(n_186),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_355),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_351),
.B(n_188),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_357),
.B(n_190),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_194),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_299),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_197),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_198),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_307),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_314),
.B(n_200),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_334),
.B(n_249),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_308),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_205),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_337),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_335),
.A2(n_240),
.B1(n_249),
.B2(n_206),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_329),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_316),
.B(n_216),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_343),
.B(n_216),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_332),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_336),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_350),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_348),
.Y(n_385)
);

OR2x6_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_224),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_333),
.A2(n_244),
.B1(n_224),
.B2(n_13),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_300),
.B(n_244),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_23),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

A2O1A1Ixp33_ASAP7_75t_L g392 ( 
.A1(n_315),
.A2(n_317),
.B(n_310),
.C(n_312),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_302),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_303),
.Y(n_395)
);

INVx3_ASAP7_75t_SL g396 ( 
.A(n_341),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_323),
.B(n_11),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_353),
.B(n_12),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_331),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_325),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_356),
.Y(n_405)
);

BUFx4f_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_361),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_304),
.B(n_24),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_320),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_325),
.B(n_25),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_325),
.B(n_26),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

OR2x6_ASAP7_75t_L g416 ( 
.A(n_345),
.B(n_29),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_320),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g419 ( 
.A1(n_306),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_344),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_338),
.Y(n_422)
);

INVx3_ASAP7_75t_SL g423 ( 
.A(n_322),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_320),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_305),
.Y(n_425)
);

OR2x6_ASAP7_75t_L g426 ( 
.A(n_347),
.B(n_152),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_318),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_320),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_301),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_395),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_383),
.A2(n_380),
.B(n_379),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_406),
.B(n_362),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_366),
.A2(n_344),
.B(n_349),
.C(n_321),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_405),
.B(n_43),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_45),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_48),
.Y(n_438)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_371),
.B(n_49),
.Y(n_439)
);

BUFx12f_ASAP7_75t_L g440 ( 
.A(n_409),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_404),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_151),
.B(n_53),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_389),
.A2(n_51),
.B(n_54),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_55),
.Y(n_444)
);

O2A1O1Ixp5_ASAP7_75t_L g445 ( 
.A1(n_365),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_368),
.B(n_60),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_61),
.C(n_62),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_397),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_381),
.A2(n_63),
.B(n_64),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_387),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_70),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_423),
.B(n_378),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_375),
.B(n_72),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_369),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_R g457 ( 
.A(n_385),
.B(n_77),
.Y(n_457)
);

OR2x6_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_78),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_382),
.B(n_81),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_406),
.B(n_363),
.Y(n_460)
);

AOI21x1_ASAP7_75t_L g461 ( 
.A1(n_390),
.A2(n_83),
.B(n_86),
.Y(n_461)
);

O2A1O1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_401),
.A2(n_373),
.B(n_399),
.C(n_392),
.Y(n_462)
);

AO32x2_ASAP7_75t_L g463 ( 
.A1(n_420),
.A2(n_87),
.A3(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_92),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_427),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_367),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_413),
.B(n_93),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_363),
.B(n_96),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_100),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_377),
.A2(n_421),
.B1(n_387),
.B2(n_403),
.Y(n_470)
);

O2A1O1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_411),
.A2(n_101),
.B(n_103),
.C(n_104),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_372),
.B(n_106),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_L g473 ( 
.A1(n_376),
.A2(n_107),
.B(n_108),
.C(n_109),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_386),
.B(n_110),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_111),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_398),
.A2(n_112),
.B(n_113),
.C(n_114),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_386),
.B(n_118),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_427),
.B(n_120),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_388),
.Y(n_480)
);

A2O1A1Ixp33_ASAP7_75t_L g481 ( 
.A1(n_391),
.A2(n_121),
.B(n_122),
.C(n_123),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g482 ( 
.A(n_393),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_417),
.A2(n_124),
.B(n_125),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_386),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_415),
.Y(n_485)
);

BUFx12f_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_414),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_466),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_433),
.A2(n_442),
.B(n_459),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_462),
.A2(n_418),
.B(n_424),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_465),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_432),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_465),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_439),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_431),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_458),
.B(n_416),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_484),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_364),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_461),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_430),
.Y(n_503)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_476),
.A2(n_419),
.B(n_428),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_458),
.B(n_416),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_448),
.Y(n_508)
);

CKINVDCx11_ASAP7_75t_R g509 ( 
.A(n_458),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_464),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_468),
.B(n_426),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_450),
.B(n_426),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_475),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_479),
.A2(n_459),
.B(n_445),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_482),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_435),
.A2(n_429),
.B(n_415),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_437),
.A2(n_449),
.B(n_483),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_441),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_446),
.A2(n_415),
.B(n_388),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_463),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_457),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_434),
.Y(n_525)
);

BUFx12f_ASAP7_75t_L g526 ( 
.A(n_434),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

NAND2x1p5_ASAP7_75t_L g528 ( 
.A(n_460),
.B(n_472),
.Y(n_528)
);

NAND2x1p5_ASAP7_75t_L g529 ( 
.A(n_436),
.B(n_388),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_438),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_454),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_469),
.A2(n_426),
.B(n_128),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_467),
.B(n_408),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_511),
.B(n_525),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_526),
.A2(n_447),
.B1(n_451),
.B2(n_452),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_493),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_514),
.A2(n_455),
.B(n_473),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_526),
.A2(n_396),
.B1(n_451),
.B2(n_402),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_SL g542 ( 
.A1(n_533),
.A2(n_408),
.B1(n_480),
.B2(n_443),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_495),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_497),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_511),
.B(n_481),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_471),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_488),
.Y(n_547)
);

INVx6_ASAP7_75t_L g548 ( 
.A(n_501),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_491),
.A2(n_477),
.B(n_129),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_500),
.A2(n_126),
.B1(n_132),
.B2(n_133),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_501),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_533),
.B(n_497),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_507),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_507),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_489),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_531),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_521),
.A2(n_138),
.B(n_139),
.Y(n_558)
);

BUFx4_ASAP7_75t_R g559 ( 
.A(n_520),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_499),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_499),
.Y(n_562)
);

BUFx2_ASAP7_75t_SL g563 ( 
.A(n_520),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_512),
.B(n_140),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_515),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_510),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_513),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_503),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_514),
.A2(n_147),
.B(n_148),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_512),
.B(n_517),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_503),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_516),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_498),
.A2(n_506),
.B1(n_496),
.B2(n_534),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_516),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_524),
.B(n_534),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_531),
.A2(n_506),
.B1(n_498),
.B2(n_534),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_498),
.A2(n_506),
.B1(n_487),
.B2(n_509),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_538),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_536),
.B(n_505),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_537),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_537),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_535),
.B(n_506),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_577),
.B(n_505),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_535),
.B(n_498),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_494),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_540),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_570),
.B(n_519),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_564),
.B(n_495),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_R g590 ( 
.A(n_565),
.B(n_515),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_561),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_565),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_540),
.B(n_505),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_545),
.A2(n_509),
.B1(n_487),
.B2(n_528),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_567),
.B(n_505),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_575),
.B(n_523),
.Y(n_596)
);

AO31x2_ASAP7_75t_L g597 ( 
.A1(n_572),
.A2(n_574),
.A3(n_527),
.B(n_556),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_547),
.B(n_516),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_567),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_543),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_541),
.A2(n_528),
.B(n_529),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_564),
.B(n_492),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_552),
.B(n_492),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_559),
.B(n_505),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_562),
.B(n_492),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_562),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_543),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_544),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_555),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_SL g610 ( 
.A(n_566),
.B(n_546),
.C(n_555),
.Y(n_610)
);

NOR3xp33_ASAP7_75t_SL g611 ( 
.A(n_556),
.B(n_487),
.C(n_532),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_545),
.B(n_522),
.Y(n_612)
);

NAND2x1p5_ASAP7_75t_L g613 ( 
.A(n_551),
.B(n_492),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_560),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_560),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_SL g616 ( 
.A(n_576),
.B(n_487),
.C(n_532),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_563),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_544),
.B(n_522),
.Y(n_618)
);

NAND3xp33_ASAP7_75t_SL g619 ( 
.A(n_542),
.B(n_528),
.C(n_529),
.Y(n_619)
);

CKINVDCx16_ASAP7_75t_R g620 ( 
.A(n_573),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_553),
.B(n_492),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_549),
.A2(n_502),
.B(n_518),
.Y(n_622)
);

NOR3xp33_ASAP7_75t_SL g623 ( 
.A(n_573),
.B(n_487),
.C(n_486),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_553),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_549),
.A2(n_504),
.B(n_518),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_554),
.Y(n_626)
);

CKINVDCx12_ASAP7_75t_R g627 ( 
.A(n_563),
.Y(n_627)
);

NAND2xp33_ASAP7_75t_R g628 ( 
.A(n_569),
.B(n_502),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_612),
.B(n_522),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_619),
.A2(n_557),
.B1(n_487),
.B2(n_550),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_597),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_612),
.B(n_522),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_602),
.Y(n_633)
);

INVx4_ASAP7_75t_R g634 ( 
.A(n_617),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_574),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_597),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_623),
.B(n_572),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_583),
.B(n_593),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_596),
.B(n_522),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_591),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_598),
.B(n_558),
.Y(n_641)
);

OR2x2_ASAP7_75t_L g642 ( 
.A(n_620),
.B(n_579),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_486),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_580),
.B(n_571),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_579),
.B(n_558),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_595),
.B(n_558),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_585),
.B(n_571),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_581),
.B(n_599),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_606),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_603),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_586),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_618),
.B(n_588),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_609),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_614),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_615),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_618),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_589),
.B(n_529),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_619),
.A2(n_504),
.B1(n_539),
.B2(n_571),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_608),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_584),
.B(n_569),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_578),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_616),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_605),
.B(n_569),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_600),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_629),
.B(n_616),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_640),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_652),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_653),
.B(n_601),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_665),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_643),
.B(n_592),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_651),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_629),
.B(n_611),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_632),
.B(n_638),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_641),
.B(n_625),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_652),
.Y(n_676)
);

INVxp67_ASAP7_75t_SL g677 ( 
.A(n_650),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_632),
.B(n_611),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_630),
.A2(n_604),
.B1(n_594),
.B2(n_610),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_665),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_641),
.B(n_625),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_638),
.B(n_622),
.Y(n_682)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_662),
.B(n_587),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_654),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_661),
.B(n_626),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_654),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_661),
.B(n_621),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_645),
.B(n_569),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_642),
.B(n_624),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

INVxp67_ASAP7_75t_SL g691 ( 
.A(n_657),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_655),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_631),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_649),
.B(n_578),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_636),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_655),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_673),
.B(n_678),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_677),
.B(n_647),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_668),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_674),
.B(n_647),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_668),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_676),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_670),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_694),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_676),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_682),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_692),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_694),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_692),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_673),
.B(n_664),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_678),
.B(n_664),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_674),
.B(n_642),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_684),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_712),
.B(n_681),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_701),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_699),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_697),
.A2(n_679),
.B1(n_663),
.B2(n_610),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_697),
.B(n_671),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_699),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_701),
.Y(n_720)
);

O2A1O1Ixp5_ASAP7_75t_R g721 ( 
.A1(n_698),
.A2(n_669),
.B(n_689),
.C(n_672),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_710),
.B(n_687),
.Y(n_722)
);

OAI33xp33_ASAP7_75t_L g723 ( 
.A1(n_713),
.A2(n_675),
.A3(n_681),
.B1(n_686),
.B2(n_696),
.B3(n_690),
.Y(n_723)
);

OAI22xp5_ASAP7_75t_L g724 ( 
.A1(n_717),
.A2(n_663),
.B1(n_708),
.B2(n_704),
.Y(n_724)
);

NOR3xp33_ASAP7_75t_L g725 ( 
.A(n_721),
.B(n_667),
.C(n_658),
.Y(n_725)
);

AOI211xp5_ASAP7_75t_L g726 ( 
.A1(n_717),
.A2(n_682),
.B(n_710),
.C(n_711),
.Y(n_726)
);

AOI21xp33_ASAP7_75t_SL g727 ( 
.A1(n_718),
.A2(n_590),
.B(n_703),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_723),
.A2(n_683),
.B(n_691),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_724),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_725),
.B(n_711),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_L g731 ( 
.A1(n_728),
.A2(n_700),
.B(n_714),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_727),
.Y(n_732)
);

NOR2x1_ASAP7_75t_L g733 ( 
.A(n_729),
.B(n_715),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_730),
.Y(n_734)
);

AOI21xp33_ASAP7_75t_L g735 ( 
.A1(n_732),
.A2(n_726),
.B(n_675),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_731),
.B(n_704),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_736),
.A2(n_720),
.B(n_703),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_734),
.A2(n_666),
.B1(n_694),
.B2(n_708),
.Y(n_738)
);

AOI211xp5_ASAP7_75t_L g739 ( 
.A1(n_737),
.A2(n_735),
.B(n_733),
.C(n_680),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_738),
.B(n_706),
.Y(n_740)
);

OAI221xp5_ASAP7_75t_SL g741 ( 
.A1(n_738),
.A2(n_722),
.B1(n_706),
.B2(n_645),
.C(n_659),
.Y(n_741)
);

NOR2x1_ASAP7_75t_L g742 ( 
.A(n_740),
.B(n_607),
.Y(n_742)
);

AND3x4_ASAP7_75t_L g743 ( 
.A(n_739),
.B(n_634),
.C(n_670),
.Y(n_743)
);

NOR2x1_ASAP7_75t_L g744 ( 
.A(n_741),
.B(n_600),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_708),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_740),
.A2(n_666),
.B1(n_633),
.B2(n_637),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_740),
.Y(n_747)
);

OAI321xp33_ASAP7_75t_L g748 ( 
.A1(n_747),
.A2(n_600),
.A3(n_648),
.B1(n_634),
.B2(n_639),
.C(n_688),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_L g749 ( 
.A1(n_746),
.A2(n_719),
.B1(n_716),
.B2(n_709),
.C(n_707),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_742),
.B(n_704),
.Y(n_750)
);

NOR3xp33_ASAP7_75t_SL g751 ( 
.A(n_743),
.B(n_627),
.C(n_702),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_745),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_744),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_745),
.Y(n_754)
);

NOR4xp25_ASAP7_75t_SL g755 ( 
.A(n_753),
.B(n_628),
.C(n_702),
.D(n_660),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_754),
.Y(n_756)
);

AND3x2_ASAP7_75t_L g757 ( 
.A(n_752),
.B(n_750),
.C(n_751),
.Y(n_757)
);

OAI211xp5_ASAP7_75t_L g758 ( 
.A1(n_749),
.A2(n_587),
.B(n_662),
.C(n_551),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_748),
.Y(n_759)
);

AOI222xp33_ASAP7_75t_L g760 ( 
.A1(n_753),
.A2(n_705),
.B1(n_644),
.B2(n_637),
.C1(n_635),
.C2(n_660),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_756),
.Y(n_761)
);

AOI22x1_ASAP7_75t_L g762 ( 
.A1(n_759),
.A2(n_551),
.B1(n_613),
.B2(n_705),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_633),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_758),
.A2(n_637),
.B1(n_635),
.B2(n_685),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_760),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_755),
.A2(n_635),
.B1(n_685),
.B2(n_644),
.Y(n_766)
);

NAND4xp75_ASAP7_75t_L g767 ( 
.A(n_756),
.B(n_649),
.C(n_539),
.D(n_490),
.Y(n_767)
);

OA22x2_ASAP7_75t_L g768 ( 
.A1(n_757),
.A2(n_644),
.B1(n_693),
.B2(n_690),
.Y(n_768)
);

AO22x2_ASAP7_75t_L g769 ( 
.A1(n_761),
.A2(n_656),
.B1(n_693),
.B2(n_695),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_765),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_763),
.B(n_687),
.Y(n_771)
);

OAI31xp33_ASAP7_75t_L g772 ( 
.A1(n_762),
.A2(n_613),
.A3(n_688),
.B(n_646),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_768),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_766),
.B(n_633),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_773),
.Y(n_775)
);

AOI22x1_ASAP7_75t_L g776 ( 
.A1(n_770),
.A2(n_769),
.B1(n_772),
.B2(n_774),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_771),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_770),
.A2(n_764),
.B(n_767),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_SL g779 ( 
.A1(n_775),
.A2(n_538),
.B1(n_548),
.B2(n_662),
.Y(n_779)
);

AOI221xp5_ASAP7_75t_L g780 ( 
.A1(n_777),
.A2(n_656),
.B1(n_633),
.B2(n_502),
.C(n_568),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_777),
.A2(n_538),
.B1(n_548),
.B2(n_662),
.Y(n_781)
);

NOR2x1_ASAP7_75t_L g782 ( 
.A(n_779),
.B(n_776),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_781),
.B(n_778),
.C(n_662),
.Y(n_783)
);

OAI31xp33_ASAP7_75t_L g784 ( 
.A1(n_783),
.A2(n_780),
.A3(n_568),
.B(n_554),
.Y(n_784)
);

XNOR2xp5_ASAP7_75t_L g785 ( 
.A(n_784),
.B(n_782),
.Y(n_785)
);

AOI31xp33_ASAP7_75t_L g786 ( 
.A1(n_785),
.A2(n_646),
.A3(n_548),
.B(n_662),
.Y(n_786)
);


endmodule