module fake_jpeg_14607_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

AND2x2_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_3),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_6),
.Y(n_13)
);

OR2x2_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_15),
.Y(n_18)
);

CKINVDCx12_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_0),
.B(n_1),
.Y(n_15)
);

NOR2x1_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_1),
.Y(n_17)
);

AND2x6_ASAP7_75t_L g20 ( 
.A(n_17),
.B(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_1),
.Y(n_26)
);

AO22x1_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_16),
.B1(n_13),
.B2(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_26),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_16),
.B(n_8),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_6),
.C(n_8),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_12),
.Y(n_32)
);

XOR2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_12),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_25),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI322xp5_ASAP7_75t_L g38 ( 
.A1(n_36),
.A2(n_2),
.A3(n_4),
.B1(n_10),
.B2(n_23),
.C1(n_30),
.C2(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_36),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);


endmodule