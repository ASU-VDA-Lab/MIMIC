module real_jpeg_1599_n_16 (n_5, n_4, n_8, n_0, n_12, n_309, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_309;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_176;
wire n_286;
wire n_300;
wire n_215;
wire n_221;
wire n_249;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_299;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_213;
wire n_128;
wire n_179;
wire n_216;
wire n_133;
wire n_202;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_43),
.B1(n_64),
.B2(n_65),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_1),
.A2(n_35),
.B1(n_37),
.B2(n_43),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_43),
.B1(n_49),
.B2(n_52),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_2),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_3),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_137),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_3),
.A2(n_49),
.B1(n_52),
.B2(n_137),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_137),
.Y(n_231)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_5),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_5),
.A2(n_49),
.B1(n_52),
.B2(n_161),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_161),
.Y(n_234)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_7),
.A2(n_49),
.B1(n_52),
.B2(n_57),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_7),
.A2(n_57),
.B1(n_64),
.B2(n_65),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_112)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_10),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_10),
.A2(n_39),
.B1(n_64),
.B2(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_10),
.A2(n_39),
.B1(n_49),
.B2(n_52),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_11),
.A2(n_35),
.B1(n_37),
.B2(n_67),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_11),
.A2(n_49),
.B1(n_52),
.B2(n_67),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_13),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_13),
.B(n_49),
.C(n_51),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_13),
.A2(n_35),
.B1(n_37),
.B2(n_152),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_13),
.B(n_88),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_13),
.B(n_47),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_13),
.B(n_30),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_13),
.A2(n_30),
.B(n_225),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_13),
.B(n_100),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_13),
.A2(n_64),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_14),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_135),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_14),
.A2(n_49),
.B1(n_52),
.B2(n_135),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_135),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_115),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_20),
.B(n_101),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_83),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g303 ( 
.A(n_21),
.B(n_74),
.CI(n_83),
.CON(n_303),
.SN(n_303)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_59),
.B2(n_73),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_45),
.B1(n_46),
.B2(n_58),
.Y(n_23)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_46),
.C(n_59),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_38),
.B(n_40),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_25),
.A2(n_38),
.B1(n_44),
.B2(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_25),
.B(n_42),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_25),
.A2(n_44),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_26),
.A2(n_41),
.B(n_112),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_26),
.A2(n_110),
.B(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_26),
.A2(n_34),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_26),
.A2(n_34),
.B1(n_158),
.B2(n_246),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_27)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OA22x2_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_28),
.A2(n_30),
.A3(n_35),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_30),
.A2(n_31),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_30),
.B(n_61),
.C(n_65),
.Y(n_153)
);

CKINVDCx6p67_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_31),
.A2(n_62),
.B(n_151),
.C(n_153),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_33),
.B(n_37),
.Y(n_226)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_34),
.A2(n_77),
.B(n_113),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_34),
.B(n_152),
.Y(n_188)
);

CKINVDCx6p67_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_35),
.B(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_44),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_45),
.A2(n_46),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_53),
.B(n_55),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_47),
.B(n_82),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_47),
.A2(n_53),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_47),
.A2(n_53),
.B1(n_190),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_56),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_48),
.A2(n_81),
.B(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_48),
.A2(n_92),
.B1(n_93),
.B2(n_130),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_48),
.A2(n_92),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_49),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_49),
.B(n_203),
.Y(n_202)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_53),
.A2(n_79),
.B(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_56),
.A2(n_92),
.B(n_94),
.Y(n_264)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_73),
.B1(n_104),
.B2(n_114),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_68),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_60),
.A2(n_63),
.B1(n_70),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_60),
.A2(n_70),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_60),
.A2(n_70),
.B1(n_134),
.B2(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_60),
.A2(n_70),
.B1(n_160),
.B2(n_260),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_65),
.B(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_97),
.B(n_99),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_70),
.A2(n_136),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B(n_95),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_84),
.A2(n_91),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_84),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_84),
.A2(n_95),
.B1(n_96),
.B2(n_167),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_85),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_85),
.A2(n_87),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_85),
.A2(n_89),
.B(n_127),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_86),
.B(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_88),
.B1(n_126),
.B2(n_155),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_86),
.A2(n_142),
.B(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_86),
.A2(n_88),
.B1(n_152),
.B2(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_86),
.A2(n_88),
.B1(n_205),
.B2(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_89),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_87),
.A2(n_144),
.B(n_156),
.Y(n_251)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_90),
.B(n_296),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_91),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B(n_94),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_100),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_300),
.B(n_304),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_289),
.B(n_299),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_178),
.B(n_288),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_162),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_120),
.B(n_162),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_139),
.C(n_147),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_121),
.B(n_139),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_131),
.B2(n_132),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_122),
.B(n_133),
.C(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_129),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_124),
.B(n_129),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_138),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_147),
.B(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_157),
.C(n_159),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_148),
.B(n_157),
.CI(n_159),
.CON(n_276),
.SN(n_276)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_151),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_154),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_177),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_166),
.B(n_169),
.C(n_177),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_175),
.Y(n_176)
);

AOI321xp33_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_271),
.A3(n_280),
.B1(n_286),
.B2(n_287),
.C(n_309),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_254),
.B(n_270),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_236),
.B(n_253),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_218),
.B(n_235),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_199),
.B(n_217),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_192),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_192),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_189),
.C(n_220),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_211),
.B(n_216),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_206),
.B(n_210),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_209),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_215),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_221),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_229),
.C(n_232),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_227),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_227),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_252),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_252),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_249),
.C(n_250),
.Y(n_267)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_256),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_265),
.B2(n_266),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_267),
.C(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_276),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g307 ( 
.A(n_276),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_277),
.A2(n_278),
.B1(n_279),
.B2(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_298),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_293),
.B2(n_294),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_295),
.C(n_297),
.Y(n_302)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_302),
.B(n_303),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g308 ( 
.A(n_303),
.Y(n_308)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);


endmodule