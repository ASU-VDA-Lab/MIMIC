module fake_jpeg_27535_n_76 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_16;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx16_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_3),
.Y(n_9)
);

INVx11_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_14),
.Y(n_24)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_1),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_11),
.B(n_14),
.C(n_13),
.Y(n_23)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_24),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_26),
.A2(n_18),
.B1(n_12),
.B2(n_14),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_29),
.A2(n_13),
.B1(n_21),
.B2(n_18),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_17),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_SL g44 ( 
.A(n_30),
.B(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_46),
.B(n_36),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_16),
.B(n_12),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_15),
.B1(n_9),
.B2(n_12),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_36),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_1),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_49),
.B(n_8),
.Y(n_62)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_53),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_56),
.Y(n_59)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_35),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_46),
.B1(n_44),
.B2(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_57),
.C(n_52),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_59),
.C(n_60),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g64 ( 
.A1(n_58),
.A2(n_56),
.A3(n_57),
.B1(n_51),
.B2(n_55),
.C(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_38),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_7),
.B(n_4),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_22),
.C(n_4),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_5),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_20),
.C(n_22),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_20),
.B1(n_37),
.B2(n_2),
.Y(n_76)
);


endmodule