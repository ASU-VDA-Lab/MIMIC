module fake_jpeg_26184_n_276 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_276);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_276;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_41),
.Y(n_45)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_19),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_53),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_19),
.B(n_32),
.C(n_18),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_24),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_60),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_36),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_22),
.B1(n_29),
.B2(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_59),
.B1(n_42),
.B2(n_39),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_22),
.B1(n_29),
.B2(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_31),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_21),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_36),
.B(n_35),
.C(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_64),
.A2(n_88),
.B(n_89),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_71),
.B1(n_79),
.B2(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_33),
.B1(n_34),
.B2(n_28),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_46),
.B1(n_47),
.B2(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_33),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_17),
.B(n_32),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_39),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_17),
.B(n_32),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_78),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_44),
.A2(n_41),
.B1(n_23),
.B2(n_18),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_44),
.A2(n_23),
.B1(n_17),
.B2(n_18),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_95),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_42),
.B1(n_61),
.B2(n_58),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_30),
.Y(n_87)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_53),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_54),
.B(n_23),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_94),
.Y(n_116)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_50),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_54),
.C(n_60),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_114),
.C(n_89),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_106),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_56),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_56),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_61),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_61),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_117),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_46),
.B1(n_37),
.B2(n_27),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_120),
.B(n_51),
.Y(n_123)
);

OA22x2_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_46),
.B1(n_35),
.B2(n_43),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_82),
.A2(n_27),
.B1(n_24),
.B2(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_51),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_117),
.B1(n_110),
.B2(n_92),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_125),
.B(n_128),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_118),
.A2(n_88),
.B(n_63),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_127),
.B(n_135),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_133),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_144),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_121),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_66),
.B(n_63),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_134),
.B(n_130),
.Y(n_175)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_76),
.B(n_90),
.C(n_72),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_111),
.A2(n_76),
.B(n_90),
.Y(n_135)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_141),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_138),
.B(n_142),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_11),
.B(n_16),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_6),
.B(n_14),
.Y(n_155)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_30),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_97),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_96),
.B(n_110),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_85),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_150),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_119),
.B1(n_111),
.B2(n_103),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_119),
.B1(n_103),
.B2(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_81),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_155),
.B(n_171),
.C(n_35),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_157),
.A2(n_172),
.B(n_178),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_159),
.A2(n_123),
.B1(n_136),
.B2(n_143),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_166),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_109),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_121),
.B1(n_108),
.B2(n_114),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_136),
.B1(n_43),
.B2(n_35),
.Y(n_202)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_168),
.B(n_170),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_107),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_135),
.A2(n_95),
.A3(n_38),
.B1(n_40),
.B2(n_43),
.C1(n_31),
.C2(n_35),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_124),
.A2(n_107),
.B(n_98),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_98),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_96),
.Y(n_174)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_133),
.A2(n_24),
.B1(n_26),
.B2(n_31),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_81),
.C(n_65),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_134),
.C(n_141),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_197),
.Y(n_214)
);

AOI22x1_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_124),
.B1(n_149),
.B2(n_147),
.Y(n_187)
);

OAI22x1_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_183),
.B1(n_189),
.B2(n_165),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_190),
.C(n_198),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_147),
.B1(n_127),
.B2(n_129),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_191),
.B1(n_169),
.B2(n_159),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_140),
.C(n_143),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_137),
.B1(n_147),
.B2(n_128),
.Y(n_191)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVxp33_ASAP7_75t_SL g193 ( 
.A(n_180),
.Y(n_193)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_202),
.B1(n_187),
.B2(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_132),
.C(n_134),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_126),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_29),
.C(n_22),
.Y(n_216)
);

OAI322xp33_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_156),
.A3(n_164),
.B1(n_162),
.B2(n_175),
.C1(n_154),
.C2(n_158),
.Y(n_204)
);

OAI322xp33_ASAP7_75t_L g228 ( 
.A1(n_204),
.A2(n_219),
.A3(n_194),
.B1(n_10),
.B2(n_14),
.C1(n_11),
.C2(n_4),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_205),
.A2(n_210),
.B1(n_212),
.B2(n_38),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_202),
.B1(n_201),
.B2(n_94),
.Y(n_231)
);

XNOR2x2_ASAP7_75t_SL g207 ( 
.A(n_188),
.B(n_156),
.Y(n_207)
);

AOI321xp33_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_213),
.A3(n_8),
.B1(n_14),
.B2(n_10),
.C(n_6),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_183),
.A2(n_153),
.B(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_209),
.B(n_211),
.Y(n_234)
);

OAI321xp33_ASAP7_75t_L g211 ( 
.A1(n_199),
.A2(n_158),
.A3(n_153),
.B1(n_180),
.B2(n_166),
.C(n_167),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_176),
.B1(n_179),
.B2(n_178),
.Y(n_212)
);

AOI321xp33_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_176),
.A3(n_21),
.B1(n_12),
.B2(n_10),
.C(n_4),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_222),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_220),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_198),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

OAI322xp33_ASAP7_75t_L g219 ( 
.A1(n_182),
.A2(n_21),
.A3(n_25),
.B1(n_29),
.B2(n_11),
.C1(n_4),
.C2(n_6),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_25),
.B1(n_95),
.B2(n_65),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_38),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_195),
.C(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_224),
.C(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_195),
.C(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_192),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_229),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_231),
.B1(n_208),
.B2(n_216),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_230),
.A2(n_237),
.B(n_205),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_7),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_94),
.C(n_43),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_239),
.B(n_242),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_209),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_246),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_235),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_245),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_208),
.B1(n_214),
.B2(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_213),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_9),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.C(n_247),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_9),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_248),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_258),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_227),
.B(n_230),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_253),
.A2(n_259),
.B(n_249),
.Y(n_261)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_0),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_223),
.C(n_233),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_242),
.A2(n_231),
.B(n_232),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_261),
.B(n_263),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_238),
.B(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_262),
.B(n_266),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_8),
.C(n_9),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_8),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_260),
.A2(n_256),
.B(n_252),
.C(n_257),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_0),
.C(n_2),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_3),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_271),
.C(n_270),
.Y(n_275)
);

HAxp5_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_269),
.CON(n_276),
.SN(n_276)
);


endmodule