module fake_jpeg_2397_n_224 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_224);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_14),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_6),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_67),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx9p33_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_86),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_65),
.Y(n_87)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_70),
.C(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_61),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_73),
.B(n_69),
.C(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_89),
.B(n_63),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_97),
.B1(n_63),
.B2(n_62),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_53),
.B1(n_77),
.B2(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_53),
.B1(n_57),
.B2(n_77),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_61),
.B1(n_62),
.B2(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_64),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_99),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_75),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_82),
.B1(n_83),
.B2(n_94),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_94),
.B1(n_95),
.B2(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_113),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_108),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_68),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_58),
.Y(n_125)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_94),
.B1(n_82),
.B2(n_76),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_119),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_80),
.B(n_72),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_55),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_121),
.A2(n_128),
.B1(n_4),
.B2(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_82),
.B1(n_89),
.B2(n_70),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_66),
.C(n_60),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_132),
.C(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_112),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_78),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_23),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_140),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_102),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_141),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_20),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_0),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_143),
.C(n_146),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_120),
.A2(n_106),
.B1(n_80),
.B2(n_25),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_50),
.C(n_47),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_130),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_157),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_2),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_152),
.A2(n_163),
.B1(n_14),
.B2(n_15),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_26),
.C(n_43),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_129),
.C(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_9),
.B(n_10),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_134),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_125),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_12),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_169),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_143),
.B(n_158),
.Y(n_169)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_122),
.C(n_30),
.D(n_31),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_SL g198 ( 
.A1(n_171),
.A2(n_176),
.A3(n_38),
.B1(n_42),
.B2(n_27),
.C1(n_36),
.C2(n_45),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_11),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_175),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_28),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_180),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_13),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_163),
.B1(n_155),
.B2(n_144),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_177),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_156),
.B(n_32),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_15),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_196),
.B1(n_166),
.B2(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_146),
.C(n_37),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_16),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_197),
.B(n_198),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_177),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_205),
.B1(n_206),
.B2(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_186),
.B1(n_185),
.B2(n_173),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_204),
.A2(n_18),
.B1(n_19),
.B2(n_39),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_186),
.B1(n_180),
.B2(n_173),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_189),
.C(n_193),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_210),
.C(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_207),
.B(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_194),
.C(n_183),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_212),
.B(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_213),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_216),
.B(n_209),
.C(n_207),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g220 ( 
.A1(n_218),
.A2(n_219),
.B(n_217),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_199),
.C(n_200),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_216),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_215),
.B(n_201),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_223),
.B(n_41),
.Y(n_224)
);


endmodule