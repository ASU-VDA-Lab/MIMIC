module real_aes_6779_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_1), .A2(n_161), .B(n_164), .C(n_244), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_2), .A2(n_190), .B(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g491 ( .A(n_3), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_4), .B(n_220), .Y(n_219) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_5), .A2(n_190), .B(n_475), .Y(n_474) );
AND2x6_ASAP7_75t_L g161 ( .A(n_6), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g257 ( .A(n_7), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_8), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_8), .B(n_41), .Y(n_126) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_9), .A2(n_189), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_10), .B(n_173), .Y(n_246) );
INVx1_ASAP7_75t_L g479 ( .A(n_11), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_12), .B(n_214), .Y(n_514) );
INVx1_ASAP7_75t_L g153 ( .A(n_13), .Y(n_153) );
INVx1_ASAP7_75t_L g526 ( .A(n_14), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_15), .A2(n_78), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_15), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_16), .A2(n_198), .B(n_279), .C(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_17), .B(n_220), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_18), .B(n_457), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_19), .B(n_190), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_20), .B(n_204), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_21), .A2(n_214), .B(n_265), .C(n_267), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_22), .B(n_220), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_23), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_24), .A2(n_200), .B(n_281), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_25), .B(n_173), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g155 ( .A(n_26), .Y(n_155) );
INVx1_ASAP7_75t_L g227 ( .A(n_27), .Y(n_227) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_28), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_29), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_30), .B(n_173), .Y(n_492) );
INVx1_ASAP7_75t_L g196 ( .A(n_31), .Y(n_196) );
INVx1_ASAP7_75t_L g469 ( .A(n_32), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_33), .A2(n_131), .B1(n_132), .B2(n_133), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_33), .Y(n_131) );
INVx2_ASAP7_75t_L g159 ( .A(n_34), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_35), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_36), .A2(n_214), .B(n_215), .C(n_217), .Y(n_213) );
INVxp67_ASAP7_75t_L g199 ( .A(n_37), .Y(n_199) );
CKINVDCx14_ASAP7_75t_R g212 ( .A(n_38), .Y(n_212) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_39), .A2(n_164), .B(n_226), .C(n_230), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_40), .A2(n_161), .B(n_164), .C(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g113 ( .A(n_41), .Y(n_113) );
INVx1_ASAP7_75t_L g468 ( .A(n_42), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_43), .A2(n_175), .B(n_255), .C(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_44), .B(n_173), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_45), .Y(n_232) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_46), .Y(n_192) );
INVx1_ASAP7_75t_L g263 ( .A(n_47), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_48), .Y(n_470) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_49), .A2(n_58), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_49), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_50), .B(n_190), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_51), .A2(n_164), .B1(n_267), .B2(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_52), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_53), .Y(n_488) );
CKINVDCx14_ASAP7_75t_R g253 ( .A(n_54), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_55), .A2(n_217), .B(n_255), .C(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_56), .Y(n_538) );
INVx1_ASAP7_75t_L g476 ( .A(n_57), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_58), .Y(n_740) );
INVx1_ASAP7_75t_L g162 ( .A(n_59), .Y(n_162) );
INVx1_ASAP7_75t_L g152 ( .A(n_60), .Y(n_152) );
INVx1_ASAP7_75t_SL g216 ( .A(n_61), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_62), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_63), .A2(n_738), .B1(n_741), .B2(n_742), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_63), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_64), .B(n_220), .Y(n_269) );
INVx1_ASAP7_75t_L g168 ( .A(n_65), .Y(n_168) );
AOI222xp33_ASAP7_75t_SL g128 ( .A1(n_66), .A2(n_129), .B1(n_130), .B2(n_136), .C1(n_729), .C2(n_731), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_SL g456 ( .A1(n_67), .A2(n_217), .B(n_457), .C(n_458), .Y(n_456) );
INVxp67_ASAP7_75t_L g459 ( .A(n_68), .Y(n_459) );
INVx1_ASAP7_75t_L g111 ( .A(n_69), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_70), .A2(n_190), .B(n_252), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_71), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_72), .A2(n_190), .B(n_276), .Y(n_275) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_73), .Y(n_472) );
INVx1_ASAP7_75t_L g532 ( .A(n_74), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_75), .A2(n_189), .B(n_191), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_76), .Y(n_224) );
INVx1_ASAP7_75t_L g277 ( .A(n_77), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_78), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_79), .A2(n_161), .B(n_164), .C(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_80), .A2(n_190), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g280 ( .A(n_81), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_82), .B(n_197), .Y(n_503) );
INVx2_ASAP7_75t_L g150 ( .A(n_83), .Y(n_150) );
INVx1_ASAP7_75t_L g245 ( .A(n_84), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_85), .B(n_457), .Y(n_504) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_86), .A2(n_161), .B(n_164), .C(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g108 ( .A(n_87), .Y(n_108) );
OR2x2_ASAP7_75t_L g123 ( .A(n_87), .B(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g443 ( .A(n_87), .B(n_125), .Y(n_443) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_88), .A2(n_164), .B(n_167), .C(n_177), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_89), .B(n_182), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_90), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_91), .A2(n_161), .B(n_164), .C(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_92), .Y(n_518) );
INVx1_ASAP7_75t_L g455 ( .A(n_93), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_94), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_95), .B(n_197), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_96), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_97), .B(n_148), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_98), .B(n_148), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g266 ( .A(n_100), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_101), .A2(n_190), .B(n_454), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_102), .A2(n_104), .B1(n_114), .B2(n_744), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g745 ( .A(n_105), .Y(n_745) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .C(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g125 ( .A(n_107), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g728 ( .A(n_108), .B(n_125), .Y(n_728) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_108), .B(n_124), .Y(n_733) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_128), .B1(n_734), .B2(n_735), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_SL g734 ( .A(n_119), .Y(n_734) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_121), .A2(n_736), .B(n_743), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_127), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_123), .Y(n_743) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_443), .B1(n_444), .B2(n_726), .Y(n_136) );
INVx2_ASAP7_75t_L g730 ( .A(n_137), .Y(n_730) );
XOR2xp5_ASAP7_75t_L g736 ( .A(n_137), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_377), .Y(n_137) );
NAND5xp2_ASAP7_75t_L g138 ( .A(n_139), .B(n_306), .C(n_336), .D(n_357), .E(n_363), .Y(n_138) );
AOI221xp5_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_236), .B1(n_270), .B2(n_272), .C(n_283), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_233), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_205), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_SL g357 ( .A1(n_144), .A2(n_221), .B(n_358), .C(n_361), .Y(n_357) );
AND2x2_ASAP7_75t_L g427 ( .A(n_144), .B(n_222), .Y(n_427) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_183), .Y(n_144) );
AND2x2_ASAP7_75t_L g285 ( .A(n_145), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g289 ( .A(n_145), .B(n_286), .Y(n_289) );
OR2x2_ASAP7_75t_L g315 ( .A(n_145), .B(n_222), .Y(n_315) );
AND2x2_ASAP7_75t_L g317 ( .A(n_145), .B(n_208), .Y(n_317) );
AND2x2_ASAP7_75t_L g335 ( .A(n_145), .B(n_207), .Y(n_335) );
INVx1_ASAP7_75t_L g368 ( .A(n_145), .Y(n_368) );
INVx2_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
BUFx2_ASAP7_75t_L g235 ( .A(n_146), .Y(n_235) );
AND2x2_ASAP7_75t_L g271 ( .A(n_146), .B(n_208), .Y(n_271) );
AND2x2_ASAP7_75t_L g424 ( .A(n_146), .B(n_222), .Y(n_424) );
AO21x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_154), .B(n_179), .Y(n_146) );
INVx3_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_147), .B(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_147), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_SL g505 ( .A(n_147), .B(n_506), .Y(n_505) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_148), .Y(n_209) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_148), .A2(n_453), .B(n_460), .Y(n_452) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g186 ( .A(n_149), .Y(n_186) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
AND2x2_ASAP7_75t_SL g182 ( .A(n_150), .B(n_151), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_163), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_156), .A2(n_182), .B(n_224), .C(n_225), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_156), .A2(n_242), .B(n_243), .Y(n_241) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_156), .A2(n_178), .B1(n_466), .B2(n_470), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_156), .A2(n_488), .B(n_489), .Y(n_487) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_156), .A2(n_532), .B(n_533), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g156 ( .A(n_157), .B(n_161), .Y(n_156) );
AND2x4_ASAP7_75t_L g190 ( .A(n_157), .B(n_161), .Y(n_190) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_160), .Y(n_157) );
INVx1_ASAP7_75t_L g201 ( .A(n_158), .Y(n_201) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
INVx1_ASAP7_75t_L g268 ( .A(n_159), .Y(n_268) );
INVx1_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_160), .Y(n_171) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_160), .Y(n_173) );
INVx3_ASAP7_75t_L g198 ( .A(n_160), .Y(n_198) );
INVx1_ASAP7_75t_L g457 ( .A(n_160), .Y(n_457) );
INVx4_ASAP7_75t_SL g178 ( .A(n_161), .Y(n_178) );
BUFx3_ASAP7_75t_L g230 ( .A(n_161), .Y(n_230) );
INVx5_ASAP7_75t_L g193 ( .A(n_164), .Y(n_193) );
AND2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
BUFx3_ASAP7_75t_L g176 ( .A(n_165), .Y(n_176) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_165), .Y(n_218) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_172), .C(n_174), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_L g244 ( .A1(n_169), .A2(n_174), .B(n_245), .C(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
OAI22xp5_ASAP7_75t_SL g467 ( .A1(n_170), .A2(n_171), .B1(n_468), .B2(n_469), .Y(n_467) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx4_ASAP7_75t_L g200 ( .A(n_171), .Y(n_200) );
INVx4_ASAP7_75t_L g214 ( .A(n_173), .Y(n_214) );
INVx2_ASAP7_75t_L g255 ( .A(n_173), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_174), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_174), .A2(n_535), .B(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g281 ( .A(n_176), .Y(n_281) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g191 ( .A1(n_178), .A2(n_192), .B(n_193), .C(n_194), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_178), .A2(n_193), .B(n_212), .C(n_213), .Y(n_211) );
O2A1O1Ixp33_ASAP7_75t_SL g252 ( .A1(n_178), .A2(n_193), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g262 ( .A1(n_178), .A2(n_193), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_SL g276 ( .A1(n_178), .A2(n_193), .B(n_277), .C(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g454 ( .A1(n_178), .A2(n_193), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_178), .A2(n_193), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_178), .A2(n_193), .B(n_523), .C(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_181), .A2(n_510), .B(n_517), .Y(n_509) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g240 ( .A(n_182), .Y(n_240) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_182), .A2(n_251), .B(n_258), .Y(n_250) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_182), .A2(n_521), .B(n_527), .Y(n_520) );
AND2x2_ASAP7_75t_L g305 ( .A(n_183), .B(n_206), .Y(n_305) );
OR2x2_ASAP7_75t_L g309 ( .A(n_183), .B(n_222), .Y(n_309) );
AND2x2_ASAP7_75t_L g334 ( .A(n_183), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g381 ( .A(n_183), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_183), .B(n_343), .Y(n_429) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_187), .B(n_202), .Y(n_183) );
INVx1_ASAP7_75t_L g287 ( .A(n_184), .Y(n_287) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_184), .A2(n_531), .B(n_537), .Y(n_530) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_SL g499 ( .A1(n_185), .A2(n_500), .B(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AO21x2_ASAP7_75t_L g464 ( .A1(n_186), .A2(n_465), .B(n_471), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_186), .B(n_472), .Y(n_471) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_186), .A2(n_487), .B(n_494), .Y(n_486) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_188), .A2(n_203), .B(n_287), .Y(n_286) );
BUFx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_195), .B(n_201), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B1(n_199), .B2(n_200), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_197), .A2(n_227), .B(n_228), .C(n_229), .Y(n_226) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_197), .A2(n_491), .B(n_492), .C(n_493), .Y(n_490) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_198), .B(n_257), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_198), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_198), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_200), .B(n_266), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_200), .B(n_280), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_200), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g229 ( .A(n_201), .Y(n_229) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
OAI322xp33_ASAP7_75t_L g430 ( .A1(n_205), .A2(n_366), .A3(n_389), .B1(n_410), .B2(n_431), .C1(n_433), .C2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_206), .B(n_286), .Y(n_433) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_221), .Y(n_206) );
AND2x2_ASAP7_75t_L g234 ( .A(n_207), .B(n_235), .Y(n_234) );
AND2x4_ASAP7_75t_L g302 ( .A(n_207), .B(n_222), .Y(n_302) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g343 ( .A(n_208), .B(n_222), .Y(n_343) );
AND2x2_ASAP7_75t_L g387 ( .A(n_208), .B(n_221), .Y(n_387) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_219), .Y(n_208) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_209), .A2(n_261), .B(n_269), .Y(n_260) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_209), .A2(n_275), .B(n_282), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_214), .B(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_218), .Y(n_515) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_220), .A2(n_474), .B(n_480), .Y(n_473) );
AND2x2_ASAP7_75t_L g270 ( .A(n_221), .B(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g288 ( .A(n_221), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_221), .B(n_317), .Y(n_441) );
INVx3_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g233 ( .A(n_222), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_222), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g355 ( .A(n_222), .B(n_286), .Y(n_355) );
AND2x2_ASAP7_75t_L g382 ( .A(n_222), .B(n_317), .Y(n_382) );
OR2x2_ASAP7_75t_L g438 ( .A(n_222), .B(n_289), .Y(n_438) );
OR2x6_ASAP7_75t_L g222 ( .A(n_223), .B(n_231), .Y(n_222) );
INVx1_ASAP7_75t_SL g324 ( .A(n_233), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_234), .B(n_355), .Y(n_356) );
AND2x2_ASAP7_75t_L g390 ( .A(n_234), .B(n_380), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_234), .B(n_313), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_234), .B(n_435), .Y(n_434) );
OAI31xp33_ASAP7_75t_L g408 ( .A1(n_236), .A2(n_270), .A3(n_409), .B(n_411), .Y(n_408) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_249), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_237), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g391 ( .A(n_237), .B(n_326), .Y(n_391) );
OR2x2_ASAP7_75t_L g398 ( .A(n_237), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g410 ( .A(n_237), .B(n_299), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g344 ( .A(n_238), .B(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g272 ( .A(n_239), .B(n_273), .Y(n_272) );
INVx4_ASAP7_75t_L g293 ( .A(n_239), .Y(n_293) );
AND2x2_ASAP7_75t_L g330 ( .A(n_239), .B(n_274), .Y(n_330) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_247), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_240), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_240), .B(n_518), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_240), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g329 ( .A(n_249), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g399 ( .A(n_249), .Y(n_399) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_259), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_250), .B(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_260), .Y(n_299) );
INVx2_ASAP7_75t_L g319 ( .A(n_250), .Y(n_319) );
AND2x2_ASAP7_75t_L g333 ( .A(n_250), .B(n_260), .Y(n_333) );
AND2x2_ASAP7_75t_L g340 ( .A(n_250), .B(n_296), .Y(n_340) );
BUFx3_ASAP7_75t_L g350 ( .A(n_250), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_250), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g295 ( .A(n_259), .Y(n_295) );
AND2x2_ASAP7_75t_L g303 ( .A(n_259), .B(n_293), .Y(n_303) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_260), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_260), .Y(n_327) );
INVx2_ASAP7_75t_L g493 ( .A(n_267), .Y(n_493) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_SL g310 ( .A(n_271), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_271), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_271), .B(n_380), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g403 ( .A(n_272), .B(n_350), .Y(n_403) );
INVx1_ASAP7_75t_SL g437 ( .A(n_272), .Y(n_437) );
INVx1_ASAP7_75t_SL g345 ( .A(n_273), .Y(n_345) );
INVx1_ASAP7_75t_SL g296 ( .A(n_274), .Y(n_296) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
OR2x2_ASAP7_75t_L g318 ( .A(n_274), .B(n_293), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_274), .B(n_293), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_274), .B(n_322), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B(n_290), .C(n_301), .Y(n_283) );
AOI31xp33_ASAP7_75t_L g400 ( .A1(n_284), .A2(n_401), .A3(n_402), .B(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_L g373 ( .A(n_285), .B(n_302), .Y(n_373) );
BUFx3_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_286), .B(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g349 ( .A(n_286), .B(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_286), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g304 ( .A(n_289), .Y(n_304) );
OAI222xp33_ASAP7_75t_L g413 ( .A1(n_289), .A2(n_414), .B1(n_417), .B2(n_418), .C1(n_419), .C2(n_420), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_297), .Y(n_290) );
INVx1_ASAP7_75t_L g419 ( .A(n_291), .Y(n_419) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_293), .B(n_296), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_293), .B(n_319), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_293), .B(n_294), .Y(n_389) );
INVx1_ASAP7_75t_L g440 ( .A(n_293), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_294), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g442 ( .A(n_294), .Y(n_442) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g322 ( .A(n_295), .Y(n_322) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_296), .Y(n_365) );
AOI32xp33_ASAP7_75t_L g301 ( .A1(n_297), .A2(n_302), .A3(n_303), .B1(n_304), .B2(n_305), .Y(n_301) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_299), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g376 ( .A(n_299), .Y(n_376) );
OR2x2_ASAP7_75t_L g417 ( .A(n_299), .B(n_318), .Y(n_417) );
INVx1_ASAP7_75t_L g353 ( .A(n_300), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_302), .B(n_313), .Y(n_338) );
INVx3_ASAP7_75t_L g347 ( .A(n_302), .Y(n_347) );
AOI322xp5_ASAP7_75t_L g363 ( .A1(n_302), .A2(n_347), .A3(n_364), .B1(n_366), .B2(n_369), .C1(n_373), .C2(n_374), .Y(n_363) );
AND2x2_ASAP7_75t_L g339 ( .A(n_303), .B(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g416 ( .A(n_303), .Y(n_416) );
A2O1A1O1Ixp25_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_311), .C(n_319), .D(n_320), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_307), .B(n_350), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g320 ( .A1(n_309), .A2(n_321), .B1(n_324), .B2(n_325), .C(n_328), .Y(n_320) );
INVx1_ASAP7_75t_SL g435 ( .A(n_309), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_316), .B(n_318), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_313), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI221xp5_ASAP7_75t_SL g405 ( .A1(n_315), .A2(n_399), .B1(n_406), .B2(n_407), .C(n_408), .Y(n_405) );
OAI222xp33_ASAP7_75t_L g436 ( .A1(n_316), .A2(n_437), .B1(n_438), .B2(n_439), .C1(n_441), .C2(n_442), .Y(n_436) );
AND2x2_ASAP7_75t_L g394 ( .A(n_317), .B(n_380), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_317), .A2(n_332), .B(n_379), .Y(n_406) );
INVx1_ASAP7_75t_L g420 ( .A(n_317), .Y(n_420) );
INVx2_ASAP7_75t_SL g323 ( .A(n_318), .Y(n_323) );
AND2x2_ASAP7_75t_L g326 ( .A(n_319), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_SL g360 ( .A(n_322), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_322), .B(n_332), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_323), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_323), .B(n_333), .Y(n_362) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI21xp5_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_331), .B(n_334), .Y(n_328) );
INVx1_ASAP7_75t_SL g346 ( .A(n_330), .Y(n_346) );
AND2x2_ASAP7_75t_L g393 ( .A(n_330), .B(n_376), .Y(n_393) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x2_ASAP7_75t_L g432 ( .A(n_332), .B(n_350), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_333), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_SL g418 ( .A(n_334), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B1(n_341), .B2(n_348), .C(n_351), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B1(n_346), .B2(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g351 ( .A1(n_345), .A2(n_352), .B1(n_354), .B2(n_356), .Y(n_351) );
OR2x2_ASAP7_75t_L g422 ( .A(n_346), .B(n_350), .Y(n_422) );
OR2x2_ASAP7_75t_L g425 ( .A(n_346), .B(n_360), .Y(n_425) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g421 ( .A1(n_367), .A2(n_422), .B1(n_423), .B2(n_425), .C(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND3xp33_ASAP7_75t_SL g377 ( .A(n_378), .B(n_392), .C(n_404), .Y(n_377) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_383), .B1(n_385), .B2(n_388), .C1(n_390), .C2(n_391), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_382), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_380), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g402 ( .A(n_382), .Y(n_402) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_395), .B2(n_397), .C(n_400), .Y(n_392) );
INVx1_ASAP7_75t_L g407 ( .A(n_393), .Y(n_407) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI21xp33_ASAP7_75t_L g426 ( .A1(n_397), .A2(n_427), .B(n_428), .Y(n_426) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
NOR5xp2_ASAP7_75t_L g404 ( .A(n_405), .B(n_413), .C(n_421), .D(n_430), .E(n_436), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp5_ASAP7_75t_SL g729 ( .A1(n_443), .A2(n_445), .B1(n_726), .B2(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_663), .Y(n_445) );
NOR4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_593), .C(n_624), .D(n_643), .Y(n_446) );
NAND4xp25_ASAP7_75t_L g447 ( .A(n_448), .B(n_551), .C(n_566), .D(n_584), .Y(n_447) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_496), .B1(n_528), .B2(n_539), .C1(n_544), .C2(n_546), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_481), .Y(n_449) );
INVx1_ASAP7_75t_L g607 ( .A(n_450), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_461), .Y(n_450) );
AND2x2_ASAP7_75t_L g482 ( .A(n_451), .B(n_473), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_451), .B(n_485), .Y(n_636) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g543 ( .A(n_452), .B(n_463), .Y(n_543) );
AND2x2_ASAP7_75t_L g552 ( .A(n_452), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g578 ( .A(n_452), .Y(n_578) );
AND2x2_ASAP7_75t_L g599 ( .A(n_452), .B(n_463), .Y(n_599) );
BUFx2_ASAP7_75t_L g622 ( .A(n_452), .Y(n_622) );
AND2x2_ASAP7_75t_L g646 ( .A(n_452), .B(n_464), .Y(n_646) );
AND2x2_ASAP7_75t_L g710 ( .A(n_452), .B(n_473), .Y(n_710) );
AND2x2_ASAP7_75t_L g611 ( .A(n_461), .B(n_542), .Y(n_611) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_462), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
OR2x2_ASAP7_75t_L g571 ( .A(n_463), .B(n_486), .Y(n_571) );
AND2x2_ASAP7_75t_L g583 ( .A(n_463), .B(n_542), .Y(n_583) );
BUFx2_ASAP7_75t_L g715 ( .A(n_463), .Y(n_715) );
INVx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g484 ( .A(n_464), .B(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g565 ( .A(n_464), .B(n_486), .Y(n_565) );
AND2x2_ASAP7_75t_L g618 ( .A(n_464), .B(n_473), .Y(n_618) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_464), .Y(n_654) );
AND2x2_ASAP7_75t_L g541 ( .A(n_473), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_SL g553 ( .A(n_473), .Y(n_553) );
INVx2_ASAP7_75t_L g564 ( .A(n_473), .Y(n_564) );
BUFx2_ASAP7_75t_L g588 ( .A(n_473), .Y(n_588) );
AND2x2_ASAP7_75t_SL g645 ( .A(n_473), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
AOI332xp33_ASAP7_75t_L g566 ( .A1(n_482), .A2(n_567), .A3(n_571), .B1(n_572), .B2(n_576), .B3(n_579), .C1(n_580), .C2(n_582), .Y(n_566) );
NAND2x1_ASAP7_75t_L g651 ( .A(n_482), .B(n_542), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_482), .B(n_556), .Y(n_702) );
A2O1A1Ixp33_ASAP7_75t_SL g584 ( .A1(n_483), .A2(n_585), .B(n_588), .C(n_589), .Y(n_584) );
AND2x2_ASAP7_75t_L g723 ( .A(n_483), .B(n_564), .Y(n_723) );
INVx3_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
OR2x2_ASAP7_75t_L g620 ( .A(n_484), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g625 ( .A(n_484), .B(n_622), .Y(n_625) );
INVx1_ASAP7_75t_L g556 ( .A(n_485), .Y(n_556) );
AND2x2_ASAP7_75t_L g659 ( .A(n_485), .B(n_618), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_485), .B(n_599), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_485), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_485), .B(n_577), .Y(n_685) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g542 ( .A(n_486), .Y(n_542) );
OAI31xp33_ASAP7_75t_L g724 ( .A1(n_496), .A2(n_645), .A3(n_652), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
AND2x2_ASAP7_75t_L g528 ( .A(n_497), .B(n_529), .Y(n_528) );
NAND2x1_ASAP7_75t_SL g547 ( .A(n_497), .B(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_497), .Y(n_634) );
AND2x2_ASAP7_75t_L g639 ( .A(n_497), .B(n_550), .Y(n_639) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_498), .A2(n_552), .B(n_554), .C(n_557), .Y(n_551) );
OR2x2_ASAP7_75t_L g568 ( .A(n_498), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g581 ( .A(n_498), .Y(n_581) );
AND2x2_ASAP7_75t_L g587 ( .A(n_498), .B(n_530), .Y(n_587) );
INVx2_ASAP7_75t_L g605 ( .A(n_498), .Y(n_605) );
AND2x2_ASAP7_75t_L g616 ( .A(n_498), .B(n_570), .Y(n_616) );
AND2x2_ASAP7_75t_L g648 ( .A(n_498), .B(n_606), .Y(n_648) );
AND2x2_ASAP7_75t_L g652 ( .A(n_498), .B(n_575), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_498), .B(n_507), .Y(n_657) );
AND2x2_ASAP7_75t_L g691 ( .A(n_498), .B(n_692), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_498), .B(n_594), .Y(n_725) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_507), .B(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g633 ( .A(n_507), .Y(n_633) );
AND2x2_ASAP7_75t_L g695 ( .A(n_507), .B(n_616), .Y(n_695) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_519), .Y(n_507) );
OR2x2_ASAP7_75t_L g549 ( .A(n_508), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g559 ( .A(n_508), .B(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_508), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g667 ( .A(n_508), .Y(n_667) );
AND2x2_ASAP7_75t_L g684 ( .A(n_508), .B(n_530), .Y(n_684) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g575 ( .A(n_509), .B(n_519), .Y(n_575) );
AND2x2_ASAP7_75t_L g604 ( .A(n_509), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g615 ( .A(n_509), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_509), .B(n_570), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_516), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g529 ( .A(n_520), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g550 ( .A(n_520), .Y(n_550) );
AND2x2_ASAP7_75t_L g606 ( .A(n_520), .B(n_570), .Y(n_606) );
INVx1_ASAP7_75t_L g708 ( .A(n_528), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_529), .Y(n_712) );
INVx2_ASAP7_75t_L g570 ( .A(n_530), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_541), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_541), .B(n_646), .Y(n_704) );
OR2x2_ASAP7_75t_L g545 ( .A(n_542), .B(n_543), .Y(n_545) );
INVx1_ASAP7_75t_SL g597 ( .A(n_542), .Y(n_597) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_548), .A2(n_601), .B1(n_603), .B2(n_607), .C(n_608), .Y(n_600) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g628 ( .A(n_549), .B(n_592), .Y(n_628) );
INVx2_ASAP7_75t_L g560 ( .A(n_550), .Y(n_560) );
INVx1_ASAP7_75t_L g586 ( .A(n_550), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_550), .B(n_570), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_550), .B(n_573), .Y(n_680) );
INVx1_ASAP7_75t_L g688 ( .A(n_550), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_552), .B(n_556), .Y(n_602) );
AND2x4_ASAP7_75t_L g577 ( .A(n_553), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g690 ( .A(n_556), .B(n_646), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_559), .B(n_591), .Y(n_590) );
INVxp67_ASAP7_75t_L g698 ( .A(n_560), .Y(n_698) );
INVxp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g598 ( .A(n_564), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g670 ( .A(n_564), .B(n_646), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_564), .B(n_583), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_565), .A2(n_599), .A3(n_606), .B1(n_631), .B2(n_634), .C1(n_635), .C2(n_637), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_565), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g696 ( .A(n_568), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g642 ( .A(n_569), .Y(n_642) );
INVx2_ASAP7_75t_L g573 ( .A(n_570), .Y(n_573) );
INVx1_ASAP7_75t_L g632 ( .A(n_570), .Y(n_632) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_571), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g668 ( .A(n_573), .B(n_581), .Y(n_668) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g580 ( .A(n_575), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g623 ( .A(n_575), .B(n_616), .Y(n_623) );
AND2x2_ASAP7_75t_L g627 ( .A(n_575), .B(n_587), .Y(n_627) );
OAI21xp33_ASAP7_75t_SL g637 ( .A1(n_576), .A2(n_638), .B(n_640), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g707 ( .A1(n_576), .A2(n_708), .B1(n_709), .B2(n_711), .Y(n_707) );
INVx3_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g582 ( .A(n_577), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_577), .B(n_597), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_579), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g719 ( .A(n_586), .Y(n_719) );
INVx4_ASAP7_75t_L g592 ( .A(n_587), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_587), .B(n_614), .Y(n_662) );
INVx1_ASAP7_75t_SL g674 ( .A(n_588), .Y(n_674) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp67_ASAP7_75t_L g687 ( .A(n_592), .B(n_688), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_595), .B(n_600), .C(n_617), .Y(n_593) );
OAI221xp5_ASAP7_75t_SL g713 ( .A1(n_595), .A2(n_633), .B1(n_712), .B2(n_714), .C(n_716), .Y(n_713) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_597), .B(n_710), .Y(n_709) );
OAI31xp33_ASAP7_75t_L g689 ( .A1(n_598), .A2(n_675), .A3(n_690), .B(n_691), .Y(n_689) );
INVx1_ASAP7_75t_L g629 ( .A(n_599), .Y(n_629) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g679 ( .A(n_604), .Y(n_679) );
AND2x2_ASAP7_75t_L g692 ( .A(n_606), .B(n_615), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_612), .Y(n_608) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVxp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_616), .B(n_719), .Y(n_718) );
OAI21xp33_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_619), .B(n_623), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B1(n_628), .B2(n_629), .C(n_630), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g693 ( .A1(n_625), .A2(n_694), .B(n_696), .C(n_699), .Y(n_693) );
CKINVDCx16_ASAP7_75t_R g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_628), .B(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx1_ASAP7_75t_L g655 ( .A(n_636), .Y(n_655) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g641 ( .A(n_639), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g683 ( .A(n_639), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_647), .B(n_649), .C(n_658), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g720 ( .A1(n_647), .A2(n_657), .B1(n_721), .B2(n_722), .C(n_724), .Y(n_720) );
INVx1_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_653), .B2(n_656), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g658 ( .A1(n_659), .A2(n_660), .B(n_661), .Y(n_658) );
INVx1_ASAP7_75t_SL g721 ( .A(n_660), .Y(n_721) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR4xp25_ASAP7_75t_L g663 ( .A(n_664), .B(n_693), .C(n_713), .D(n_720), .Y(n_663) );
OAI211xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_669), .B(n_671), .C(n_689), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_668), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_675), .B(n_677), .C(n_681), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g700 ( .A(n_678), .Y(n_700) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
OR2x2_ASAP7_75t_L g711 ( .A(n_679), .B(n_712), .Y(n_711) );
OAI21xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B(n_686), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_701), .B1(n_703), .B2(n_705), .C(n_707), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_710), .B(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_738), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
endmodule