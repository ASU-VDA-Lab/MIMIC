module fake_jpeg_21686_n_192 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_1),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_56),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_25),
.B1(n_26),
.B2(n_15),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_52),
.B1(n_16),
.B2(n_14),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_25),
.B1(n_15),
.B2(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_23),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_17),
.B1(n_2),
.B2(n_3),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_28),
.B1(n_16),
.B2(n_14),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_41),
.B1(n_32),
.B2(n_35),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_45),
.B(n_40),
.Y(n_66)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_96),
.A3(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_76),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_62),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_77),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_89),
.Y(n_99)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_80),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_22),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_30),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_87),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_27),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

OR2x4_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_32),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_93),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_35),
.B1(n_39),
.B2(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_91),
.A2(n_94),
.B1(n_49),
.B2(n_34),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_39),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_39),
.B1(n_34),
.B2(n_33),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_31),
.B1(n_44),
.B2(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_31),
.B1(n_64),
.B2(n_4),
.Y(n_106)
);

AO22x2_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_94),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_67),
.C(n_77),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_93),
.C(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_82),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_79),
.Y(n_121)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_66),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_125),
.C(n_102),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_133),
.B1(n_134),
.B2(n_80),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_101),
.B1(n_106),
.B2(n_99),
.Y(n_146)
);

CKINVDCx10_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_76),
.C(n_111),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_74),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_103),
.B1(n_108),
.B2(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_143),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_111),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_116),
.Y(n_144)
);

OAI322xp33_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_124),
.A3(n_107),
.B1(n_126),
.B2(n_128),
.C1(n_133),
.C2(n_118),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_116),
.C(n_114),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_132),
.C(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_148),
.B(n_104),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_144),
.Y(n_167)
);

OA21x2_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_130),
.B(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_154),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_107),
.B(n_97),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_159),
.A2(n_161),
.B1(n_146),
.B2(n_107),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_83),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_75),
.C(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_164),
.B(n_165),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_167),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_170),
.B(n_152),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_156),
.C(n_157),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_162),
.C(n_169),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_157),
.B1(n_152),
.B2(n_156),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_177),
.B1(n_6),
.B2(n_7),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_169),
.A2(n_158),
.B1(n_150),
.B2(n_78),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_168),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_179),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_171),
.C(n_172),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_181),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_9),
.B(n_12),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_6),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_178),
.B(n_9),
.Y(n_186)
);

AO21x1_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_183),
.B(n_7),
.Y(n_189)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_187),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_188),
.B(n_75),
.Y(n_191)
);

BUFx24_ASAP7_75t_SL g192 ( 
.A(n_191),
.Y(n_192)
);


endmodule