module fake_jpeg_13207_n_349 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_44),
.Y(n_123)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_45),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_50),
.Y(n_82)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_18),
.B(n_14),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_54),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_13),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_13),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_68),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_61),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_24),
.B(n_11),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_69),
.B(n_71),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_70),
.Y(n_110)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_73),
.Y(n_100)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_74),
.B(n_75),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_38),
.B1(n_20),
.B2(n_19),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_76),
.A2(n_87),
.B1(n_83),
.B2(n_119),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_38),
.B1(n_35),
.B2(n_20),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_77),
.A2(n_78),
.B1(n_89),
.B2(n_83),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_35),
.B1(n_25),
.B2(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_36),
.B1(n_16),
.B2(n_39),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_43),
.A2(n_36),
.B1(n_16),
.B2(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_16),
.B1(n_34),
.B2(n_15),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_16),
.B1(n_34),
.B2(n_15),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_55),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_30),
.B1(n_28),
.B2(n_40),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_88),
.B(n_98),
.C(n_115),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_46),
.A2(n_26),
.B1(n_25),
.B2(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_29),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_96),
.B(n_102),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_40),
.B1(n_22),
.B2(n_11),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_0),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_107),
.B1(n_112),
.B2(n_126),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_11),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_109),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_45),
.B(n_0),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_67),
.B(n_5),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_5),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_60),
.B(n_5),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_102),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_44),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_128),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_66),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_68),
.A2(n_7),
.B1(n_9),
.B2(n_71),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_127),
.A2(n_129),
.B1(n_123),
.B2(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_9),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_65),
.A2(n_9),
.B1(n_23),
.B2(n_33),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_130),
.B(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_125),
.C(n_106),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_147),
.Y(n_189)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_148),
.Y(n_183)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_89),
.B1(n_96),
.B2(n_77),
.Y(n_141)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_113),
.B(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_142),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_87),
.A2(n_98),
.B1(n_88),
.B2(n_83),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_144),
.A2(n_145),
.B1(n_157),
.B2(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_146),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_125),
.C(n_121),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_82),
.B(n_91),
.C(n_118),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_149),
.A2(n_175),
.B(n_152),
.C(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_156),
.Y(n_198)
);

BUFx4f_ASAP7_75t_SL g152 ( 
.A(n_110),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_152),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_154),
.B1(n_161),
.B2(n_166),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_78),
.A2(n_95),
.B1(n_114),
.B2(n_92),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_111),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_158),
.B(n_160),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_163),
.Y(n_199)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_84),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_116),
.A2(n_118),
.B1(n_105),
.B2(n_95),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_93),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_165),
.Y(n_204)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_92),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_168),
.B(n_171),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_110),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_175),
.B(n_172),
.Y(n_192)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_122),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_172),
.Y(n_179)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_174),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_81),
.Y(n_175)
);

NOR2x1_ASAP7_75t_R g203 ( 
.A(n_177),
.B(n_133),
.Y(n_203)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_187),
.B(n_190),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_177),
.A2(n_137),
.B(n_141),
.C(n_153),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_196),
.Y(n_218)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_149),
.A3(n_162),
.B1(n_143),
.B2(n_176),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_206),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_179),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_147),
.A2(n_150),
.B1(n_132),
.B2(n_165),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g245 ( 
.A(n_201),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_189),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_205),
.A2(n_208),
.B1(n_195),
.B2(n_214),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_139),
.B(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_210),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_160),
.A2(n_167),
.B1(n_159),
.B2(n_135),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_152),
.B(n_158),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_181),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_148),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_156),
.B(n_130),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_201),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_147),
.B(n_169),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_214),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_144),
.A2(n_145),
.B1(n_157),
.B2(n_153),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_205),
.B1(n_188),
.B2(n_184),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_217),
.B(n_178),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_211),
.B(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_219),
.A2(n_226),
.B1(n_235),
.B2(n_237),
.Y(n_271)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_223),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_191),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_215),
.A2(n_182),
.B1(n_203),
.B2(n_184),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_229),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_200),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_194),
.B(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_198),
.B(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_232),
.B(n_236),
.Y(n_257)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_233),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_186),
.Y(n_234)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_202),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_180),
.A2(n_210),
.B1(n_199),
.B2(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_240),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_195),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_241),
.B(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_237),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_246),
.Y(n_264)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_269),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_266),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_255),
.B(n_261),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_178),
.B(n_228),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_260),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_218),
.A2(n_228),
.B(n_245),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_225),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_220),
.B1(n_230),
.B2(n_222),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_242),
.Y(n_266)
);

OAI22x1_ASAP7_75t_L g269 ( 
.A1(n_216),
.A2(n_226),
.B1(n_223),
.B2(n_243),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_272),
.B(n_275),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_273),
.A2(n_266),
.B1(n_267),
.B2(n_248),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_280),
.C(n_289),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_225),
.B1(n_222),
.B2(n_241),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_286),
.B1(n_287),
.B2(n_290),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_251),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_279),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_238),
.C(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_252),
.B(n_246),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_284),
.Y(n_303)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_250),
.B(n_251),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_292),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_221),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_268),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_269),
.C(n_259),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_296),
.B(n_308),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_254),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_298),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_269),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_258),
.A3(n_262),
.B1(n_255),
.B2(n_267),
.C1(n_271),
.C2(n_254),
.Y(n_300)
);

OAI322xp33_ASAP7_75t_L g310 ( 
.A1(n_300),
.A2(n_274),
.A3(n_288),
.B1(n_276),
.B2(n_247),
.C1(n_264),
.C2(n_285),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_273),
.A2(n_271),
.B1(n_248),
.B2(n_264),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_270),
.C(n_260),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_275),
.Y(n_309)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_309),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_310),
.A2(n_318),
.B1(n_322),
.B2(n_240),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_284),
.B(n_291),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_311),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_272),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_314),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_279),
.B1(n_274),
.B2(n_284),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_316),
.B1(n_319),
.B2(n_303),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_247),
.B1(n_270),
.B2(n_260),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_268),
.Y(n_318)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_260),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_320),
.B(n_293),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_282),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_295),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_233),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_324),
.Y(n_336)
);

OAI21x1_ASAP7_75t_SL g333 ( 
.A1(n_325),
.A2(n_332),
.B(n_320),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_321),
.B(n_298),
.C(n_308),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_327),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_296),
.C(n_293),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_304),
.B1(n_301),
.B2(n_299),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_331),
.A2(n_317),
.B1(n_304),
.B2(n_301),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_333),
.B(n_338),
.Y(n_340)
);

A2O1A1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_329),
.A2(n_310),
.B(n_311),
.C(n_316),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_337),
.C(n_328),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_329),
.A2(n_312),
.B(n_320),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_342),
.B(n_327),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_336),
.B(n_330),
.Y(n_341)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_341),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_334),
.B(n_317),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_340),
.B(n_335),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_326),
.C(n_323),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_345),
.C(n_324),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_313),
.Y(n_349)
);


endmodule