module fake_jpeg_20648_n_232 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_32),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_14),
.B1(n_24),
.B2(n_18),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_15),
.B1(n_24),
.B2(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_14),
.B1(n_24),
.B2(n_20),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_40),
.B1(n_46),
.B2(n_34),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_20),
.B1(n_14),
.B2(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_26),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_50),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_26),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_58),
.Y(n_72)
);

AO22x2_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_39),
.B1(n_33),
.B2(n_37),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_54),
.B1(n_57),
.B2(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_33),
.B1(n_30),
.B2(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_48),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_33),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_65),
.C(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_27),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_47),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_64),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_45),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_51),
.B(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_37),
.B1(n_45),
.B2(n_44),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_70),
.A2(n_73),
.B1(n_75),
.B2(n_81),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_37),
.B1(n_45),
.B2(n_30),
.Y(n_75)
);

OAI32xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_30),
.A3(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_27),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_43),
.B1(n_15),
.B2(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_28),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_28),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_84),
.Y(n_95)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_52),
.B1(n_63),
.B2(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_78),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_90),
.B(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_92),
.B(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_52),
.B1(n_66),
.B2(n_59),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_102),
.B1(n_67),
.B2(n_84),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_76),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_52),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_61),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_25),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_67),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_21),
.B1(n_16),
.B2(n_19),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_67),
.B(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_110),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_98),
.B1(n_104),
.B2(n_112),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_71),
.C(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_108),
.C(n_95),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_74),
.C(n_79),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_75),
.B1(n_82),
.B2(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_69),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_113),
.B(n_118),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_117),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_84),
.B(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_80),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_87),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_111),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_128),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_87),
.B(n_86),
.Y(n_123)
);

AO21x2_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_86),
.B(n_106),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_91),
.B(n_1),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_99),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_132),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_108),
.C(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_140),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_136),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_86),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_103),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_109),
.B(n_18),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_151),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_114),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_132),
.B(n_86),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_140),
.A2(n_141),
.B1(n_124),
.B2(n_139),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_150),
.B1(n_159),
.B2(n_152),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_91),
.B1(n_109),
.B2(n_85),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_127),
.A2(n_123),
.B(n_136),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_158),
.B(n_16),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_7),
.B(n_11),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_85),
.B1(n_16),
.B2(n_13),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_160),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_126),
.B1(n_134),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_166),
.B1(n_167),
.B2(n_143),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_135),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_143),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_135),
.C(n_131),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_145),
.C(n_142),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_123),
.B1(n_125),
.B2(n_122),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_125),
.B1(n_43),
.B2(n_15),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_160),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_168),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_174),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_155),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_177),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_22),
.C(n_17),
.Y(n_196)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_148),
.A3(n_167),
.B1(n_144),
.B2(n_170),
.C(n_172),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_188),
.B(n_10),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_187),
.Y(n_193)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_143),
.A3(n_149),
.B1(n_157),
.B2(n_35),
.C1(n_22),
.C2(n_25),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_164),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_186),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_162),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

AO221x1_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_166),
.B1(n_22),
.B2(n_43),
.C(n_29),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_197),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_163),
.B(n_10),
.Y(n_194)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_194),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_198),
.C(n_22),
.Y(n_207)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_29),
.B(n_28),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_186),
.C(n_184),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_181),
.A2(n_9),
.B(n_10),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_8),
.B(n_12),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_189),
.C(n_185),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_195),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_8),
.Y(n_204)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_204),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_197),
.C(n_35),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_7),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_209),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_193),
.A2(n_29),
.B1(n_9),
.B2(n_15),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_215),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_198),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_207),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_213),
.A2(n_201),
.B1(n_35),
.B2(n_2),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_197),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_9),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_4),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_206),
.B(n_0),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_211),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_218),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_223),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_222),
.B(n_217),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_0),
.C(n_1),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_226),
.Y(n_228)
);

AOI321xp33_ASAP7_75t_L g227 ( 
.A1(n_225),
.A2(n_220),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_227),
.A2(n_224),
.B(n_1),
.Y(n_229)
);

OAI321xp33_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_0),
.A3(n_2),
.B1(n_3),
.B2(n_228),
.C(n_202),
.Y(n_230)
);

NOR2xp67_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_0),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_3),
.Y(n_232)
);


endmodule