module fake_jpeg_28563_n_35 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_8),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_3),
.B(n_0),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_7),
.A2(n_2),
.B(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_11),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_11),
.A2(n_1),
.B1(n_9),
.B2(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

AO221x1_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_27),
.B1(n_14),
.B2(n_10),
.C(n_23),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_17),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_23),
.C(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

OAI321xp33_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_25),
.A3(n_15),
.B1(n_8),
.B2(n_6),
.C(n_4),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_28),
.A3(n_25),
.B1(n_30),
.B2(n_15),
.C1(n_12),
.C2(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_34),
.B1(n_10),
.B2(n_27),
.Y(n_35)
);


endmodule