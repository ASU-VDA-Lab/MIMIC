module fake_ariane_2613_n_712 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_712);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_712;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_367;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_264;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_354;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_500;
wire n_665;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_672;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_222;
wire n_703;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_491;
wire n_181;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_452;
wire n_217;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_212;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_378;
wire n_203;
wire n_436;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_0),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_11),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_142),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_88),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_27),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_105),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_119),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_22),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_100),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_114),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g171 ( 
.A(n_127),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_51),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_42),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_59),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_69),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_10),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_99),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_40),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_33),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_73),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_116),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_47),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_139),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_35),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_96),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_72),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_102),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_83),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_58),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_132),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_56),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_75),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_84),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_4),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_57),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_91),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_65),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_86),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_104),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_26),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_38),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_93),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_126),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_39),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_16),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_44),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_82),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_54),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_61),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_95),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_48),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_28),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_21),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_49),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_5),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_120),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_20),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_146),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_115),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_98),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_19),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_101),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_62),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_150),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_85),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_18),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_13),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_24),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_89),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_45),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_23),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_97),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_230),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_179),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_230),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_190),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_183),
.B(n_153),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_204),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_154),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_210),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_155),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_246),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_224),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_254),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_R g273 ( 
.A(n_232),
.B(n_25),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_167),
.Y(n_274)
);

BUFx6f_ASAP7_75t_SL g275 ( 
.A(n_161),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_157),
.B(n_1),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_200),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_209),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_159),
.B(n_1),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_163),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_163),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_174),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_166),
.B(n_2),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_180),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_180),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

BUFx6f_ASAP7_75t_SL g289 ( 
.A(n_160),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_172),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_175),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_239),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_189),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_176),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_177),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_184),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_202),
.Y(n_298)
);

NOR2xp67_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_3),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_236),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_227),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_198),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_251),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_158),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_162),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_201),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_207),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_164),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_208),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_211),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_219),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_221),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_231),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_169),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_237),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_240),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_185),
.Y(n_327)
);

OA21x2_ASAP7_75t_L g328 ( 
.A1(n_264),
.A2(n_182),
.B(n_165),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_156),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_297),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_327),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_276),
.A2(n_194),
.B(n_182),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_327),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_256),
.Y(n_342)
);

OA21x2_ASAP7_75t_L g343 ( 
.A1(n_290),
.A2(n_216),
.B(n_194),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_259),
.A2(n_187),
.B1(n_191),
.B2(n_168),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_193),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_277),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_311),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_255),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_291),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_257),
.B(n_214),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_263),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_L g356 ( 
.A(n_273),
.B(n_185),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_310),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_L g360 ( 
.A(n_313),
.B(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_300),
.B(n_171),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_315),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_325),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_320),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_274),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_262),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_282),
.B(n_283),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_324),
.Y(n_374)
);

OA21x2_ASAP7_75t_L g375 ( 
.A1(n_326),
.A2(n_233),
.B(n_218),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_284),
.B(n_218),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_266),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_281),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_285),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_316),
.B(n_206),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_289),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

BUFx4f_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_378),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_378),
.B(n_308),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_364),
.B(n_309),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_333),
.B(n_286),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_342),
.Y(n_398)
);

AND2x6_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_244),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_364),
.B(n_312),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_331),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_334),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_332),
.B(n_336),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_287),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_365),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_352),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_323),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_342),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_368),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_375),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_288),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_331),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_374),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_362),
.B(n_278),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_345),
.B(n_280),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_372),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_377),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_349),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_372),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_381),
.A2(n_293),
.B1(n_307),
.B2(n_298),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_346),
.B(n_244),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_371),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_420),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_434),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_403),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_348),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_398),
.B(n_353),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_348),
.Y(n_447)
);

AND2x6_ASAP7_75t_L g448 ( 
.A(n_404),
.B(n_245),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_410),
.B(n_382),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_436),
.A2(n_339),
.B1(n_328),
.B2(n_356),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_355),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g453 ( 
.A1(n_426),
.A2(n_265),
.B1(n_270),
.B2(n_269),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_385),
.Y(n_454)
);

NOR2xp67_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_267),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_437),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_395),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_385),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_432),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_358),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_396),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_400),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_406),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_407),
.Y(n_471)
);

AO22x2_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_272),
.B1(n_271),
.B2(n_363),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_411),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_390),
.B(n_370),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_397),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_386),
.Y(n_478)
);

NAND2x1p5_ASAP7_75t_L g479 ( 
.A(n_409),
.B(n_369),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_414),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_424),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_415),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_415),
.Y(n_483)
);

NAND2x1p5_ASAP7_75t_L g484 ( 
.A(n_416),
.B(n_361),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_435),
.A2(n_292),
.B1(n_367),
.B2(n_366),
.Y(n_486)
);

OAI221xp5_ASAP7_75t_L g487 ( 
.A1(n_425),
.A2(n_299),
.B1(n_401),
.B2(n_391),
.C(n_431),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_390),
.A2(n_178),
.B1(n_170),
.B2(n_360),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_417),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_449),
.B(n_423),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_447),
.B(n_419),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_452),
.B(n_454),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_419),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_462),
.B(n_393),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_455),
.B(n_408),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_440),
.B(n_399),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_440),
.B(n_445),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_475),
.B(n_402),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_443),
.B(n_399),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_488),
.B(n_402),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_SL g502 ( 
.A(n_446),
.B(n_275),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_442),
.B(n_438),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_444),
.B(n_422),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_458),
.B(n_173),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_450),
.B(n_418),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_SL g507 ( 
.A(n_441),
.B(n_289),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_459),
.B(n_186),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_484),
.B(n_489),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_486),
.B(n_188),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_SL g511 ( 
.A(n_478),
.B(n_192),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_479),
.B(n_195),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_463),
.B(n_245),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_451),
.B(n_247),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_464),
.B(n_196),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_465),
.B(n_197),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_470),
.B(n_199),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_487),
.B(n_203),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_461),
.B(n_456),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_480),
.B(n_212),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_481),
.B(n_215),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_467),
.B(n_468),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_469),
.B(n_471),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_473),
.B(n_217),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_460),
.B(n_220),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_SL g526 ( 
.A(n_457),
.B(n_222),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_498),
.A2(n_483),
.B(n_482),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_492),
.Y(n_528)
);

AO31x2_ASAP7_75t_L g529 ( 
.A1(n_506),
.A2(n_490),
.A3(n_485),
.B(n_476),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_497),
.A2(n_477),
.B(n_474),
.Y(n_530)
);

O2A1O1Ixp33_ASAP7_75t_SL g531 ( 
.A1(n_491),
.A2(n_247),
.B(n_448),
.C(n_338),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_519),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_522),
.A2(n_472),
.B(n_448),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_494),
.B(n_448),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_500),
.B(n_453),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_523),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_513),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_507),
.Y(n_538)
);

AO31x2_ASAP7_75t_L g539 ( 
.A1(n_518),
.A2(n_514),
.A3(n_525),
.B(n_508),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_504),
.B(n_6),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_493),
.B(n_7),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_510),
.B(n_8),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_496),
.B(n_8),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_502),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_503),
.B(n_13),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_501),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_509),
.B(n_229),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_14),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_512),
.A2(n_30),
.B(n_29),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_524),
.B(n_15),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_526),
.B(n_15),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_517),
.A2(n_32),
.B(n_31),
.Y(n_554)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_511),
.B(n_341),
.C(n_340),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_515),
.Y(n_556)
);

BUFx2_ASAP7_75t_R g557 ( 
.A(n_516),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_533),
.A2(n_521),
.B(n_520),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_538),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_532),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g561 ( 
.A1(n_527),
.A2(n_37),
.B(n_36),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_528),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_536),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_537),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_544),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g566 ( 
.A1(n_530),
.A2(n_90),
.B(n_152),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_543),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_546),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_548),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

AOI221xp5_ASAP7_75t_L g572 ( 
.A1(n_542),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.C(n_50),
.Y(n_572)
);

AO21x2_ASAP7_75t_L g573 ( 
.A1(n_534),
.A2(n_53),
.B(n_55),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_556),
.Y(n_574)
);

INVx1_ASAP7_75t_SL g575 ( 
.A(n_547),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_552),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_547),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_545),
.A2(n_553),
.B1(n_541),
.B2(n_549),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_550),
.B(n_557),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_554),
.A2(n_68),
.B(n_70),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_531),
.A2(n_71),
.B(n_74),
.Y(n_582)
);

OR2x6_ASAP7_75t_L g583 ( 
.A(n_535),
.B(n_77),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_529),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_551),
.Y(n_585)
);

OA21x2_ASAP7_75t_L g586 ( 
.A1(n_555),
.A2(n_78),
.B(n_80),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_584),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_562),
.B(n_539),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_571),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_563),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_565),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_568),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_570),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_585),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_577),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_578),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_566),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_573),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_567),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_586),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_559),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_564),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_564),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_569),
.Y(n_607)
);

OR2x2_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_145),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_580),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_581),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_560),
.B(n_81),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_582),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_106),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_607),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_590),
.Y(n_617)
);

BUFx10_ASAP7_75t_L g618 ( 
.A(n_609),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_590),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_599),
.B(n_579),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_609),
.B(n_601),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_591),
.Y(n_622)
);

OR2x6_ASAP7_75t_L g623 ( 
.A(n_614),
.B(n_576),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_601),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g625 ( 
.A(n_595),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_602),
.B(n_576),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_592),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_592),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_596),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_596),
.B(n_561),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_613),
.B(n_109),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_615),
.B(n_572),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_615),
.B(n_110),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_588),
.B(n_111),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_587),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_605),
.B(n_117),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_593),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_606),
.Y(n_639)
);

CKINVDCx11_ASAP7_75t_R g640 ( 
.A(n_611),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_635),
.B(n_594),
.Y(n_641)
);

NOR2x1_ASAP7_75t_SL g642 ( 
.A(n_623),
.B(n_626),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_625),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_620),
.B(n_593),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_617),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_619),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_622),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_624),
.B(n_608),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_638),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_627),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_639),
.B(n_604),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_598),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_629),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_628),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_636),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_634),
.B(n_589),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_640),
.B(n_600),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_630),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_621),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_631),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_618),
.B(n_597),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_637),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_643),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_653),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_652),
.B(n_612),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_645),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_659),
.B(n_616),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_650),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_654),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_645),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_649),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_649),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_646),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_661),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_647),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_657),
.B(n_610),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_674),
.B(n_642),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_663),
.B(n_641),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_666),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_666),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_670),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_671),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_676),
.B(n_664),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_677),
.Y(n_684)
);

AO221x2_ASAP7_75t_L g685 ( 
.A1(n_678),
.A2(n_667),
.B1(n_672),
.B2(n_673),
.C(n_648),
.Y(n_685)
);

AO221x2_ASAP7_75t_L g686 ( 
.A1(n_679),
.A2(n_675),
.B1(n_658),
.B2(n_660),
.C(n_662),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_680),
.Y(n_687)
);

AO221x2_ASAP7_75t_L g688 ( 
.A1(n_681),
.A2(n_655),
.B1(n_644),
.B2(n_668),
.C(n_669),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_687),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_685),
.B(n_682),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_684),
.B(n_683),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_686),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_688),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_689),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_690),
.A2(n_693),
.B(n_692),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_691),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_694),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_697),
.B(n_695),
.Y(n_698)
);

NOR2x1_ASAP7_75t_L g699 ( 
.A(n_698),
.B(n_696),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_699),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_700),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_R g702 ( 
.A(n_701),
.B(n_121),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_702),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_703),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_704),
.Y(n_705)
);

AOI31xp33_ASAP7_75t_L g706 ( 
.A1(n_705),
.A2(n_656),
.A3(n_124),
.B(n_125),
.Y(n_706)
);

INVxp33_ASAP7_75t_L g707 ( 
.A(n_706),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_707),
.Y(n_708)
);

AOI221xp5_ASAP7_75t_L g709 ( 
.A1(n_707),
.A2(n_651),
.B1(n_665),
.B2(n_129),
.C(n_130),
.Y(n_709)
);

INVxp67_ASAP7_75t_SL g710 ( 
.A(n_708),
.Y(n_710)
);

AOI221xp5_ASAP7_75t_L g711 ( 
.A1(n_710),
.A2(n_709),
.B1(n_128),
.B2(n_131),
.C(n_134),
.Y(n_711)
);

AOI211xp5_ASAP7_75t_L g712 ( 
.A1(n_711),
.A2(n_140),
.B(n_141),
.C(n_144),
.Y(n_712)
);


endmodule