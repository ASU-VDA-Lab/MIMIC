module fake_jpeg_29592_n_417 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_417);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_417;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_46),
.B(n_48),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_51),
.B(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_56),
.B(n_80),
.Y(n_132)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_6),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_7),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_70),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_7),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_75),
.B(n_42),
.Y(n_127)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_82),
.B(n_83),
.Y(n_109)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_85),
.Y(n_121)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_86),
.B(n_37),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_52),
.B1(n_63),
.B2(n_68),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_89),
.A2(n_94),
.B1(n_96),
.B2(n_112),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_56),
.A2(n_23),
.B1(n_43),
.B2(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_90),
.A2(n_98),
.B1(n_107),
.B2(n_108),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_34),
.B1(n_43),
.B2(n_30),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_69),
.A2(n_34),
.B1(n_43),
.B2(n_30),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_23),
.B1(n_43),
.B2(n_30),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_53),
.A2(n_23),
.B1(n_34),
.B2(n_22),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_59),
.A2(n_34),
.B1(n_22),
.B2(n_35),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_45),
.A2(n_22),
.B1(n_40),
.B2(n_39),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_48),
.A2(n_39),
.B(n_35),
.C(n_40),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_116),
.A2(n_0),
.B(n_103),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_49),
.A2(n_44),
.B1(n_42),
.B2(n_41),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_31),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_16),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_55),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_16),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_64),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_133),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_65),
.B(n_35),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_48),
.B(n_21),
.C(n_54),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_136),
.Y(n_188)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

BUFx4f_ASAP7_75t_SL g185 ( 
.A(n_137),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_140),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_145),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_87),
.A2(n_71),
.B1(n_85),
.B2(n_73),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_143),
.A2(n_168),
.B1(n_179),
.B2(n_135),
.Y(n_196)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g215 ( 
.A(n_144),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_131),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_91),
.B1(n_130),
.B2(n_125),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_162),
.B1(n_141),
.B2(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_152),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_21),
.B1(n_16),
.B2(n_37),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_104),
.B(n_37),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_54),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_37),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_37),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_160),
.Y(n_192)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_79),
.C(n_21),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_12),
.Y(n_223)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx4_ASAP7_75t_SL g214 ( 
.A(n_158),
.Y(n_214)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_16),
.Y(n_160)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_165),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_103),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_175),
.Y(n_205)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

AO22x1_ASAP7_75t_SL g166 ( 
.A1(n_95),
.A2(n_24),
.B1(n_0),
.B2(n_2),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_166),
.A2(n_181),
.B1(n_122),
.B2(n_114),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_170),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_24),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_171),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_101),
.B(n_7),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_173),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_99),
.B(n_5),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_177),
.Y(n_221)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g176 ( 
.A1(n_105),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_180),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_9),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_9),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_99),
.A2(n_11),
.B1(n_1),
.B2(n_3),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_11),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_111),
.B(n_124),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_184),
.A2(n_209),
.B1(n_212),
.B2(n_217),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_186),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_196),
.Y(n_231)
);

CKINVDCx12_ASAP7_75t_R g195 ( 
.A(n_144),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_195),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_216),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_151),
.B(n_135),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_202),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_138),
.A2(n_120),
.B(n_119),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_199),
.A2(n_203),
.B(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_148),
.B(n_93),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_138),
.A2(n_136),
.B(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_93),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_206),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_153),
.B(n_122),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_120),
.B1(n_92),
.B2(n_119),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_167),
.A2(n_92),
.B1(n_124),
.B2(n_13),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_149),
.A2(n_157),
.B(n_164),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_154),
.B(n_4),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_224),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_166),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_166),
.B(n_14),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_230),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_191),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_191),
.B(n_181),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_232),
.B(n_205),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_233),
.B(n_217),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_188),
.A2(n_176),
.B1(n_175),
.B2(n_171),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_253),
.B1(n_205),
.B2(n_209),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_235),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_183),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_236),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_187),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_237),
.B(n_240),
.Y(n_283)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_156),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_239),
.B(n_241),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_201),
.B(n_142),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_192),
.B(n_204),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_159),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_243),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_201),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_248),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_197),
.B(n_223),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_139),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_258),
.C(n_199),
.Y(n_263)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_188),
.A2(n_176),
.B(n_140),
.C(n_147),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_251),
.A2(n_210),
.B(n_194),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_187),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_252),
.B(n_255),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_203),
.A2(n_176),
.B1(n_169),
.B2(n_168),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_180),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_193),
.B(n_144),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_257),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_206),
.B(n_174),
.C(n_165),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_224),
.A2(n_193),
.B(n_222),
.C(n_219),
.Y(n_259)
);

OA21x2_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_220),
.B(n_211),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_207),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_260),
.B(n_236),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_250),
.A2(n_193),
.B(n_216),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_274),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_263),
.B(n_272),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_266),
.A2(n_271),
.B1(n_288),
.B2(n_251),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_267),
.B(n_235),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_216),
.B1(n_205),
.B2(n_184),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_221),
.B(n_220),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_289),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_231),
.A2(n_226),
.B(n_257),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_244),
.A2(n_225),
.B1(n_228),
.B2(n_241),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_239),
.B1(n_233),
.B2(n_234),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_244),
.Y(n_307)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_284),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_248),
.B(n_207),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_290),
.C(n_232),
.Y(n_294)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_287),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_231),
.A2(n_210),
.B1(n_194),
.B2(n_213),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_213),
.C(n_200),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_225),
.B(n_230),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_292),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_296),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_294),
.B(n_307),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_251),
.B(n_246),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_295),
.A2(n_275),
.B(n_265),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_231),
.B1(n_266),
.B2(n_276),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_297),
.A2(n_316),
.B1(n_289),
.B2(n_317),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_228),
.C(n_232),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_299),
.B(n_305),
.C(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_261),
.B(n_240),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_300),
.B(n_301),
.Y(n_328)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_303),
.B(n_314),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_261),
.B(n_242),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_304),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_259),
.C(n_258),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_263),
.B(n_259),
.C(n_260),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_264),
.B(n_255),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_309),
.B(n_292),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_265),
.B1(n_282),
.B2(n_275),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_229),
.B1(n_256),
.B2(n_254),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_311),
.A2(n_315),
.B1(n_273),
.B2(n_288),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_264),
.B(n_227),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_274),
.B1(n_283),
.B2(n_270),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_283),
.A2(n_252),
.B1(n_243),
.B2(n_237),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_321),
.A2(n_313),
.B1(n_298),
.B2(n_295),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_325),
.A2(n_342),
.B1(n_316),
.B2(n_319),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_294),
.C(n_308),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_327),
.C(n_332),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_263),
.C(n_290),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_302),
.B(n_272),
.CI(n_270),
.CON(n_329),
.SN(n_329)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_329),
.B(n_331),
.Y(n_350)
);

AO21x1_ASAP7_75t_L g359 ( 
.A1(n_330),
.A2(n_306),
.B(n_269),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_290),
.C(n_299),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_279),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_313),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_275),
.B1(n_278),
.B2(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_278),
.B1(n_291),
.B2(n_285),
.Y(n_336)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_336),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_293),
.A2(n_262),
.B1(n_284),
.B2(n_277),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g351 ( 
.A1(n_337),
.A2(n_295),
.B1(n_301),
.B2(n_312),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_272),
.C(n_282),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_279),
.C(n_298),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_306),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_313),
.A2(n_280),
.B(n_268),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_341),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_310),
.A2(n_280),
.B1(n_277),
.B2(n_269),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_345),
.B(n_357),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_332),
.B(n_302),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_346),
.B(n_349),
.C(n_360),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_347),
.A2(n_351),
.B1(n_342),
.B2(n_324),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_322),
.B(n_309),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_352),
.B(n_354),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_353),
.A2(n_321),
.B1(n_341),
.B2(n_333),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_325),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_330),
.B(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_355),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_359),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_227),
.C(n_303),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_247),
.C(n_200),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_338),
.B(n_247),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_361),
.B(n_338),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_366),
.A2(n_343),
.B1(n_371),
.B2(n_324),
.Y(n_381)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_359),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_367),
.B(n_368),
.Y(n_380)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_340),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_371),
.Y(n_382)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_347),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_372),
.B(n_374),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_348),
.B(n_320),
.C(n_326),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_373),
.B(n_360),
.C(n_327),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_339),
.Y(n_388)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_376),
.B(n_344),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_373),
.B(n_348),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_384),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_383),
.C(n_386),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_381),
.B(n_385),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_365),
.B(n_346),
.C(n_349),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_365),
.B(n_323),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_323),
.C(n_345),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_376),
.B(n_358),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_362),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_388),
.B(n_386),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_378),
.B(n_364),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_394),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_382),
.A2(n_370),
.B(n_362),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_392),
.A2(n_195),
.B(n_158),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_388),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_372),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_395),
.B(n_396),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_369),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_379),
.B(n_375),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_385),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_403),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_397),
.A2(n_368),
.B(n_363),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_404),
.B(n_405),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_363),
.C(n_367),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_358),
.C(n_334),
.Y(n_405)
);

AOI322xp5_ASAP7_75t_L g410 ( 
.A1(n_406),
.A2(n_185),
.A3(n_215),
.B1(n_161),
.B2(n_186),
.C1(n_329),
.C2(n_214),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_400),
.A2(n_391),
.B(n_396),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_408),
.A2(n_411),
.B(n_404),
.Y(n_412)
);

AO21x1_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_185),
.B(n_215),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_399),
.A2(n_390),
.B(n_329),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_SL g415 ( 
.A(n_412),
.B(n_413),
.C(n_414),
.Y(n_415)
);

AOI332xp33_ASAP7_75t_L g414 ( 
.A1(n_407),
.A2(n_405),
.A3(n_185),
.B1(n_214),
.B2(n_186),
.B3(n_155),
.C1(n_13),
.C2(n_14),
.Y(n_414)
);

AOI321xp33_ASAP7_75t_SL g416 ( 
.A1(n_415),
.A2(n_409),
.A3(n_185),
.B1(n_214),
.B2(n_186),
.C(n_13),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_416),
.B(n_12),
.Y(n_417)
);


endmodule