module fake_jpeg_7354_n_248 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_248);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_248;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_30),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_16),
.B1(n_19),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_60),
.B1(n_62),
.B2(n_24),
.Y(n_68)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_26),
.Y(n_69)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_64),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_19),
.B1(n_16),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_61),
.B1(n_32),
.B2(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_30),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_30),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_33),
.A2(n_22),
.B1(n_25),
.B2(n_23),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_33),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_32),
.C(n_20),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_40),
.C(n_17),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_74),
.B1(n_55),
.B2(n_53),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_68),
.A2(n_58),
.B1(n_55),
.B2(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_56),
.B(n_41),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_34),
.B1(n_38),
.B2(n_42),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_34),
.B1(n_26),
.B2(n_24),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_83),
.C(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_87),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_40),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_51),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_65),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_82),
.B1(n_47),
.B2(n_46),
.Y(n_134)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_90),
.B(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_91),
.A2(n_104),
.B1(n_82),
.B2(n_46),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_52),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_107),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_103),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_67),
.A2(n_55),
.B1(n_57),
.B2(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_43),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_43),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_39),
.C(n_64),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_85),
.B1(n_81),
.B2(n_84),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_135),
.B1(n_97),
.B2(n_90),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_92),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_86),
.B(n_43),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_119),
.A2(n_126),
.B(n_131),
.Y(n_152)
);

OAI32xp33_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_86),
.A3(n_78),
.B1(n_17),
.B2(n_39),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_91),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_123),
.B(n_104),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_2),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_17),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_109),
.C(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_92),
.B(n_98),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_130),
.Y(n_139)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_17),
.B(n_4),
.C(n_5),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_96),
.A2(n_31),
.B(n_5),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_47),
.B1(n_65),
.B2(n_44),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_136),
.A2(n_150),
.B(n_152),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_137),
.B(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_102),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_108),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_150),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_145),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_130),
.B1(n_131),
.B2(n_114),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_124),
.B(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_149),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_124),
.B(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_106),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_93),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_114),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_140),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_94),
.C(n_99),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_133),
.C(n_121),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_127),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_126),
.B1(n_44),
.B2(n_103),
.C(n_70),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_141),
.A2(n_115),
.B1(n_134),
.B2(n_123),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_175),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_135),
.B1(n_133),
.B2(n_122),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_146),
.A2(n_148),
.B1(n_137),
.B2(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_177),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_173),
.C(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_120),
.C(n_126),
.Y(n_173)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

OAI321xp33_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_156),
.A3(n_103),
.B1(n_70),
.B2(n_7),
.C(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_31),
.Y(n_177)
);

OAI22x1_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_103),
.B1(n_44),
.B2(n_31),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_178),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_31),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_31),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_185),
.C(n_186),
.Y(n_198)
);

AOI222xp33_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_152),
.B1(n_149),
.B2(n_143),
.C1(n_151),
.C2(n_139),
.Y(n_181)
);

AOI31xp67_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_184),
.A3(n_161),
.B(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_166),
.B(n_3),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_3),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_187)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_164),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_6),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_195),
.C(n_168),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_6),
.C(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_163),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g199 ( 
.A(n_197),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_169),
.B1(n_160),
.B2(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_194),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_208),
.C(n_195),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_165),
.C(n_170),
.Y(n_208)
);

OA21x2_ASAP7_75t_SL g209 ( 
.A1(n_181),
.A2(n_179),
.B(n_159),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_10),
.Y(n_222)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_214),
.C(n_218),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_219),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_188),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_215),
.B(n_217),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_182),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_185),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_165),
.C(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_221),
.Y(n_223)
);

OAI21x1_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_200),
.B(n_211),
.Y(n_226)
);

INVx11_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_214),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_226),
.B(n_199),
.Y(n_233)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_212),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_207),
.B1(n_206),
.B2(n_202),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_230),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_231),
.A2(n_232),
.B(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_235),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_228),
.B(n_11),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_11),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_223),
.C(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_238),
.B(n_240),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_223),
.B(n_227),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_239),
.A2(n_225),
.B(n_12),
.C(n_13),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_11),
.C(n_12),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_245),
.B(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_243),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_247),
.Y(n_248)
);


endmodule