module fake_ibex_1610_n_2563 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_417, n_471, n_265, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_465, n_48, n_325, n_57, n_301, n_434, n_296, n_120, n_168, n_155, n_315, n_441, n_13, n_122, n_116, n_370, n_431, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_22, n_136, n_261, n_459, n_30, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_52, n_448, n_99, n_466, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_420, n_483, n_141, n_222, n_186, n_349, n_454, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_429, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_480, n_416, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_447, n_26, n_188, n_200, n_444, n_199, n_410, n_308, n_463, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_479, n_225, n_360, n_272, n_23, n_468, n_223, n_381, n_382, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_482, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_460, n_476, n_461, n_313, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_344, n_393, n_436, n_428, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_424, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_425, n_2563);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_417;
input n_471;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_434;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_116;
input n_370;
input n_431;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_22;
input n_136;
input n_261;
input n_459;
input n_30;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_141;
input n_222;
input n_186;
input n_349;
input n_454;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_429;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_480;
input n_416;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_199;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_479;
input n_225;
input n_360;
input n_272;
input n_23;
input n_468;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_460;
input n_476;
input n_461;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_344;
input n_393;
input n_436;
input n_428;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_424;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;
input n_425;

output n_2563;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_622;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_1722;
wire n_911;
wire n_2023;
wire n_652;
wire n_781;
wire n_802;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_884;
wire n_667;
wire n_2396;
wire n_850;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_2475;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_2192;
wire n_1766;
wire n_550;
wire n_1922;
wire n_2032;
wire n_557;
wire n_641;
wire n_1937;
wire n_2311;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_523;
wire n_787;
wire n_2448;
wire n_614;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_538;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_2421;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_646;
wire n_2558;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_530;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_662;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_2480;
wire n_1445;
wire n_573;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_554;
wire n_553;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_2373;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_2275;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2112;
wire n_1753;
wire n_564;
wire n_562;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_592;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_2541;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2509;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_2401;
wire n_1787;
wire n_2511;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_606;
wire n_737;
wire n_2445;
wire n_1571;
wire n_1980;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_2224;
wire n_1862;
wire n_2470;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_2499;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_1591;
wire n_583;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_2101;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2456;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_1831;
wire n_608;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2390;
wire n_2423;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_2176;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_591;
wire n_1933;
wire n_2522;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_2554;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_2468;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_2549;
wire n_2461;
wire n_2006;
wire n_2440;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2441;
wire n_2358;
wire n_2490;
wire n_594;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_2062;
wire n_2277;
wire n_585;
wire n_1982;
wire n_2252;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_660;
wire n_524;
wire n_2294;
wire n_1977;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_576;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_1279;
wire n_2505;
wire n_931;
wire n_827;
wire n_607;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_488;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_2434;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_517;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2095;
wire n_555;
wire n_2486;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_502;
wire n_1705;
wire n_633;
wire n_2304;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_863;
wire n_597;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_486;
wire n_1870;
wire n_2484;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_2507;
wire n_1528;
wire n_1495;
wire n_2463;
wire n_717;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_1512;
wire n_2496;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_485;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_2459;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_588;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_2450;
wire n_528;
wire n_836;
wire n_1475;
wire n_2465;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2524;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_2545;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_510;
wire n_972;
wire n_1815;
wire n_2500;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_2442;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1349;
wire n_1331;
wire n_2127;
wire n_1323;
wire n_578;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2562;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_2446;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_598;
wire n_2141;
wire n_1422;
wire n_508;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2380;
wire n_2420;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_636;
wire n_1259;
wire n_490;
wire n_2108;
wire n_2535;
wire n_595;
wire n_1001;
wire n_570;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_487;
wire n_2528;
wire n_2548;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_625;
wire n_2113;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2320;
wire n_2268;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2447;
wire n_1057;
wire n_1473;
wire n_516;
wire n_2125;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_950;
wire n_512;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2531;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_700;
wire n_1779;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_2272;
wire n_535;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_2546;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2417;
wire n_505;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_599;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_2518;
wire n_1909;
wire n_2543;
wire n_2381;
wire n_621;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_2508;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1518;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2487;
wire n_632;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2513;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_898;
wire n_928;
wire n_1285;
wire n_967;
wire n_2561;
wire n_736;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_569;
wire n_2483;
wire n_2305;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_987;
wire n_750;
wire n_1299;
wire n_2096;
wire n_2129;
wire n_665;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_2492;
wire n_910;
wire n_2291;
wire n_635;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_704;
wire n_2357;
wire n_2148;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2302;
wire n_2560;
wire n_2092;
wire n_566;
wire n_581;
wire n_1365;
wire n_1472;
wire n_2443;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_548;
wire n_1158;
wire n_2066;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_509;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_2538;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_519;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2435;
wire n_1665;
wire n_1091;
wire n_1780;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_2282;
wire n_970;
wire n_491;
wire n_2430;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;

INVx1_ASAP7_75t_L g484 ( 
.A(n_358),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_54),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_3),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_11),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_327),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_110),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_83),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_483),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_198),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_28),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_125),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_357),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_60),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_35),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_390),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_346),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_80),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_63),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_482),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_292),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

BUFx5_ASAP7_75t_L g505 ( 
.A(n_210),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_480),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_213),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_441),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_337),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_259),
.Y(n_511)
);

NOR2xp67_ASAP7_75t_L g512 ( 
.A(n_307),
.B(n_375),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_170),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_377),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_436),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_445),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_376),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_265),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_395),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_105),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_188),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_195),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_229),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_58),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_472),
.Y(n_525)
);

NOR2xp67_ASAP7_75t_L g526 ( 
.A(n_59),
.B(n_56),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_40),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_211),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_241),
.B(n_72),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_417),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_356),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_433),
.Y(n_532)
);

CKINVDCx16_ASAP7_75t_R g533 ( 
.A(n_124),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_274),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_16),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_268),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_213),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_197),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g539 ( 
.A(n_91),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_367),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_481),
.Y(n_541)
);

NOR2xp67_ASAP7_75t_L g542 ( 
.A(n_347),
.B(n_0),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_374),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_25),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_191),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_269),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_95),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_313),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_30),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_361),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_212),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_149),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_91),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_0),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_368),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_113),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_391),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_438),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_354),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_330),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_479),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_45),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_261),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_12),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_135),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_385),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_124),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g568 ( 
.A(n_348),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_147),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_379),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_8),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_383),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_85),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_454),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_19),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_426),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_353),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_143),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_63),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_205),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_338),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_69),
.Y(n_582)
);

NOR2xp67_ASAP7_75t_L g583 ( 
.A(n_33),
.B(n_428),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_425),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_148),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_268),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_362),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_406),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_280),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_447),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_217),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_372),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_401),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_199),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_269),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_209),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_291),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_474),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_388),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_199),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_169),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_83),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_317),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_6),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_125),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_352),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_456),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_408),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_135),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_458),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_84),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_238),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_336),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_94),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_95),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_113),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_276),
.Y(n_617)
);

BUFx5_ASAP7_75t_L g618 ( 
.A(n_28),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_418),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_51),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_313),
.Y(n_621)
);

BUFx5_ASAP7_75t_L g622 ( 
.A(n_396),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_381),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_462),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_450),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_320),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_222),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_181),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_137),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_31),
.B(n_355),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_328),
.Y(n_631)
);

BUFx5_ASAP7_75t_L g632 ( 
.A(n_96),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_109),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_461),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_47),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_116),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_241),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_373),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_136),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_20),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_297),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_107),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_434),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_402),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_392),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_386),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_419),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_265),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_257),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_172),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_382),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_100),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_259),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_370),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_477),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_175),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_138),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_85),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_473),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_452),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_108),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_183),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_467),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_344),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_98),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_415),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_345),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_332),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_9),
.Y(n_669)
);

INVx1_ASAP7_75t_SL g670 ( 
.A(n_165),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_254),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_440),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_248),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_453),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_98),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_81),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_136),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_221),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_57),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_350),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_311),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_18),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_210),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_475),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_176),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_331),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_53),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_277),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_465),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_317),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_236),
.Y(n_691)
);

CKINVDCx16_ASAP7_75t_R g692 ( 
.A(n_364),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_304),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_397),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_173),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_273),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_79),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_257),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_400),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_300),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_109),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_323),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_366),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_389),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_302),
.Y(n_705)
);

INVx4_ASAP7_75t_R g706 ( 
.A(n_252),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_306),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_378),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_282),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_181),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_478),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_283),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_252),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_369),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_179),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_306),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_335),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_420),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_93),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_321),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_142),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_318),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_283),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_254),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_114),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_192),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_207),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_476),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_188),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_190),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_360),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_174),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_166),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_184),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_464),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_227),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_206),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_39),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_179),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_387),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_154),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_371),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_228),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_359),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_287),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_469),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_151),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_37),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_204),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_140),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_233),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_326),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_284),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_73),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_78),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_77),
.Y(n_756)
);

BUFx2_ASAP7_75t_L g757 ( 
.A(n_123),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_182),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_163),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_351),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_221),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_128),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_466),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_277),
.Y(n_764)
);

BUFx2_ASAP7_75t_SL g765 ( 
.A(n_66),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_86),
.Y(n_766)
);

NOR2xp67_ASAP7_75t_L g767 ( 
.A(n_94),
.B(n_140),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_250),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_444),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_411),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_300),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_449),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_203),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_12),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_76),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_304),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_303),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_87),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_116),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_380),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_468),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_168),
.Y(n_782)
);

CKINVDCx16_ASAP7_75t_R g783 ( 
.A(n_11),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_L g784 ( 
.A(n_159),
.B(n_96),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_260),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_251),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_203),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_244),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_443),
.Y(n_789)
);

INVxp67_ASAP7_75t_SL g790 ( 
.A(n_455),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_349),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_78),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_228),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_131),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_298),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_212),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_58),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_37),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_121),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_23),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_33),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_235),
.Y(n_802)
);

BUFx10_ASAP7_75t_L g803 ( 
.A(n_384),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_314),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_119),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_296),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_4),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_191),
.Y(n_808)
);

OAI22x1_ASAP7_75t_R g809 ( 
.A1(n_493),
.A2(n_649),
.B1(n_676),
.B2(n_616),
.Y(n_809)
);

XNOR2x2_ASAP7_75t_L g810 ( 
.A(n_628),
.B(n_1),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_539),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_505),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_539),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_564),
.B(n_1),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_659),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_645),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_606),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_519),
.B(n_2),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_508),
.B(n_4),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_564),
.B(n_5),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_487),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_580),
.Y(n_822)
);

BUFx12f_ASAP7_75t_L g823 ( 
.A(n_595),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_523),
.B(n_5),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_580),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_803),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_595),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_652),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_608),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_698),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_595),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_698),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_700),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_588),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_736),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_736),
.B(n_6),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_608),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_505),
.Y(n_838)
);

INVx5_ASAP7_75t_L g839 ( 
.A(n_803),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_640),
.A2(n_757),
.B1(n_568),
.B2(n_692),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_777),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_777),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_608),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_532),
.B(n_7),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_533),
.B(n_7),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_803),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_783),
.B(n_8),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_604),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_637),
.B(n_9),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_701),
.B(n_10),
.Y(n_850)
);

BUFx12f_ASAP7_75t_L g851 ( 
.A(n_741),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_669),
.B(n_10),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_608),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_644),
.Y(n_854)
);

INVx4_ASAP7_75t_L g855 ( 
.A(n_498),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_505),
.Y(n_856)
);

CKINVDCx16_ASAP7_75t_R g857 ( 
.A(n_610),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_604),
.Y(n_858)
);

OA21x2_ASAP7_75t_L g859 ( 
.A1(n_504),
.A2(n_324),
.B(n_322),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_762),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_513),
.A2(n_650),
.B1(n_665),
.B2(n_518),
.Y(n_861)
);

BUFx2_ASAP7_75t_L g862 ( 
.A(n_513),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_489),
.B(n_13),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_627),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_741),
.B(n_14),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_494),
.B(n_15),
.Y(n_866)
);

BUFx8_ASAP7_75t_SL g867 ( 
.A(n_496),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_627),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_633),
.Y(n_869)
);

CKINVDCx8_ASAP7_75t_R g870 ( 
.A(n_765),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_518),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_505),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_497),
.B(n_16),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_505),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_741),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_644),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_633),
.B(n_17),
.Y(n_877)
);

INVx4_ASAP7_75t_L g878 ( 
.A(n_499),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_650),
.A2(n_20),
.B1(n_17),
.B2(n_19),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_491),
.Y(n_880)
);

OAI22x1_ASAP7_75t_L g881 ( 
.A1(n_665),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_573),
.B(n_21),
.Y(n_882)
);

AO22x1_ASAP7_75t_L g883 ( 
.A1(n_808),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_618),
.B(n_24),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_511),
.B(n_26),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_671),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_726),
.Y(n_887)
);

AND2x6_ASAP7_75t_L g888 ( 
.A(n_731),
.B(n_325),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_726),
.B(n_26),
.Y(n_889)
);

AND2x6_ASAP7_75t_L g890 ( 
.A(n_504),
.B(n_329),
.Y(n_890)
);

INVx5_ASAP7_75t_L g891 ( 
.A(n_644),
.Y(n_891)
);

AND2x6_ASAP7_75t_L g892 ( 
.A(n_559),
.B(n_584),
.Y(n_892)
);

BUFx12f_ASAP7_75t_L g893 ( 
.A(n_806),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_730),
.B(n_27),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_730),
.B(n_27),
.Y(n_895)
);

OAI22x1_ASAP7_75t_R g896 ( 
.A1(n_496),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_520),
.B(n_29),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_644),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_734),
.Y(n_899)
);

OAI22x1_ASAP7_75t_R g900 ( 
.A1(n_527),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_502),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_734),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_537),
.B(n_32),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_549),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_559),
.A2(n_593),
.B(n_584),
.Y(n_905)
);

INVx5_ASAP7_75t_L g906 ( 
.A(n_593),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_738),
.B(n_34),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_737),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_618),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_549),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_737),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_905),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_812),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_839),
.B(n_510),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_838),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_839),
.B(n_510),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_856),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_872),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_874),
.Y(n_919)
);

CKINVDCx6p67_ASAP7_75t_R g920 ( 
.A(n_857),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_813),
.B(n_806),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_909),
.Y(n_922)
);

BUFx6f_ASAP7_75t_SL g923 ( 
.A(n_814),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_L g924 ( 
.A(n_888),
.B(n_622),
.Y(n_924)
);

AO22x2_ASAP7_75t_L g925 ( 
.A1(n_814),
.A2(n_745),
.B1(n_545),
.B2(n_548),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_877),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_839),
.B(n_668),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_817),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_813),
.B(n_808),
.Y(n_929)
);

INVxp33_ASAP7_75t_SL g930 ( 
.A(n_811),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_817),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_817),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_L g933 ( 
.A(n_815),
.B(n_799),
.C(n_797),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_817),
.Y(n_934)
);

INVx4_ASAP7_75t_L g935 ( 
.A(n_888),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_827),
.B(n_831),
.Y(n_936)
);

AO21x2_ASAP7_75t_L g937 ( 
.A1(n_863),
.A2(n_488),
.B(n_484),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_827),
.B(n_514),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_826),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_855),
.B(n_686),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_888),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_877),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_821),
.B(n_686),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_821),
.B(n_618),
.Y(n_944)
);

NOR2x1_ASAP7_75t_L g945 ( 
.A(n_846),
.B(n_495),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_884),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_889),
.Y(n_947)
);

BUFx10_ASAP7_75t_L g948 ( 
.A(n_871),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_892),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_878),
.B(n_485),
.Y(n_950)
);

OR2x2_ASAP7_75t_SL g951 ( 
.A(n_871),
.B(n_745),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_901),
.B(n_507),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_901),
.B(n_509),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_867),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_889),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_831),
.B(n_792),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_865),
.B(n_491),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_894),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_823),
.B(n_515),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_851),
.B(n_517),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_829),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_829),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_892),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_875),
.B(n_531),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_894),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_892),
.Y(n_966)
);

BUFx6f_ASAP7_75t_SL g967 ( 
.A(n_820),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_829),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_892),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_893),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_906),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_816),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_837),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_837),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_895),
.Y(n_975)
);

INVx1_ASAP7_75t_SL g976 ( 
.A(n_828),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_837),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_816),
.B(n_800),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_837),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_843),
.Y(n_980)
);

INVxp33_ASAP7_75t_L g981 ( 
.A(n_828),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_843),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_843),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_906),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_906),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_895),
.Y(n_986)
);

BUFx10_ASAP7_75t_L g987 ( 
.A(n_834),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_822),
.B(n_825),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_820),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_824),
.B(n_618),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_843),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_836),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_853),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_853),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_906),
.Y(n_995)
);

INVx1_ASAP7_75t_SL g996 ( 
.A(n_845),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_853),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_850),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_853),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_854),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_854),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_854),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_830),
.B(n_832),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_876),
.Y(n_1004)
);

OAI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_879),
.A2(n_490),
.B1(n_492),
.B2(n_486),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_SL g1006 ( 
.A(n_847),
.B(n_516),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_833),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_876),
.Y(n_1008)
);

INVx8_ASAP7_75t_L g1009 ( 
.A(n_888),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_876),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_876),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_898),
.Y(n_1012)
);

OAI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_840),
.A2(n_527),
.B1(n_616),
.B2(n_535),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_861),
.B(n_525),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_835),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_841),
.B(n_526),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_898),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_842),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_819),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_819),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_L g1021 ( 
.A(n_890),
.B(n_622),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_890),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_898),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_908),
.B(n_618),
.Y(n_1024)
);

CKINVDCx11_ASAP7_75t_R g1025 ( 
.A(n_870),
.Y(n_1025)
);

NAND2xp33_ASAP7_75t_L g1026 ( 
.A(n_890),
.B(n_622),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_908),
.B(n_500),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_849),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_898),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_849),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_867),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_818),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_880),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_848),
.B(n_529),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_859),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_910),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_904),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_911),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_818),
.B(n_530),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_858),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_904),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_844),
.B(n_543),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_904),
.Y(n_1043)
);

INVx6_ASAP7_75t_L g1044 ( 
.A(n_891),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_904),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_891),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_883),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_844),
.B(n_852),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_864),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_891),
.Y(n_1050)
);

NOR2x1p5_ASAP7_75t_L g1051 ( 
.A(n_809),
.B(n_544),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_868),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_869),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_886),
.Y(n_1054)
);

AND2x6_ASAP7_75t_L g1055 ( 
.A(n_852),
.B(n_555),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_887),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_899),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_863),
.A2(n_646),
.B(n_631),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_890),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_866),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_902),
.Y(n_1061)
);

NOR2x1p5_ASAP7_75t_L g1062 ( 
.A(n_866),
.B(n_554),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_873),
.B(n_618),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_890),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_873),
.B(n_618),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_885),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_885),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_897),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_882),
.B(n_907),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_903),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_907),
.B(n_557),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_903),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_810),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_881),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_860),
.Y(n_1075)
);

NAND2xp33_ASAP7_75t_SL g1076 ( 
.A(n_896),
.B(n_550),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_900),
.B(n_560),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_905),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_905),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_839),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_905),
.Y(n_1081)
);

AOI21x1_ASAP7_75t_L g1082 ( 
.A1(n_905),
.A2(n_646),
.B(n_631),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_862),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_813),
.B(n_501),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_812),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_905),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_877),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1053),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1053),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1054),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1067),
.A2(n_632),
.B1(n_552),
.B2(n_556),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1019),
.B(n_558),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_935),
.B(n_506),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_943),
.A2(n_590),
.B1(n_598),
.B2(n_587),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_1005),
.B(n_724),
.C(n_670),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_933),
.B(n_36),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1072),
.B(n_540),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1072),
.B(n_541),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_935),
.B(n_566),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1020),
.B(n_574),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1072),
.B(n_1028),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1030),
.B(n_1066),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_1067),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1054),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_941),
.B(n_581),
.Y(n_1105)
);

NAND2xp33_ASAP7_75t_L g1106 ( 
.A(n_1009),
.B(n_1055),
.Y(n_1106)
);

OAI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1075),
.A2(n_590),
.B1(n_599),
.B2(n_598),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1068),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_L g1109 ( 
.A(n_1013),
.B(n_759),
.C(n_751),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1070),
.B(n_1060),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_1068),
.B(n_561),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_1068),
.B(n_570),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_941),
.B(n_572),
.Y(n_1113)
);

OR2x6_ASAP7_75t_L g1114 ( 
.A(n_1051),
.B(n_767),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1048),
.B(n_592),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1060),
.B(n_576),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1063),
.B(n_577),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1057),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1063),
.B(n_624),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1057),
.Y(n_1120)
);

BUFx8_ASAP7_75t_L g1121 ( 
.A(n_970),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_950),
.B(n_625),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_956),
.B(n_634),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1065),
.B(n_626),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1024),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_924),
.B(n_521),
.C(n_503),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_946),
.B(n_789),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1065),
.B(n_651),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_943),
.B(n_654),
.Y(n_1129)
);

OAI22xp33_ASAP7_75t_SL g1130 ( 
.A1(n_1047),
.A2(n_524),
.B1(n_528),
.B2(n_522),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_938),
.B(n_1071),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_912),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_990),
.B(n_655),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_976),
.B(n_534),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1049),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_990),
.B(n_663),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_948),
.B(n_672),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_936),
.B(n_638),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_912),
.Y(n_1139)
);

AND2x6_ASAP7_75t_SL g1140 ( 
.A(n_954),
.B(n_553),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_944),
.B(n_680),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_948),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1049),
.Y(n_1143)
);

NAND2x1_ASAP7_75t_L g1144 ( 
.A(n_989),
.B(n_706),
.Y(n_1144)
);

AO221x1_ASAP7_75t_L g1145 ( 
.A1(n_970),
.A2(n_619),
.B1(n_643),
.B2(n_623),
.C(n_599),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_948),
.B(n_694),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_SL g1147 ( 
.A(n_987),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1069),
.B(n_699),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1075),
.A2(n_1074),
.B(n_926),
.C(n_1014),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_1032),
.B(n_703),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1049),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1032),
.B(n_704),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_998),
.B(n_708),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1062),
.B(n_714),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_921),
.B(n_718),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_929),
.B(n_720),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_972),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_940),
.B(n_978),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1032),
.B(n_728),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_981),
.B(n_939),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_925),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_925),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1025),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_1039),
.B(n_647),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_925),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1078),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1042),
.B(n_660),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_925),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1038),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_1025),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1055),
.B(n_742),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_992),
.B(n_744),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_992),
.B(n_769),
.Y(n_1173)
);

AND2x4_ASAP7_75t_SL g1174 ( 
.A(n_920),
.B(n_619),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_992),
.B(n_781),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1007),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1040),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1083),
.B(n_536),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_949),
.B(n_664),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_923),
.A2(n_643),
.B1(n_689),
.B2(n_623),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_987),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_SL g1182 ( 
.A(n_930),
.B(n_689),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1007),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_939),
.B(n_607),
.Y(n_1184)
);

OR2x2_ASAP7_75t_L g1185 ( 
.A(n_996),
.B(n_920),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_923),
.A2(n_770),
.B1(n_763),
.B2(n_546),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_952),
.B(n_632),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_953),
.B(n_632),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_930),
.B(n_763),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_SL g1190 ( 
.A(n_1047),
.B(n_770),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_1027),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1084),
.B(n_790),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_942),
.B(n_613),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_942),
.B(n_538),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_945),
.B(n_791),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1078),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1040),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_SL g1198 ( 
.A(n_987),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_942),
.B(n_666),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1052),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_947),
.B(n_667),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1074),
.B(n_784),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1052),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_947),
.B(n_547),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_947),
.B(n_551),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_955),
.B(n_565),
.Y(n_1206)
);

INVxp33_ASAP7_75t_L g1207 ( 
.A(n_1033),
.Y(n_1207)
);

OAI221xp5_ASAP7_75t_L g1208 ( 
.A1(n_955),
.A2(n_1087),
.B1(n_975),
.B2(n_986),
.C(n_965),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1015),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_955),
.B(n_567),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_957),
.Y(n_1211)
);

INVxp67_ASAP7_75t_L g1212 ( 
.A(n_923),
.Y(n_1212)
);

OA21x2_ASAP7_75t_L g1213 ( 
.A1(n_1079),
.A2(n_746),
.B(n_684),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1015),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_958),
.B(n_571),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_958),
.B(n_579),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_954),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_958),
.B(n_582),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_967),
.A2(n_594),
.B1(n_596),
.B2(n_591),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1018),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1018),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_951),
.A2(n_602),
.B1(n_605),
.B2(n_601),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_965),
.B(n_674),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_965),
.B(n_609),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_975),
.B(n_611),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_975),
.B(n_614),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_986),
.B(n_615),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_986),
.B(n_617),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1087),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1087),
.Y(n_1230)
);

NAND2xp33_ASAP7_75t_SL g1231 ( 
.A(n_967),
.B(n_796),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_967),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_937),
.B(n_642),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_924),
.B(n_658),
.C(n_653),
.Y(n_1234)
);

AOI221xp5_ASAP7_75t_L g1235 ( 
.A1(n_957),
.A2(n_562),
.B1(n_575),
.B2(n_569),
.C(n_563),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1056),
.Y(n_1236)
);

AO221x1_ASAP7_75t_L g1237 ( 
.A1(n_1006),
.A2(n_676),
.B1(n_722),
.B2(n_649),
.C(n_535),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_959),
.B(n_960),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_914),
.B(n_702),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_937),
.B(n_679),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1080),
.B(n_681),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1056),
.B(n_683),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1061),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_964),
.B(n_711),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_927),
.B(n_690),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_988),
.B(n_693),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_916),
.B(n_717),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1003),
.B(n_735),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1022),
.B(n_740),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1016),
.B(n_695),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1016),
.B(n_752),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1016),
.B(n_705),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1034),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1034),
.B(n_707),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_951),
.A2(n_716),
.B1(n_719),
.B2(n_712),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1034),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_915),
.B(n_723),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_971),
.Y(n_1258)
);

INVx8_ASAP7_75t_L g1259 ( 
.A(n_1064),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_971),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_984),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1085),
.B(n_725),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1085),
.B(n_727),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_985),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1058),
.B(n_729),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1058),
.B(n_732),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1077),
.B(n_733),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1022),
.B(n_760),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1081),
.B(n_1086),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_995),
.Y(n_1270)
);

INVx8_ASAP7_75t_L g1271 ( 
.A(n_1064),
.Y(n_1271)
);

INVxp67_ASAP7_75t_L g1272 ( 
.A(n_1031),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_913),
.B(n_743),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_963),
.B(n_772),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_995),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1073),
.B(n_749),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_SL g1277 ( 
.A(n_1076),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1036),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1036),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_917),
.B(n_753),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1076),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1082),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1059),
.B(n_780),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_918),
.B(n_768),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_918),
.B(n_774),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1046),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_919),
.B(n_922),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_922),
.B(n_776),
.Y(n_1288)
);

NOR3xp33_ASAP7_75t_L g1289 ( 
.A(n_1021),
.B(n_786),
.C(n_785),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1046),
.Y(n_1290)
);

NOR3xp33_ASAP7_75t_L g1291 ( 
.A(n_1021),
.B(n_788),
.C(n_586),
.Y(n_1291)
);

INVxp67_ASAP7_75t_L g1292 ( 
.A(n_1026),
.Y(n_1292)
);

OAI221xp5_ASAP7_75t_L g1293 ( 
.A1(n_1026),
.A2(n_578),
.B1(n_600),
.B2(n_597),
.C(n_589),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1059),
.B(n_1064),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1035),
.B(n_603),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1035),
.A2(n_620),
.B1(n_621),
.B2(n_612),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1035),
.A2(n_754),
.B1(n_782),
.B2(n_750),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_966),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1050),
.B(n_629),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1050),
.B(n_635),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_966),
.B(n_969),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1044),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1044),
.B(n_639),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1044),
.A2(n_648),
.B1(n_656),
.B2(n_641),
.Y(n_1304)
);

INVx2_ASAP7_75t_L g1305 ( 
.A(n_1037),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_SL g1306 ( 
.A(n_928),
.B(n_549),
.Y(n_1306)
);

INVxp67_ASAP7_75t_L g1307 ( 
.A(n_1041),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_928),
.B(n_585),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1043),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1043),
.B(n_661),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1045),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_931),
.B(n_662),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1045),
.B(n_750),
.Y(n_1313)
);

NAND2x1_ASAP7_75t_L g1314 ( 
.A(n_932),
.B(n_585),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_934),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_934),
.B(n_673),
.Y(n_1316)
);

OAI21xp33_ASAP7_75t_L g1317 ( 
.A1(n_1102),
.A2(n_677),
.B(n_675),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1103),
.B(n_678),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1142),
.B(n_1110),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1282),
.A2(n_630),
.B(n_542),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1229),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1101),
.B(n_682),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1103),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1295),
.A2(n_583),
.B(n_512),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_L g1325 ( 
.A(n_1185),
.Y(n_1325)
);

NOR3xp33_ASAP7_75t_L g1326 ( 
.A(n_1107),
.B(n_687),
.C(n_685),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1121),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1181),
.B(n_688),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1109),
.A2(n_696),
.B(n_697),
.C(n_691),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1207),
.B(n_754),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1229),
.Y(n_1331)
);

NOR2x2_ASAP7_75t_L g1332 ( 
.A(n_1182),
.B(n_782),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1178),
.Y(n_1333)
);

OAI21xp33_ASAP7_75t_L g1334 ( 
.A1(n_1134),
.A2(n_710),
.B(n_709),
.Y(n_1334)
);

INVx3_ASAP7_75t_L g1335 ( 
.A(n_1275),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1132),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1158),
.A2(n_1099),
.B(n_1294),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1238),
.B(n_787),
.Y(n_1338)
);

NAND2xp33_ASAP7_75t_L g1339 ( 
.A(n_1259),
.B(n_585),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1286),
.Y(n_1340)
);

NOR2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1163),
.B(n_787),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1295),
.A2(n_715),
.B(n_721),
.C(n_713),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1292),
.A2(n_1240),
.B(n_1233),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1191),
.B(n_739),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1189),
.B(n_794),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1161),
.A2(n_796),
.B1(n_798),
.B2(n_794),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1212),
.B(n_585),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1149),
.A2(n_748),
.B(n_755),
.C(n_747),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1135),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1230),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1191),
.B(n_756),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1092),
.B(n_758),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1092),
.B(n_761),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1121),
.Y(n_1354)
);

NOR3xp33_ASAP7_75t_L g1355 ( 
.A(n_1107),
.B(n_766),
.C(n_764),
.Y(n_1355)
);

A2O1A1Ixp33_ASAP7_75t_L g1356 ( 
.A1(n_1100),
.A2(n_773),
.B(n_775),
.C(n_771),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1176),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_SL g1358 ( 
.A(n_1147),
.B(n_798),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1265),
.A2(n_779),
.B(n_778),
.Y(n_1359)
);

INVx2_ASAP7_75t_SL g1360 ( 
.A(n_1174),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1094),
.B(n_793),
.Y(n_1361)
);

O2A1O1Ixp5_ASAP7_75t_L g1362 ( 
.A1(n_1127),
.A2(n_802),
.B(n_807),
.C(n_801),
.Y(n_1362)
);

CKINVDCx8_ASAP7_75t_R g1363 ( 
.A(n_1140),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_L g1364 ( 
.A(n_1297),
.B(n_962),
.C(n_961),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1179),
.A2(n_962),
.B(n_961),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1232),
.B(n_636),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1105),
.A2(n_973),
.B(n_968),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1232),
.B(n_657),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1160),
.B(n_657),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1289),
.B(n_795),
.C(n_657),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1231),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1183),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1105),
.A2(n_973),
.B(n_968),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1108),
.Y(n_1374)
);

A2O1A1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1115),
.A2(n_804),
.B(n_805),
.C(n_795),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1143),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1198),
.Y(n_1377)
);

A2O1A1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1115),
.A2(n_804),
.B(n_805),
.C(n_795),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1289),
.B(n_804),
.C(n_795),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1211),
.B(n_804),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1162),
.A2(n_805),
.B1(n_977),
.B2(n_974),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1151),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1109),
.A2(n_980),
.B(n_982),
.C(n_979),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1170),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1116),
.B(n_38),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_L g1386 ( 
.A(n_1130),
.B(n_991),
.C(n_983),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1301),
.A2(n_994),
.B(n_993),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1180),
.B(n_40),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1209),
.A2(n_1029),
.B(n_997),
.C(n_999),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1132),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1132),
.Y(n_1391)
);

BUFx2_ASAP7_75t_L g1392 ( 
.A(n_1313),
.Y(n_1392)
);

AOI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1274),
.A2(n_997),
.B(n_994),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1198),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1129),
.B(n_1219),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_L g1396 ( 
.A(n_1114),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1123),
.B(n_41),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1122),
.B(n_41),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1169),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_1001),
.B(n_1002),
.C(n_1000),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1122),
.B(n_1117),
.Y(n_1401)
);

AND2x6_ASAP7_75t_L g1402 ( 
.A(n_1165),
.B(n_1001),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1119),
.B(n_42),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1177),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1197),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1272),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1291),
.A2(n_1004),
.B1(n_1008),
.B2(n_1002),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1124),
.B(n_42),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1220),
.B(n_43),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_1011),
.B(n_1010),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1200),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1221),
.A2(n_1029),
.B(n_1017),
.C(n_1023),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1250),
.B(n_44),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1236),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1243),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1298),
.A2(n_1023),
.B(n_1012),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1291),
.A2(n_47),
.B1(n_44),
.B2(n_46),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1125),
.A2(n_334),
.B(n_333),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1186),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1252),
.B(n_46),
.Y(n_1420)
);

OAI21xp33_ASAP7_75t_L g1421 ( 
.A1(n_1296),
.A2(n_1148),
.B(n_1190),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_SL g1422 ( 
.A1(n_1093),
.A2(n_340),
.B(n_341),
.C(n_339),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1168),
.A2(n_50),
.B1(n_48),
.B2(n_49),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1293),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_1424)
);

AOI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1274),
.A2(n_343),
.B(n_342),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1296),
.B(n_51),
.Y(n_1426)
);

BUFx4_ASAP7_75t_SL g1427 ( 
.A(n_1217),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1299),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1091),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1254),
.B(n_52),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1203),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1137),
.B(n_55),
.Y(n_1432)
);

OAI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1091),
.A2(n_1213),
.B(n_1287),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1276),
.B(n_57),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1271),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1223),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1223),
.A2(n_64),
.B(n_61),
.C(n_62),
.Y(n_1437)
);

BUFx4f_ASAP7_75t_L g1438 ( 
.A(n_1114),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1097),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1128),
.B(n_64),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1260),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1098),
.B(n_1242),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1133),
.B(n_65),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1153),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1300),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1139),
.A2(n_1196),
.B(n_1166),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1136),
.B(n_66),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1278),
.Y(n_1448)
);

BUFx8_ASAP7_75t_L g1449 ( 
.A(n_1277),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1146),
.B(n_67),
.Y(n_1450)
);

OAI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1213),
.A2(n_365),
.B(n_363),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1279),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1126),
.A2(n_1234),
.B(n_1208),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1277),
.Y(n_1454)
);

AOI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1249),
.A2(n_1283),
.B(n_1268),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1248),
.B(n_67),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1248),
.B(n_68),
.Y(n_1457)
);

NAND3xp33_ASAP7_75t_L g1458 ( 
.A(n_1235),
.B(n_68),
.C(n_69),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1131),
.B(n_70),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1131),
.B(n_71),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1192),
.B(n_71),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1154),
.B(n_73),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1253),
.B(n_74),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1222),
.A2(n_79),
.B1(n_75),
.B2(n_77),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1256),
.B(n_80),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1144),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1303),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1194),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1255),
.A2(n_86),
.B(n_82),
.C(n_84),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1241),
.Y(n_1470)
);

O2A1O1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1127),
.A2(n_88),
.B(n_82),
.C(n_87),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1257),
.B(n_88),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1204),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1262),
.B(n_89),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_R g1475 ( 
.A(n_1281),
.B(n_1106),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1199),
.A2(n_394),
.B(n_393),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1201),
.A2(n_399),
.B(n_398),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1205),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1263),
.B(n_90),
.Y(n_1479)
);

INVx3_ASAP7_75t_SL g1480 ( 
.A(n_1114),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1304),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1258),
.A2(n_404),
.B(n_403),
.Y(n_1482)
);

OAI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1261),
.A2(n_407),
.B(n_405),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1164),
.B(n_90),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1167),
.B(n_92),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1206),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1095),
.A2(n_97),
.B(n_92),
.C(n_93),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1167),
.B(n_97),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1210),
.Y(n_1489)
);

BUFx4f_ASAP7_75t_L g1490 ( 
.A(n_1267),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1088),
.Y(n_1491)
);

AND2x2_ASAP7_75t_SL g1492 ( 
.A(n_1095),
.B(n_99),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_L g1493 ( 
.A1(n_1215),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1244),
.B(n_102),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1264),
.A2(n_410),
.B(n_409),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1187),
.A2(n_413),
.B(n_412),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1188),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1141),
.B(n_103),
.Y(n_1498)
);

O2A1O1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1216),
.A2(n_106),
.B(n_104),
.C(n_105),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1290),
.Y(n_1500)
);

OAI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1089),
.A2(n_416),
.B(n_414),
.Y(n_1501)
);

OAI321xp33_ASAP7_75t_L g1502 ( 
.A1(n_1202),
.A2(n_106),
.A3(n_107),
.B1(n_108),
.B2(n_110),
.C(n_111),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1246),
.B(n_111),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1155),
.B(n_112),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1156),
.B(n_1184),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1218),
.Y(n_1506)
);

OAI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1090),
.A2(n_422),
.B(n_421),
.Y(n_1507)
);

AOI21xp5_ASAP7_75t_L g1508 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1173),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1224),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1225),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_R g1511 ( 
.A(n_1171),
.B(n_112),
.Y(n_1511)
);

AOI21xp33_ASAP7_75t_L g1512 ( 
.A1(n_1239),
.A2(n_427),
.B(n_424),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1111),
.A2(n_430),
.B(n_429),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1237),
.B(n_114),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1112),
.A2(n_435),
.B(n_432),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1150),
.B(n_1159),
.C(n_1152),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1251),
.B(n_1193),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1157),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1251),
.B(n_115),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1271),
.Y(n_1520)
);

CKINVDCx10_ASAP7_75t_R g1521 ( 
.A(n_1202),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1104),
.Y(n_1522)
);

OAI321xp33_ASAP7_75t_L g1523 ( 
.A1(n_1202),
.A2(n_117),
.A3(n_118),
.B1(n_119),
.B2(n_120),
.C(n_121),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1118),
.B(n_117),
.Y(n_1524)
);

NOR2x1p5_ASAP7_75t_L g1525 ( 
.A(n_1145),
.B(n_118),
.Y(n_1525)
);

O2A1O1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1226),
.A2(n_123),
.B(n_120),
.C(n_122),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1227),
.B(n_122),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_1228),
.B(n_1138),
.Y(n_1528)
);

INVxp67_ASAP7_75t_L g1529 ( 
.A(n_1273),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1120),
.B(n_126),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1239),
.B(n_126),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1270),
.Y(n_1532)
);

INVx4_ASAP7_75t_L g1533 ( 
.A(n_1271),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1245),
.B(n_127),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1312),
.A2(n_439),
.B(n_437),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1312),
.A2(n_446),
.B(n_442),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1310),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1138),
.B(n_1280),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1302),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1113),
.A2(n_451),
.B(n_448),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1096),
.A2(n_1247),
.B1(n_1285),
.B2(n_1284),
.Y(n_1541)
);

NOR2xp67_ASAP7_75t_L g1542 ( 
.A(n_1195),
.B(n_129),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1288),
.B(n_130),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1316),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1309),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1307),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1307),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1547)
);

BUFx8_ASAP7_75t_L g1548 ( 
.A(n_1305),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1314),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1311),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1315),
.B(n_133),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1306),
.A2(n_138),
.B(n_134),
.C(n_137),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1308),
.A2(n_142),
.B(n_139),
.C(n_141),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1102),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1110),
.Y(n_1555)
);

INVx2_ASAP7_75t_SL g1556 ( 
.A(n_1548),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1446),
.A2(n_459),
.B(n_457),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1548),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1554),
.B(n_141),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1442),
.A2(n_463),
.B(n_460),
.Y(n_1560)
);

INVxp67_ASAP7_75t_SL g1561 ( 
.A(n_1555),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1508),
.A2(n_1337),
.B(n_1401),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1357),
.B(n_143),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1435),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1392),
.B(n_144),
.Y(n_1565)
);

AO31x2_ASAP7_75t_L g1566 ( 
.A1(n_1375),
.A2(n_144),
.A3(n_145),
.B(n_146),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1406),
.B(n_145),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1410),
.A2(n_471),
.B(n_470),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1435),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1333),
.B(n_1325),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1463),
.A2(n_1323),
.B1(n_1457),
.B2(n_1456),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1463),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1372),
.B(n_150),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1419),
.B(n_152),
.Y(n_1574)
);

NOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1354),
.B(n_153),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1325),
.B(n_153),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1427),
.Y(n_1577)
);

OR2x6_ASAP7_75t_L g1578 ( 
.A(n_1394),
.B(n_155),
.Y(n_1578)
);

OR2x6_ASAP7_75t_L g1579 ( 
.A(n_1327),
.B(n_1520),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1365),
.A2(n_156),
.B(n_157),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1414),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1415),
.Y(n_1582)
);

AOI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1383),
.A2(n_156),
.B(n_157),
.Y(n_1583)
);

INVx5_ASAP7_75t_L g1584 ( 
.A(n_1520),
.Y(n_1584)
);

AOI221x1_ASAP7_75t_L g1585 ( 
.A1(n_1324),
.A2(n_1451),
.B1(n_1320),
.B2(n_1536),
.C(n_1535),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1345),
.B(n_158),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1448),
.B(n_160),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1452),
.B(n_161),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1393),
.A2(n_162),
.B(n_163),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1433),
.A2(n_162),
.B(n_164),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1336),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1358),
.Y(n_1592)
);

NAND2x1p5_ASAP7_75t_L g1593 ( 
.A(n_1533),
.B(n_165),
.Y(n_1593)
);

OAI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1359),
.A2(n_166),
.B(n_167),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1405),
.Y(n_1595)
);

AOI21xp33_ASAP7_75t_L g1596 ( 
.A1(n_1421),
.A2(n_167),
.B(n_168),
.Y(n_1596)
);

AOI21x1_ASAP7_75t_L g1597 ( 
.A1(n_1425),
.A2(n_169),
.B(n_170),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1546),
.Y(n_1598)
);

A2O1A1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1504),
.A2(n_171),
.B(n_173),
.C(n_174),
.Y(n_1599)
);

OR2x6_ASAP7_75t_L g1600 ( 
.A(n_1377),
.B(n_319),
.Y(n_1600)
);

AO31x2_ASAP7_75t_L g1601 ( 
.A1(n_1378),
.A2(n_1348),
.A3(n_1409),
.B(n_1436),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1346),
.B(n_177),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1468),
.B(n_178),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1473),
.B(n_180),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1318),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1444),
.B(n_182),
.Y(n_1606)
);

OAI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1359),
.A2(n_183),
.B(n_184),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1478),
.B(n_185),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1486),
.B(n_185),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1449),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1481),
.A2(n_1318),
.B1(n_1426),
.B2(n_1398),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1342),
.A2(n_186),
.B(n_187),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1489),
.B(n_187),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1362),
.A2(n_189),
.B(n_190),
.Y(n_1614)
);

CKINVDCx14_ASAP7_75t_R g1615 ( 
.A(n_1384),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1501),
.A2(n_189),
.B(n_192),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1517),
.A2(n_193),
.B(n_194),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1491),
.Y(n_1618)
);

A2O1A1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1503),
.A2(n_196),
.B(n_197),
.C(n_198),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1346),
.B(n_200),
.Y(n_1620)
);

CKINVDCx20_ASAP7_75t_R g1621 ( 
.A(n_1449),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1522),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1368),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1326),
.B(n_201),
.Y(n_1624)
);

OAI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1507),
.A2(n_201),
.B(n_202),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1426),
.A2(n_205),
.B(n_206),
.Y(n_1626)
);

OAI22x1_ASAP7_75t_L g1627 ( 
.A1(n_1341),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1506),
.B(n_208),
.Y(n_1628)
);

BUFx2_ASAP7_75t_SL g1629 ( 
.A(n_1377),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1399),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1404),
.Y(n_1631)
);

O2A1O1Ixp5_ASAP7_75t_L g1632 ( 
.A1(n_1324),
.A2(n_214),
.B(n_215),
.C(n_216),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1330),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1509),
.B(n_219),
.Y(n_1634)
);

INVx8_ASAP7_75t_L g1635 ( 
.A(n_1368),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1510),
.B(n_223),
.Y(n_1636)
);

OAI22x1_ASAP7_75t_L g1637 ( 
.A1(n_1525),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_1637)
);

OAI22x1_ASAP7_75t_L g1638 ( 
.A1(n_1371),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_1638)
);

INVx1_ASAP7_75t_SL g1639 ( 
.A(n_1328),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1537),
.A2(n_230),
.B(n_231),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1428),
.B(n_232),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1397),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1483),
.A2(n_1495),
.B(n_1387),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1445),
.B(n_234),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1411),
.A2(n_237),
.B(n_238),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_SL g1646 ( 
.A1(n_1492),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1355),
.B(n_239),
.Y(n_1647)
);

OA22x2_ASAP7_75t_L g1648 ( 
.A1(n_1388),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1395),
.B(n_245),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_1328),
.Y(n_1650)
);

A2O1A1Ixp33_ASAP7_75t_L g1651 ( 
.A1(n_1527),
.A2(n_246),
.B(n_247),
.C(n_249),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1524),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1431),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1441),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1335),
.Y(n_1655)
);

OAI22x1_ASAP7_75t_L g1656 ( 
.A1(n_1464),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_1656)
);

AND2x6_ASAP7_75t_L g1657 ( 
.A(n_1335),
.B(n_253),
.Y(n_1657)
);

INVx4_ASAP7_75t_L g1658 ( 
.A(n_1340),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1338),
.B(n_253),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1439),
.B(n_255),
.Y(n_1660)
);

OAI21xp33_ASAP7_75t_L g1661 ( 
.A1(n_1334),
.A2(n_255),
.B(n_256),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1467),
.B(n_258),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_L g1663 ( 
.A1(n_1344),
.A2(n_262),
.B(n_263),
.Y(n_1663)
);

INVx5_ASAP7_75t_L g1664 ( 
.A(n_1402),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1521),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1547),
.A2(n_264),
.B(n_266),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1516),
.B(n_264),
.Y(n_1667)
);

NAND3xp33_ASAP7_75t_SL g1668 ( 
.A(n_1363),
.B(n_266),
.C(n_267),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1511),
.B(n_270),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1519),
.A2(n_270),
.B(n_271),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1505),
.A2(n_1543),
.B(n_1420),
.C(n_1430),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1390),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1403),
.A2(n_271),
.B(n_272),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1370),
.A2(n_272),
.B(n_273),
.Y(n_1674)
);

INVx2_ASAP7_75t_SL g1675 ( 
.A(n_1360),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1413),
.A2(n_274),
.B(n_275),
.C(n_276),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1530),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1408),
.A2(n_275),
.B(n_278),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_SL g1679 ( 
.A(n_1319),
.B(n_279),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1440),
.A2(n_281),
.B(n_282),
.Y(n_1680)
);

OR2x6_ASAP7_75t_L g1681 ( 
.A(n_1545),
.B(n_319),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1396),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1322),
.Y(n_1683)
);

AOI221x1_ASAP7_75t_L g1684 ( 
.A1(n_1535),
.A2(n_285),
.B1(n_286),
.B2(n_288),
.C(n_289),
.Y(n_1684)
);

BUFx3_ASAP7_75t_L g1685 ( 
.A(n_1396),
.Y(n_1685)
);

BUFx10_ASAP7_75t_L g1686 ( 
.A(n_1432),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1350),
.B(n_285),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1454),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1529),
.B(n_289),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1356),
.B(n_290),
.Y(n_1690)
);

INVx5_ASAP7_75t_L g1691 ( 
.A(n_1402),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1438),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1443),
.A2(n_1447),
.B(n_1416),
.Y(n_1693)
);

OAI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1379),
.A2(n_292),
.B(n_293),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1352),
.B(n_293),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1353),
.B(n_294),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1470),
.B(n_294),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_SL g1698 ( 
.A1(n_1496),
.A2(n_295),
.B(n_296),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1490),
.B(n_299),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1351),
.B(n_301),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1461),
.Y(n_1701)
);

BUFx4f_ASAP7_75t_L g1702 ( 
.A(n_1480),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1434),
.B(n_1317),
.Y(n_1703)
);

AO31x2_ASAP7_75t_L g1704 ( 
.A1(n_1437),
.A2(n_303),
.A3(n_305),
.B(n_307),
.Y(n_1704)
);

AOI211x1_ASAP7_75t_L g1705 ( 
.A1(n_1458),
.A2(n_305),
.B(n_308),
.C(n_309),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1459),
.B(n_308),
.Y(n_1706)
);

AOI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1493),
.A2(n_310),
.B(n_311),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1498),
.A2(n_312),
.B(n_314),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1329),
.A2(n_312),
.B1(n_315),
.B2(n_316),
.C(n_318),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1453),
.A2(n_315),
.B(n_316),
.Y(n_1710)
);

OAI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1453),
.A2(n_1531),
.B(n_1460),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1361),
.B(n_1490),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1531),
.B(n_1364),
.Y(n_1713)
);

INVx2_ASAP7_75t_SL g1714 ( 
.A(n_1438),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1462),
.B(n_1465),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1340),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1547),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1500),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1514),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1472),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1475),
.B(n_1484),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1389),
.A2(n_1412),
.B(n_1400),
.Y(n_1722)
);

AO31x2_ASAP7_75t_L g1723 ( 
.A1(n_1381),
.A2(n_1544),
.A3(n_1429),
.B(n_1497),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1466),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1532),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1494),
.B(n_1450),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1518),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1391),
.Y(n_1728)
);

OAI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1485),
.A2(n_1488),
.B(n_1385),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1367),
.A2(n_1373),
.B(n_1513),
.Y(n_1730)
);

AO21x1_ASAP7_75t_L g1731 ( 
.A1(n_1512),
.A2(n_1429),
.B(n_1499),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_L g1732 ( 
.A1(n_1515),
.A2(n_1540),
.B(n_1476),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1518),
.Y(n_1733)
);

NOR4xp25_ASAP7_75t_L g1734 ( 
.A(n_1487),
.B(n_1469),
.C(n_1502),
.D(n_1523),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1374),
.Y(n_1735)
);

AOI21xp33_ASAP7_75t_L g1736 ( 
.A1(n_1526),
.A2(n_1424),
.B(n_1471),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1474),
.B(n_1479),
.Y(n_1737)
);

INVx6_ASAP7_75t_SL g1738 ( 
.A(n_1386),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1417),
.B(n_1423),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_SL g1740 ( 
.A1(n_1339),
.A2(n_1534),
.B(n_1551),
.Y(n_1740)
);

OAI21x1_ASAP7_75t_L g1741 ( 
.A1(n_1477),
.A2(n_1349),
.B(n_1376),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1321),
.B(n_1331),
.Y(n_1742)
);

BUFx12f_ASAP7_75t_L g1743 ( 
.A(n_1549),
.Y(n_1743)
);

OAI21x1_ASAP7_75t_L g1744 ( 
.A1(n_1349),
.A2(n_1382),
.B(n_1376),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1380),
.A2(n_1369),
.B(n_1552),
.C(n_1553),
.Y(n_1745)
);

OAI22x1_ASAP7_75t_L g1746 ( 
.A1(n_1347),
.A2(n_1366),
.B1(n_1542),
.B2(n_1382),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1402),
.A2(n_1539),
.B1(n_1550),
.B2(n_1407),
.Y(n_1747)
);

AO31x2_ASAP7_75t_L g1748 ( 
.A1(n_1422),
.A2(n_1375),
.A3(n_1378),
.B(n_1348),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1455),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1750)
);

OAI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_SL g1754 ( 
.A(n_1358),
.B(n_1182),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_1336),
.Y(n_1755)
);

INVx6_ASAP7_75t_L g1756 ( 
.A(n_1548),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1554),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1548),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1554),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1538),
.A2(n_1528),
.B(n_1401),
.C(n_1442),
.Y(n_1761)
);

O2A1O1Ixp5_ASAP7_75t_L g1762 ( 
.A1(n_1541),
.A2(n_1324),
.B(n_1320),
.C(n_1534),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1763)
);

OAI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1435),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1330),
.A2(n_1107),
.B1(n_1189),
.B2(n_1182),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1554),
.B(n_1142),
.Y(n_1770)
);

BUFx12f_ASAP7_75t_L g1771 ( 
.A(n_1327),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1554),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1336),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1442),
.A2(n_924),
.B(n_1269),
.Y(n_1776)
);

CKINVDCx11_ASAP7_75t_R g1777 ( 
.A(n_1363),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1555),
.B(n_1060),
.Y(n_1778)
);

A2O1A1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1538),
.A2(n_1528),
.B(n_1401),
.C(n_1442),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1554),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1555),
.Y(n_1782)
);

AO31x2_ASAP7_75t_L g1783 ( 
.A1(n_1375),
.A2(n_1378),
.A3(n_1348),
.B(n_1295),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1785)
);

AOI221xp5_ASAP7_75t_L g1786 ( 
.A1(n_1329),
.A2(n_1554),
.B1(n_1326),
.B2(n_1355),
.C(n_1356),
.Y(n_1786)
);

BUFx3_ASAP7_75t_L g1787 ( 
.A(n_1548),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1555),
.B(n_1060),
.Y(n_1788)
);

OA22x2_ASAP7_75t_L g1789 ( 
.A1(n_1346),
.A2(n_1297),
.B1(n_1237),
.B2(n_1180),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1555),
.B(n_1060),
.Y(n_1790)
);

A2O1A1Ixp33_ASAP7_75t_L g1791 ( 
.A1(n_1538),
.A2(n_1528),
.B(n_1401),
.C(n_1442),
.Y(n_1791)
);

INVx3_ASAP7_75t_L g1792 ( 
.A(n_1435),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_SL g1795 ( 
.A(n_1554),
.B(n_1142),
.Y(n_1795)
);

AND2x2_ASAP7_75t_SL g1796 ( 
.A(n_1358),
.B(n_1174),
.Y(n_1796)
);

BUFx2_ASAP7_75t_L g1797 ( 
.A(n_1548),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1554),
.Y(n_1798)
);

INVx6_ASAP7_75t_L g1799 ( 
.A(n_1548),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1800)
);

O2A1O1Ixp5_ASAP7_75t_L g1801 ( 
.A1(n_1541),
.A2(n_1324),
.B(n_1320),
.C(n_1534),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1554),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1508),
.A2(n_1442),
.B(n_1401),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_SL g1806 ( 
.A1(n_1418),
.A2(n_1483),
.B(n_1482),
.Y(n_1806)
);

INVx4_ASAP7_75t_L g1807 ( 
.A(n_1354),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1419),
.B(n_1182),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1810)
);

AOI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1330),
.A2(n_1107),
.B1(n_1189),
.B2(n_1182),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1555),
.B(n_1060),
.Y(n_1813)
);

INVx3_ASAP7_75t_L g1814 ( 
.A(n_1435),
.Y(n_1814)
);

AOI221x1_ASAP7_75t_L g1815 ( 
.A1(n_1324),
.A2(n_1451),
.B1(n_1320),
.B2(n_1536),
.C(n_1535),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_SL g1817 ( 
.A(n_1554),
.B(n_1142),
.Y(n_1817)
);

BUFx8_ASAP7_75t_L g1818 ( 
.A(n_1327),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1554),
.B(n_1102),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1554),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1343),
.A2(n_1433),
.B(n_1337),
.Y(n_1822)
);

AOI21xp33_ASAP7_75t_L g1823 ( 
.A1(n_1611),
.A2(n_1715),
.B(n_1713),
.Y(n_1823)
);

BUFx8_ASAP7_75t_L g1824 ( 
.A(n_1797),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1584),
.B(n_1556),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1756),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1752),
.B(n_1768),
.Y(n_1827)
);

BUFx2_ASAP7_75t_L g1828 ( 
.A(n_1558),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1584),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1787),
.Y(n_1830)
);

BUFx2_ASAP7_75t_SL g1831 ( 
.A(n_1610),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1782),
.B(n_1778),
.Y(n_1832)
);

BUFx10_ASAP7_75t_L g1833 ( 
.A(n_1756),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1561),
.Y(n_1834)
);

INVx4_ASAP7_75t_L g1835 ( 
.A(n_1584),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1769),
.B(n_1775),
.Y(n_1836)
);

AO21x1_ASAP7_75t_L g1837 ( 
.A1(n_1710),
.A2(n_1590),
.B(n_1611),
.Y(n_1837)
);

NAND2x1p5_ASAP7_75t_L g1838 ( 
.A(n_1584),
.B(n_1664),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1751),
.A2(n_1785),
.B(n_1764),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1767),
.B(n_1811),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1769),
.B(n_1775),
.Y(n_1841)
);

BUFx4f_ASAP7_75t_L g1842 ( 
.A(n_1756),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1780),
.B(n_1784),
.Y(n_1843)
);

OA21x2_ASAP7_75t_L g1844 ( 
.A1(n_1585),
.A2(n_1815),
.B(n_1804),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1761),
.A2(n_1791),
.B(n_1779),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1793),
.Y(n_1846)
);

NOR2xp67_ASAP7_75t_L g1847 ( 
.A(n_1759),
.B(n_1807),
.Y(n_1847)
);

OA21x2_ASAP7_75t_L g1848 ( 
.A1(n_1803),
.A2(n_1822),
.B(n_1810),
.Y(n_1848)
);

AO21x2_ASAP7_75t_L g1849 ( 
.A1(n_1804),
.A2(n_1810),
.B(n_1822),
.Y(n_1849)
);

OAI21x1_ASAP7_75t_L g1850 ( 
.A1(n_1730),
.A2(n_1562),
.B(n_1732),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_1577),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1794),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1788),
.B(n_1790),
.Y(n_1853)
);

BUFx12f_ASAP7_75t_L g1854 ( 
.A(n_1777),
.Y(n_1854)
);

BUFx4_ASAP7_75t_SL g1855 ( 
.A(n_1621),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1799),
.Y(n_1856)
);

OAI21x1_ASAP7_75t_SL g1857 ( 
.A1(n_1698),
.A2(n_1571),
.B(n_1594),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1800),
.Y(n_1858)
);

CKINVDCx20_ASAP7_75t_R g1859 ( 
.A(n_1818),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1813),
.B(n_1800),
.Y(n_1860)
);

OAI21x1_ASAP7_75t_L g1861 ( 
.A1(n_1693),
.A2(n_1597),
.B(n_1722),
.Y(n_1861)
);

NOR2x1_ASAP7_75t_R g1862 ( 
.A(n_1799),
.B(n_1665),
.Y(n_1862)
);

NAND2x1p5_ASAP7_75t_L g1863 ( 
.A(n_1664),
.B(n_1691),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1722),
.A2(n_1741),
.B(n_1557),
.Y(n_1864)
);

INVx3_ASAP7_75t_SL g1865 ( 
.A(n_1799),
.Y(n_1865)
);

AO21x2_ASAP7_75t_L g1866 ( 
.A1(n_1711),
.A2(n_1596),
.B(n_1729),
.Y(n_1866)
);

AO21x2_ASAP7_75t_L g1867 ( 
.A1(n_1711),
.A2(n_1596),
.B(n_1729),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1564),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1717),
.A2(n_1789),
.B1(n_1739),
.B2(n_1786),
.Y(n_1869)
);

INVx5_ASAP7_75t_L g1870 ( 
.A(n_1657),
.Y(n_1870)
);

OAI21x1_ASAP7_75t_L g1871 ( 
.A1(n_1744),
.A2(n_1589),
.B(n_1580),
.Y(n_1871)
);

CKINVDCx20_ASAP7_75t_R g1872 ( 
.A(n_1818),
.Y(n_1872)
);

OAI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1568),
.A2(n_1625),
.B(n_1616),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1564),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1569),
.Y(n_1875)
);

INVx4_ASAP7_75t_L g1876 ( 
.A(n_1807),
.Y(n_1876)
);

AOI22x1_ASAP7_75t_L g1877 ( 
.A1(n_1746),
.A2(n_1805),
.B1(n_1637),
.B2(n_1560),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1809),
.B(n_1812),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1569),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1816),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1816),
.B(n_1819),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1819),
.B(n_1820),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1766),
.Y(n_1883)
);

OA21x2_ASAP7_75t_L g1884 ( 
.A1(n_1684),
.A2(n_1801),
.B(n_1762),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1808),
.B(n_1820),
.Y(n_1885)
);

INVx4_ASAP7_75t_L g1886 ( 
.A(n_1579),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_SL g1887 ( 
.A(n_1754),
.B(n_1646),
.C(n_1666),
.Y(n_1887)
);

CKINVDCx6p67_ASAP7_75t_R g1888 ( 
.A(n_1771),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_SL g1889 ( 
.A(n_1796),
.B(n_1702),
.Y(n_1889)
);

BUFx3_ASAP7_75t_L g1890 ( 
.A(n_1766),
.Y(n_1890)
);

BUFx3_ASAP7_75t_L g1891 ( 
.A(n_1792),
.Y(n_1891)
);

OR2x6_ASAP7_75t_L g1892 ( 
.A(n_1629),
.B(n_1579),
.Y(n_1892)
);

OAI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1805),
.A2(n_1671),
.B(n_1750),
.Y(n_1893)
);

NOR2xp67_ASAP7_75t_L g1894 ( 
.A(n_1682),
.B(n_1714),
.Y(n_1894)
);

AO21x2_ASAP7_75t_L g1895 ( 
.A1(n_1731),
.A2(n_1583),
.B(n_1736),
.Y(n_1895)
);

BUFx8_ASAP7_75t_SL g1896 ( 
.A(n_1702),
.Y(n_1896)
);

NAND3xp33_ASAP7_75t_L g1897 ( 
.A(n_1705),
.B(n_1632),
.C(n_1651),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1792),
.Y(n_1898)
);

BUFx6f_ASAP7_75t_L g1899 ( 
.A(n_1591),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1579),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1753),
.A2(n_1763),
.B(n_1757),
.Y(n_1901)
);

AO31x2_ASAP7_75t_L g1902 ( 
.A1(n_1713),
.A2(n_1571),
.A3(n_1677),
.B(n_1652),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1786),
.B(n_1683),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1758),
.B(n_1760),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1781),
.B(n_1798),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1765),
.A2(n_1776),
.B(n_1773),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_1814),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1814),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1605),
.B(n_1772),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1802),
.Y(n_1910)
);

BUFx2_ASAP7_75t_R g1911 ( 
.A(n_1688),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1712),
.B(n_1719),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1821),
.B(n_1570),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1743),
.Y(n_1914)
);

AO21x2_ASAP7_75t_L g1915 ( 
.A1(n_1583),
.A2(n_1736),
.B(n_1707),
.Y(n_1915)
);

BUFx2_ASAP7_75t_L g1916 ( 
.A(n_1615),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_L g1917 ( 
.A(n_1599),
.B(n_1619),
.C(n_1676),
.Y(n_1917)
);

OA21x2_ASAP7_75t_L g1918 ( 
.A1(n_1674),
.A2(n_1694),
.B(n_1626),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1635),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1581),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1598),
.B(n_1697),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1718),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1559),
.Y(n_1923)
);

BUFx4f_ASAP7_75t_L g1924 ( 
.A(n_1578),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1726),
.B(n_1582),
.Y(n_1925)
);

A2O1A1Ixp33_ASAP7_75t_L g1926 ( 
.A1(n_1594),
.A2(n_1607),
.B(n_1612),
.C(n_1617),
.Y(n_1926)
);

INVx2_ASAP7_75t_SL g1927 ( 
.A(n_1685),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_SL g1928 ( 
.A1(n_1607),
.A2(n_1640),
.B(n_1645),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1635),
.Y(n_1929)
);

AND2x4_ASAP7_75t_L g1930 ( 
.A(n_1595),
.B(n_1664),
.Y(n_1930)
);

OA21x2_ASAP7_75t_L g1931 ( 
.A1(n_1626),
.A2(n_1640),
.B(n_1645),
.Y(n_1931)
);

BUFx2_ASAP7_75t_R g1932 ( 
.A(n_1692),
.Y(n_1932)
);

BUFx2_ASAP7_75t_SL g1933 ( 
.A(n_1657),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1691),
.B(n_1701),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1691),
.B(n_1720),
.Y(n_1935)
);

INVx1_ASAP7_75t_SL g1936 ( 
.A(n_1639),
.Y(n_1936)
);

INVx4_ASAP7_75t_L g1937 ( 
.A(n_1600),
.Y(n_1937)
);

OAI21x1_ASAP7_75t_L g1938 ( 
.A1(n_1747),
.A2(n_1706),
.B(n_1740),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_SL g1939 ( 
.A1(n_1679),
.A2(n_1612),
.B(n_1572),
.Y(n_1939)
);

BUFx2_ASAP7_75t_L g1940 ( 
.A(n_1578),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1700),
.B(n_1618),
.Y(n_1941)
);

OAI21x1_ASAP7_75t_SL g1942 ( 
.A1(n_1572),
.A2(n_1614),
.B(n_1641),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1789),
.A2(n_1667),
.B1(n_1648),
.B2(n_1620),
.Y(n_1943)
);

BUFx2_ASAP7_75t_SL g1944 ( 
.A(n_1657),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1658),
.Y(n_1945)
);

NAND3xp33_ASAP7_75t_L g1946 ( 
.A(n_1709),
.B(n_1633),
.C(n_1670),
.Y(n_1946)
);

AO21x2_ASAP7_75t_L g1947 ( 
.A1(n_1737),
.A2(n_1614),
.B(n_1734),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1660),
.B(n_1650),
.Y(n_1948)
);

AOI22xp33_ASAP7_75t_L g1949 ( 
.A1(n_1648),
.A2(n_1602),
.B1(n_1574),
.B2(n_1647),
.Y(n_1949)
);

BUFx12f_ASAP7_75t_L g1950 ( 
.A(n_1578),
.Y(n_1950)
);

AO21x2_ASAP7_75t_L g1951 ( 
.A1(n_1649),
.A2(n_1703),
.B(n_1745),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1644),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1727),
.B(n_1655),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1709),
.A2(n_1661),
.B(n_1649),
.C(n_1663),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1622),
.B(n_1659),
.Y(n_1955)
);

OAI21xp5_ASAP7_75t_L g1956 ( 
.A1(n_1603),
.A2(n_1628),
.B(n_1636),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1559),
.B(n_1634),
.Y(n_1957)
);

OAI21x1_ASAP7_75t_L g1958 ( 
.A1(n_1563),
.A2(n_1587),
.B(n_1573),
.Y(n_1958)
);

OAI21x1_ASAP7_75t_L g1959 ( 
.A1(n_1742),
.A2(n_1687),
.B(n_1588),
.Y(n_1959)
);

NAND2x1p5_ASAP7_75t_L g1960 ( 
.A(n_1634),
.B(n_1658),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1644),
.Y(n_1961)
);

OAI21x1_ASAP7_75t_L g1962 ( 
.A1(n_1742),
.A2(n_1687),
.B(n_1587),
.Y(n_1962)
);

O2A1O1Ixp33_ASAP7_75t_L g1963 ( 
.A1(n_1690),
.A2(n_1608),
.B(n_1628),
.C(n_1613),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1603),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1604),
.Y(n_1965)
);

OAI21x1_ASAP7_75t_L g1966 ( 
.A1(n_1662),
.A2(n_1721),
.B(n_1673),
.Y(n_1966)
);

AO21x2_ASAP7_75t_L g1967 ( 
.A1(n_1695),
.A2(n_1696),
.B(n_1662),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1604),
.A2(n_1613),
.B(n_1609),
.Y(n_1968)
);

CKINVDCx16_ASAP7_75t_R g1969 ( 
.A(n_1600),
.Y(n_1969)
);

OA21x2_ASAP7_75t_L g1970 ( 
.A1(n_1678),
.A2(n_1680),
.B(n_1708),
.Y(n_1970)
);

OAI21x1_ASAP7_75t_L g1971 ( 
.A1(n_1608),
.A2(n_1609),
.B(n_1593),
.Y(n_1971)
);

OA21x2_ASAP7_75t_L g1972 ( 
.A1(n_1690),
.A2(n_1735),
.B(n_1642),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_L g1973 ( 
.A(n_1592),
.B(n_1675),
.Y(n_1973)
);

OA21x2_ASAP7_75t_L g1974 ( 
.A1(n_1642),
.A2(n_1654),
.B(n_1653),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1689),
.A2(n_1817),
.B(n_1795),
.Y(n_1975)
);

INVx1_ASAP7_75t_SL g1976 ( 
.A(n_1576),
.Y(n_1976)
);

BUFx2_ASAP7_75t_R g1977 ( 
.A(n_1724),
.Y(n_1977)
);

AOI21xp33_ASAP7_75t_L g1978 ( 
.A1(n_1623),
.A2(n_1635),
.B(n_1770),
.Y(n_1978)
);

OAI21x1_ASAP7_75t_L g1979 ( 
.A1(n_1630),
.A2(n_1725),
.B(n_1631),
.Y(n_1979)
);

NOR2x1_ASAP7_75t_L g1980 ( 
.A(n_1600),
.B(n_1681),
.Y(n_1980)
);

NAND3xp33_ASAP7_75t_L g1981 ( 
.A(n_1699),
.B(n_1575),
.C(n_1669),
.Y(n_1981)
);

AO21x2_ASAP7_75t_L g1982 ( 
.A1(n_1586),
.A2(n_1624),
.B(n_1749),
.Y(n_1982)
);

OA21x2_ASAP7_75t_L g1983 ( 
.A1(n_1749),
.A2(n_1606),
.B(n_1704),
.Y(n_1983)
);

INVx5_ASAP7_75t_L g1984 ( 
.A(n_1657),
.Y(n_1984)
);

BUFx12f_ASAP7_75t_L g1985 ( 
.A(n_1681),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1565),
.B(n_1567),
.Y(n_1986)
);

BUFx2_ASAP7_75t_L g1987 ( 
.A(n_1681),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1686),
.B(n_1733),
.Y(n_1988)
);

INVx2_ASAP7_75t_SL g1989 ( 
.A(n_1716),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1656),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1672),
.A2(n_1728),
.B(n_1774),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1704),
.Y(n_1992)
);

INVx2_ASAP7_75t_SL g1993 ( 
.A(n_1627),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1755),
.B(n_1601),
.Y(n_1994)
);

INVx3_ASAP7_75t_SL g1995 ( 
.A(n_1755),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1738),
.A2(n_1748),
.B(n_1601),
.Y(n_1996)
);

AO21x2_ASAP7_75t_L g1997 ( 
.A1(n_1601),
.A2(n_1748),
.B(n_1783),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1668),
.B(n_1723),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1638),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1566),
.Y(n_2000)
);

INVx4_ASAP7_75t_L g2001 ( 
.A(n_1566),
.Y(n_2001)
);

AND2x4_ASAP7_75t_L g2002 ( 
.A(n_1783),
.B(n_1748),
.Y(n_2002)
);

A2O1A1Ixp33_ASAP7_75t_L g2003 ( 
.A1(n_1805),
.A2(n_1779),
.B(n_1791),
.C(n_1761),
.Y(n_2003)
);

CKINVDCx20_ASAP7_75t_R g2004 ( 
.A(n_1610),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1571),
.A2(n_1717),
.B1(n_1779),
.B2(n_1761),
.Y(n_2005)
);

NOR2x1_ASAP7_75t_SL g2006 ( 
.A(n_1584),
.B(n_1664),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1778),
.B(n_1788),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1752),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1611),
.B(n_1571),
.Y(n_2009)
);

BUFx2_ASAP7_75t_R g2010 ( 
.A(n_1577),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1752),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1752),
.Y(n_2012)
);

INVx3_ASAP7_75t_L g2013 ( 
.A(n_1584),
.Y(n_2013)
);

OA21x2_ASAP7_75t_L g2014 ( 
.A1(n_1585),
.A2(n_1815),
.B(n_1643),
.Y(n_2014)
);

OR3x4_ASAP7_75t_SL g2015 ( 
.A(n_1561),
.B(n_1332),
.C(n_1363),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_1577),
.Y(n_2016)
);

AO21x2_ASAP7_75t_L g2017 ( 
.A1(n_1806),
.A2(n_1764),
.B(n_1751),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_L g2018 ( 
.A(n_1767),
.B(n_1419),
.Y(n_2018)
);

INVx2_ASAP7_75t_SL g2019 ( 
.A(n_1756),
.Y(n_2019)
);

INVx3_ASAP7_75t_L g2020 ( 
.A(n_1584),
.Y(n_2020)
);

OA21x2_ASAP7_75t_L g2021 ( 
.A1(n_1585),
.A2(n_1815),
.B(n_1643),
.Y(n_2021)
);

INVxp67_ASAP7_75t_L g2022 ( 
.A(n_1752),
.Y(n_2022)
);

BUFx4f_ASAP7_75t_L g2023 ( 
.A(n_1756),
.Y(n_2023)
);

BUFx2_ASAP7_75t_L g2024 ( 
.A(n_1797),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1752),
.B(n_1768),
.Y(n_2025)
);

INVxp67_ASAP7_75t_SL g2026 ( 
.A(n_1752),
.Y(n_2026)
);

NAND2x1p5_ASAP7_75t_L g2027 ( 
.A(n_1584),
.B(n_1435),
.Y(n_2027)
);

AO21x1_ASAP7_75t_L g2028 ( 
.A1(n_1710),
.A2(n_1590),
.B(n_1611),
.Y(n_2028)
);

INVx3_ASAP7_75t_SL g2029 ( 
.A(n_1756),
.Y(n_2029)
);

AO21x2_ASAP7_75t_L g2030 ( 
.A1(n_1806),
.A2(n_1764),
.B(n_1751),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1846),
.Y(n_2031)
);

CKINVDCx5p33_ASAP7_75t_R g2032 ( 
.A(n_1855),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1904),
.Y(n_2033)
);

CKINVDCx20_ASAP7_75t_R g2034 ( 
.A(n_2004),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1905),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2026),
.B(n_1846),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1836),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1881),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1843),
.B(n_1878),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_2005),
.A2(n_1869),
.B1(n_2018),
.B2(n_1840),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1843),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1878),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1923),
.Y(n_2043)
);

BUFx3_ASAP7_75t_L g2044 ( 
.A(n_2027),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1882),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2025),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2025),
.B(n_1853),
.Y(n_2047)
);

CKINVDCx20_ASAP7_75t_R g2048 ( 
.A(n_2004),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_2025),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1869),
.A2(n_2018),
.B1(n_1840),
.B2(n_1887),
.Y(n_2050)
);

BUFx2_ASAP7_75t_R g2051 ( 
.A(n_1896),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_1824),
.Y(n_2052)
);

BUFx3_ASAP7_75t_L g2053 ( 
.A(n_2027),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1827),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2007),
.B(n_2022),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1841),
.Y(n_2056)
);

CKINVDCx5p33_ASAP7_75t_R g2057 ( 
.A(n_1855),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1923),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1885),
.A2(n_1845),
.B1(n_1943),
.B2(n_2009),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_SL g2060 ( 
.A1(n_1924),
.A2(n_1985),
.B1(n_1969),
.B2(n_1937),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1852),
.B(n_1858),
.Y(n_2061)
);

BUFx12f_ASAP7_75t_L g2062 ( 
.A(n_1854),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1858),
.B(n_1880),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1859),
.Y(n_2064)
);

OAI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_1926),
.A2(n_1954),
.B(n_2003),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1885),
.A2(n_1943),
.B1(n_1924),
.B2(n_1823),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_1829),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2022),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1880),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2003),
.B(n_1903),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1860),
.Y(n_2071)
);

BUFx3_ASAP7_75t_L g2072 ( 
.A(n_1829),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1835),
.Y(n_2073)
);

BUFx3_ASAP7_75t_L g2074 ( 
.A(n_1919),
.Y(n_2074)
);

NAND2x1p5_ASAP7_75t_L g2075 ( 
.A(n_1870),
.B(n_1984),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1832),
.B(n_1834),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1920),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1892),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_1824),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1910),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1902),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2008),
.Y(n_2082)
);

BUFx8_ASAP7_75t_L g2083 ( 
.A(n_1854),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1824),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1913),
.B(n_2011),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_1916),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_1919),
.Y(n_2087)
);

NAND2x1p5_ASAP7_75t_L g2088 ( 
.A(n_1870),
.B(n_1984),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_2012),
.B(n_1976),
.Y(n_2089)
);

INVxp67_ASAP7_75t_SL g2090 ( 
.A(n_1960),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1835),
.Y(n_2091)
);

INVx3_ASAP7_75t_L g2092 ( 
.A(n_1838),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_1902),
.Y(n_2093)
);

AO21x1_ASAP7_75t_L g2094 ( 
.A1(n_1957),
.A2(n_2001),
.B(n_1999),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1870),
.B(n_1984),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_1986),
.B(n_1936),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1952),
.B(n_1961),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1964),
.B(n_1965),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1909),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1925),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1990),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1941),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1955),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1993),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_1921),
.B(n_1948),
.Y(n_2105)
);

AOI22xp33_ASAP7_75t_SL g2106 ( 
.A1(n_1985),
.A2(n_1937),
.B1(n_1950),
.B2(n_1987),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1980),
.A2(n_1926),
.B1(n_1957),
.B2(n_1960),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1979),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_1929),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_1994),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_1994),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1838),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1974),
.Y(n_2113)
);

INVx4_ASAP7_75t_L g2114 ( 
.A(n_1892),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2013),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_2013),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1912),
.B(n_1949),
.Y(n_2117)
);

INVxp67_ASAP7_75t_L g2118 ( 
.A(n_1940),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2020),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_1929),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2020),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1876),
.B(n_1922),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1825),
.B(n_1989),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1856),
.B(n_1865),
.Y(n_2124)
);

AND2x4_ASAP7_75t_L g2125 ( 
.A(n_1870),
.B(n_1984),
.Y(n_2125)
);

OR2x6_ASAP7_75t_L g2126 ( 
.A(n_1933),
.B(n_1944),
.Y(n_2126)
);

HB1xp67_ASAP7_75t_L g2127 ( 
.A(n_1994),
.Y(n_2127)
);

AOI22xp33_ASAP7_75t_SL g2128 ( 
.A1(n_1950),
.A2(n_1942),
.B1(n_1939),
.B2(n_1886),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_SL g2129 ( 
.A1(n_2006),
.A2(n_1857),
.B(n_1928),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1849),
.B(n_1947),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1947),
.B(n_1956),
.Y(n_2131)
);

AO21x1_ASAP7_75t_L g2132 ( 
.A1(n_2001),
.A2(n_1992),
.B(n_1998),
.Y(n_2132)
);

BUFx2_ASAP7_75t_L g2133 ( 
.A(n_1886),
.Y(n_2133)
);

CKINVDCx11_ASAP7_75t_R g2134 ( 
.A(n_1859),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1856),
.B(n_1865),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2024),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2029),
.B(n_1842),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1988),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2029),
.B(n_1842),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1988),
.Y(n_2140)
);

OR2x2_ASAP7_75t_L g2141 ( 
.A(n_1828),
.B(n_1830),
.Y(n_2141)
);

OAI222xp33_ASAP7_75t_L g2142 ( 
.A1(n_2000),
.A2(n_1963),
.B1(n_1877),
.B2(n_1900),
.C1(n_1872),
.C2(n_2015),
.Y(n_2142)
);

AOI22xp5_ASAP7_75t_L g2143 ( 
.A1(n_1889),
.A2(n_1946),
.B1(n_1981),
.B2(n_1847),
.Y(n_2143)
);

OAI21x1_ASAP7_75t_L g2144 ( 
.A1(n_1850),
.A2(n_1871),
.B(n_1991),
.Y(n_2144)
);

OR2x2_ASAP7_75t_L g2145 ( 
.A(n_1831),
.B(n_1826),
.Y(n_2145)
);

NOR2xp33_ASAP7_75t_L g2146 ( 
.A(n_1917),
.B(n_2019),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_1934),
.B(n_1935),
.Y(n_2147)
);

BUFx8_ASAP7_75t_L g2148 ( 
.A(n_1914),
.Y(n_2148)
);

OR2x2_ASAP7_75t_L g2149 ( 
.A(n_1875),
.B(n_1890),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1968),
.B(n_1848),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_1894),
.Y(n_2151)
);

AO21x2_ASAP7_75t_L g2152 ( 
.A1(n_1893),
.A2(n_1906),
.B(n_1901),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1971),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1971),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1959),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1962),
.Y(n_2156)
);

OA21x2_ASAP7_75t_L g2157 ( 
.A1(n_1861),
.A2(n_1864),
.B(n_1873),
.Y(n_2157)
);

CKINVDCx11_ASAP7_75t_R g2158 ( 
.A(n_1872),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1927),
.Y(n_2159)
);

OR2x2_ASAP7_75t_L g2160 ( 
.A(n_1875),
.B(n_1890),
.Y(n_2160)
);

BUFx6f_ASAP7_75t_SL g2161 ( 
.A(n_1914),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_1973),
.Y(n_2162)
);

BUFx3_ASAP7_75t_L g2163 ( 
.A(n_2023),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1868),
.Y(n_2164)
);

OAI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1931),
.A2(n_1897),
.B1(n_1972),
.B2(n_1918),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_1899),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1868),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2039),
.B(n_2002),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2061),
.B(n_2002),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2061),
.B(n_2002),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2063),
.B(n_1848),
.Y(n_2171)
);

HB1xp67_ASAP7_75t_L g2172 ( 
.A(n_2076),
.Y(n_2172)
);

AND2x2_ASAP7_75t_L g2173 ( 
.A(n_2031),
.B(n_1997),
.Y(n_2173)
);

BUFx3_ASAP7_75t_L g2174 ( 
.A(n_2044),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_2044),
.Y(n_2175)
);

INVx4_ASAP7_75t_L g2176 ( 
.A(n_2126),
.Y(n_2176)
);

AOI22xp33_ASAP7_75t_L g2177 ( 
.A1(n_2040),
.A2(n_2028),
.B1(n_1837),
.B2(n_1982),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_2053),
.Y(n_2178)
);

CKINVDCx5p33_ASAP7_75t_R g2179 ( 
.A(n_2134),
.Y(n_2179)
);

OAI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_2066),
.A2(n_1975),
.B1(n_1978),
.B2(n_2023),
.C(n_2015),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2047),
.B(n_2017),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2071),
.Y(n_2182)
);

INVxp67_ASAP7_75t_L g2183 ( 
.A(n_2136),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2069),
.B(n_2017),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2113),
.Y(n_2185)
);

BUFx3_ASAP7_75t_L g2186 ( 
.A(n_2053),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_SL g2187 ( 
.A1(n_2114),
.A2(n_1945),
.B1(n_1918),
.B2(n_1891),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2068),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2082),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2038),
.Y(n_2190)
);

AND2x4_ASAP7_75t_L g2191 ( 
.A(n_2110),
.B(n_1996),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2041),
.B(n_2030),
.Y(n_2192)
);

NOR2x1_ASAP7_75t_L g2193 ( 
.A(n_2114),
.B(n_1945),
.Y(n_2193)
);

INVxp67_ASAP7_75t_L g2194 ( 
.A(n_2141),
.Y(n_2194)
);

BUFx2_ASAP7_75t_L g2195 ( 
.A(n_2043),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2089),
.Y(n_2196)
);

BUFx3_ASAP7_75t_L g2197 ( 
.A(n_2074),
.Y(n_2197)
);

NAND2x1_ASAP7_75t_L g2198 ( 
.A(n_2126),
.B(n_1930),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_R g2199 ( 
.A(n_2034),
.B(n_1851),
.Y(n_2199)
);

INVx4_ASAP7_75t_L g2200 ( 
.A(n_2126),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_2054),
.B(n_1967),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2033),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_2034),
.B(n_1888),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2042),
.B(n_1839),
.Y(n_2204)
);

OAI22xp33_ASAP7_75t_L g2205 ( 
.A1(n_2107),
.A2(n_1907),
.B1(n_1891),
.B2(n_1918),
.Y(n_2205)
);

INVx3_ASAP7_75t_L g2206 ( 
.A(n_2095),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2036),
.B(n_1983),
.Y(n_2207)
);

OAI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_2050),
.A2(n_1907),
.B1(n_1874),
.B2(n_1908),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_2045),
.B(n_1983),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2035),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2085),
.Y(n_2211)
);

INVx4_ASAP7_75t_R g2212 ( 
.A(n_2052),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2036),
.B(n_1983),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2056),
.B(n_1951),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2046),
.B(n_1951),
.Y(n_2215)
);

INVx4_ASAP7_75t_SL g2216 ( 
.A(n_2095),
.Y(n_2216)
);

INVx1_ASAP7_75t_SL g2217 ( 
.A(n_2134),
.Y(n_2217)
);

INVxp67_ASAP7_75t_SL g2218 ( 
.A(n_2043),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2049),
.B(n_1844),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_2037),
.B(n_1866),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_2108),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_2110),
.B(n_1866),
.Y(n_2222)
);

BUFx2_ASAP7_75t_L g2223 ( 
.A(n_2058),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2058),
.Y(n_2224)
);

INVx3_ASAP7_75t_L g2225 ( 
.A(n_2125),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2111),
.B(n_1867),
.Y(n_2226)
);

OAI222xp33_ASAP7_75t_L g2227 ( 
.A1(n_2066),
.A2(n_1863),
.B1(n_1908),
.B2(n_1898),
.C1(n_1879),
.C2(n_1883),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2152),
.Y(n_2228)
);

BUFx2_ASAP7_75t_SL g2229 ( 
.A(n_2161),
.Y(n_2229)
);

BUFx3_ASAP7_75t_L g2230 ( 
.A(n_2074),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_2127),
.B(n_1938),
.Y(n_2231)
);

BUFx3_ASAP7_75t_L g2232 ( 
.A(n_2087),
.Y(n_2232)
);

INVx4_ASAP7_75t_L g2233 ( 
.A(n_2075),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2055),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2099),
.Y(n_2235)
);

INVxp67_ASAP7_75t_L g2236 ( 
.A(n_2122),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2077),
.B(n_1867),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_2067),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2103),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2102),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_L g2241 ( 
.A1(n_2117),
.A2(n_1970),
.B1(n_1915),
.B2(n_1895),
.Y(n_2241)
);

HB1xp67_ASAP7_75t_L g2242 ( 
.A(n_2067),
.Y(n_2242)
);

HB1xp67_ASAP7_75t_L g2243 ( 
.A(n_2072),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2075),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2100),
.Y(n_2245)
);

HB1xp67_ASAP7_75t_L g2246 ( 
.A(n_2072),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2097),
.Y(n_2247)
);

BUFx2_ASAP7_75t_L g2248 ( 
.A(n_2166),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2080),
.Y(n_2249)
);

INVx4_ASAP7_75t_R g2250 ( 
.A(n_2079),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_2065),
.B(n_2014),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2097),
.Y(n_2252)
);

INVx3_ASAP7_75t_L g2253 ( 
.A(n_2088),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2096),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_2149),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2060),
.A2(n_1883),
.B1(n_1898),
.B2(n_1874),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2065),
.B(n_2021),
.Y(n_2257)
);

HB1xp67_ASAP7_75t_L g2258 ( 
.A(n_2160),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2131),
.B(n_2021),
.Y(n_2259)
);

HB1xp67_ASAP7_75t_L g2260 ( 
.A(n_2073),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_2181),
.B(n_2081),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2185),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2181),
.B(n_2171),
.Y(n_2263)
);

BUFx3_ASAP7_75t_L g2264 ( 
.A(n_2197),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2234),
.B(n_2059),
.Y(n_2265)
);

AOI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_2180),
.A2(n_2059),
.B1(n_2107),
.B2(n_2146),
.Y(n_2266)
);

BUFx4_ASAP7_75t_SL g2267 ( 
.A(n_2179),
.Y(n_2267)
);

OR2x6_ASAP7_75t_SL g2268 ( 
.A(n_2179),
.B(n_2032),
.Y(n_2268)
);

AND2x2_ASAP7_75t_L g2269 ( 
.A(n_2251),
.B(n_2257),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2251),
.B(n_2093),
.Y(n_2270)
);

HB1xp67_ASAP7_75t_L g2271 ( 
.A(n_2255),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2257),
.B(n_2093),
.Y(n_2272)
);

BUFx3_ASAP7_75t_L g2273 ( 
.A(n_2197),
.Y(n_2273)
);

HB1xp67_ASAP7_75t_L g2274 ( 
.A(n_2258),
.Y(n_2274)
);

AOI22xp33_ASAP7_75t_SL g2275 ( 
.A1(n_2176),
.A2(n_2078),
.B1(n_2090),
.B2(n_2133),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2169),
.B(n_2150),
.Y(n_2276)
);

AND2x2_ASAP7_75t_L g2277 ( 
.A(n_2169),
.B(n_2170),
.Y(n_2277)
);

OR2x6_ASAP7_75t_SL g2278 ( 
.A(n_2256),
.B(n_2057),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2170),
.B(n_2101),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_2195),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2249),
.Y(n_2281)
);

INVx1_ASAP7_75t_SL g2282 ( 
.A(n_2199),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_2231),
.B(n_2153),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2191),
.B(n_2154),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2249),
.Y(n_2285)
);

INVxp67_ASAP7_75t_L g2286 ( 
.A(n_2242),
.Y(n_2286)
);

HB1xp67_ASAP7_75t_L g2287 ( 
.A(n_2223),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2196),
.B(n_2190),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2201),
.Y(n_2289)
);

INVxp67_ASAP7_75t_SL g2290 ( 
.A(n_2218),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2176),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_2254),
.B(n_2182),
.Y(n_2292)
);

INVx3_ASAP7_75t_L g2293 ( 
.A(n_2176),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2219),
.B(n_2130),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2239),
.B(n_2105),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2221),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2184),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2240),
.B(n_2118),
.Y(n_2298)
);

NAND2x1p5_ASAP7_75t_L g2299 ( 
.A(n_2200),
.B(n_2073),
.Y(n_2299)
);

HB1xp67_ASAP7_75t_L g2300 ( 
.A(n_2224),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2184),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2214),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2209),
.B(n_2165),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2168),
.B(n_2132),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_2230),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2202),
.B(n_2118),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2210),
.B(n_2138),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2173),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2191),
.B(n_2155),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2168),
.B(n_2156),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2245),
.B(n_2172),
.Y(n_2311)
);

AND2x4_ASAP7_75t_L g2312 ( 
.A(n_2191),
.B(n_2144),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_2229),
.Y(n_2313)
);

HB1xp67_ASAP7_75t_L g2314 ( 
.A(n_2243),
.Y(n_2314)
);

BUFx2_ASAP7_75t_L g2315 ( 
.A(n_2248),
.Y(n_2315)
);

AND2x4_ASAP7_75t_SL g2316 ( 
.A(n_2233),
.B(n_2147),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2192),
.B(n_2157),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2192),
.B(n_2157),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2269),
.B(n_2222),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2269),
.B(n_2222),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_2282),
.B(n_2217),
.Y(n_2321)
);

INVx3_ASAP7_75t_R g2322 ( 
.A(n_2315),
.Y(n_2322)
);

OR2x2_ASAP7_75t_L g2323 ( 
.A(n_2297),
.B(n_2207),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2271),
.B(n_2188),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2281),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2297),
.B(n_2207),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2314),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2263),
.B(n_2226),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2262),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2263),
.B(n_2226),
.Y(n_2330)
);

AND2x2_ASAP7_75t_L g2331 ( 
.A(n_2303),
.B(n_2259),
.Y(n_2331)
);

OR2x2_ASAP7_75t_L g2332 ( 
.A(n_2301),
.B(n_2213),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2289),
.B(n_2259),
.Y(n_2333)
);

AND2x4_ASAP7_75t_L g2334 ( 
.A(n_2312),
.B(n_2228),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2281),
.Y(n_2335)
);

HB1xp67_ASAP7_75t_L g2336 ( 
.A(n_2274),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2303),
.B(n_2215),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2285),
.Y(n_2338)
);

CKINVDCx5p33_ASAP7_75t_R g2339 ( 
.A(n_2267),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2285),
.Y(n_2340)
);

HB1xp67_ASAP7_75t_L g2341 ( 
.A(n_2280),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2296),
.Y(n_2342)
);

AND2x2_ASAP7_75t_L g2343 ( 
.A(n_2304),
.B(n_2215),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2289),
.B(n_2237),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2292),
.B(n_2189),
.Y(n_2345)
);

INVx3_ASAP7_75t_L g2346 ( 
.A(n_2312),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2304),
.B(n_2276),
.Y(n_2347)
);

NAND2x1_ASAP7_75t_SL g2348 ( 
.A(n_2291),
.B(n_2200),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_2276),
.B(n_2220),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2279),
.B(n_2235),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2294),
.B(n_2220),
.Y(n_2351)
);

AND3x2_ASAP7_75t_L g2352 ( 
.A(n_2286),
.B(n_2203),
.C(n_2238),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_2313),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2279),
.B(n_2311),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2294),
.B(n_2237),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2264),
.Y(n_2356)
);

INVxp67_ASAP7_75t_SL g2357 ( 
.A(n_2290),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2270),
.B(n_2204),
.Y(n_2358)
);

HB1xp67_ASAP7_75t_L g2359 ( 
.A(n_2327),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2356),
.B(n_2313),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2346),
.B(n_2312),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_2346),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2325),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2324),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2325),
.Y(n_2365)
);

AOI21xp33_ASAP7_75t_L g2366 ( 
.A1(n_2336),
.A2(n_2104),
.B(n_2146),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2341),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2346),
.B(n_2284),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2347),
.B(n_2261),
.Y(n_2369)
);

NAND3xp33_ASAP7_75t_L g2370 ( 
.A(n_2352),
.B(n_2266),
.C(n_2183),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2335),
.Y(n_2371)
);

INVx1_ASAP7_75t_L g2372 ( 
.A(n_2335),
.Y(n_2372)
);

OAI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2357),
.A2(n_2275),
.B(n_2142),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2329),
.Y(n_2374)
);

OR2x2_ASAP7_75t_L g2375 ( 
.A(n_2319),
.B(n_2308),
.Y(n_2375)
);

NAND2x1p5_ASAP7_75t_L g2376 ( 
.A(n_2356),
.B(n_2200),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2319),
.B(n_2317),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2347),
.B(n_2261),
.Y(n_2378)
);

NAND4xp75_ASAP7_75t_L g2379 ( 
.A(n_2321),
.B(n_2193),
.C(n_2084),
.D(n_2094),
.Y(n_2379)
);

HB1xp67_ASAP7_75t_L g2380 ( 
.A(n_2322),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_2348),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2346),
.B(n_2284),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2329),
.Y(n_2383)
);

AND2x4_ASAP7_75t_L g2384 ( 
.A(n_2334),
.B(n_2284),
.Y(n_2384)
);

HB1xp67_ASAP7_75t_L g2385 ( 
.A(n_2322),
.Y(n_2385)
);

AND2x4_ASAP7_75t_L g2386 ( 
.A(n_2334),
.B(n_2284),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2320),
.B(n_2317),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_2329),
.Y(n_2388)
);

AND2x2_ASAP7_75t_L g2389 ( 
.A(n_2320),
.B(n_2318),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2343),
.B(n_2270),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2353),
.B(n_2264),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2350),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2338),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2343),
.B(n_2272),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2328),
.B(n_2318),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2331),
.B(n_2272),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2323),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_2331),
.B(n_2355),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2355),
.B(n_2288),
.Y(n_2399)
);

OR2x2_ASAP7_75t_L g2400 ( 
.A(n_2375),
.B(n_2354),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2377),
.B(n_2328),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2397),
.B(n_2337),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2375),
.Y(n_2403)
);

OR2x2_ASAP7_75t_L g2404 ( 
.A(n_2399),
.B(n_2330),
.Y(n_2404)
);

OAI22xp33_ASAP7_75t_L g2405 ( 
.A1(n_2380),
.A2(n_2278),
.B1(n_2305),
.B2(n_2273),
.Y(n_2405)
);

OAI33xp33_ASAP7_75t_L g2406 ( 
.A1(n_2364),
.A2(n_2345),
.A3(n_2295),
.B1(n_2194),
.B2(n_2344),
.B3(n_2333),
.Y(n_2406)
);

INVx1_ASAP7_75t_SL g2407 ( 
.A(n_2391),
.Y(n_2407)
);

AOI222xp33_ASAP7_75t_L g2408 ( 
.A1(n_2370),
.A2(n_2236),
.B1(n_2211),
.B2(n_2140),
.C1(n_2306),
.C2(n_2298),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2359),
.B(n_2367),
.Y(n_2409)
);

NOR2xp33_ASAP7_75t_L g2410 ( 
.A(n_2392),
.B(n_2162),
.Y(n_2410)
);

INVx2_ASAP7_75t_L g2411 ( 
.A(n_2374),
.Y(n_2411)
);

AND2x2_ASAP7_75t_L g2412 ( 
.A(n_2377),
.B(n_2330),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_L g2413 ( 
.A(n_2398),
.B(n_2337),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2385),
.B(n_2273),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2363),
.Y(n_2415)
);

OR2x2_ASAP7_75t_L g2416 ( 
.A(n_2369),
.B(n_2323),
.Y(n_2416)
);

OAI32xp33_ASAP7_75t_L g2417 ( 
.A1(n_2376),
.A2(n_2278),
.A3(n_2268),
.B1(n_2305),
.B2(n_2299),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2363),
.Y(n_2418)
);

OR2x2_ASAP7_75t_L g2419 ( 
.A(n_2378),
.B(n_2326),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2365),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2387),
.B(n_2351),
.Y(n_2421)
);

OAI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2360),
.A2(n_2128),
.B1(n_2299),
.B2(n_2060),
.Y(n_2422)
);

AOI21xp33_ASAP7_75t_L g2423 ( 
.A1(n_2373),
.A2(n_2145),
.B(n_2151),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2374),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2387),
.B(n_2351),
.Y(n_2425)
);

O2A1O1Ixp5_ASAP7_75t_L g2426 ( 
.A1(n_2362),
.A2(n_2198),
.B(n_2142),
.C(n_2233),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2365),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2389),
.B(n_2358),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2371),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2389),
.B(n_2358),
.Y(n_2430)
);

AOI211xp5_ASAP7_75t_L g2431 ( 
.A1(n_2366),
.A2(n_2227),
.B(n_2205),
.C(n_2339),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2395),
.B(n_2349),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2396),
.B(n_2268),
.Y(n_2433)
);

OAI22xp5_ASAP7_75t_L g2434 ( 
.A1(n_2376),
.A2(n_2128),
.B1(n_2299),
.B2(n_2316),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2390),
.B(n_2086),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2415),
.Y(n_2436)
);

XOR2x2_ASAP7_75t_L g2437 ( 
.A(n_2433),
.B(n_2083),
.Y(n_2437)
);

AOI21xp5_ASAP7_75t_L g2438 ( 
.A1(n_2417),
.A2(n_2381),
.B(n_2376),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2411),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2418),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2420),
.Y(n_2441)
);

O2A1O1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_2422),
.A2(n_2048),
.B(n_2159),
.C(n_2307),
.Y(n_2442)
);

OAI21xp5_ASAP7_75t_L g2443 ( 
.A1(n_2426),
.A2(n_2379),
.B(n_2048),
.Y(n_2443)
);

NOR2x1_ASAP7_75t_L g2444 ( 
.A(n_2405),
.B(n_2379),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2416),
.B(n_2419),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2427),
.Y(n_2446)
);

INVxp67_ASAP7_75t_L g2447 ( 
.A(n_2407),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2429),
.Y(n_2448)
);

OAI22xp5_ASAP7_75t_L g2449 ( 
.A1(n_2405),
.A2(n_2381),
.B1(n_2362),
.B2(n_2368),
.Y(n_2449)
);

NAND3x1_ASAP7_75t_L g2450 ( 
.A(n_2433),
.B(n_2362),
.C(n_2293),
.Y(n_2450)
);

O2A1O1Ixp33_ASAP7_75t_SL g2451 ( 
.A1(n_2414),
.A2(n_2394),
.B(n_2246),
.C(n_2250),
.Y(n_2451)
);

AOI221xp5_ASAP7_75t_L g2452 ( 
.A1(n_2406),
.A2(n_2395),
.B1(n_2361),
.B2(n_2371),
.C(n_2393),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2403),
.Y(n_2453)
);

OAI22xp33_ASAP7_75t_L g2454 ( 
.A1(n_2434),
.A2(n_2293),
.B1(n_2291),
.B2(n_2326),
.Y(n_2454)
);

AOI22xp33_ASAP7_75t_L g2455 ( 
.A1(n_2423),
.A2(n_2361),
.B1(n_2382),
.B2(n_2368),
.Y(n_2455)
);

NOR3xp33_ASAP7_75t_L g2456 ( 
.A(n_2443),
.B(n_1862),
.C(n_2158),
.Y(n_2456)
);

AOI21xp5_ASAP7_75t_L g2457 ( 
.A1(n_2451),
.A2(n_2414),
.B(n_2408),
.Y(n_2457)
);

OAI211xp5_ASAP7_75t_L g2458 ( 
.A1(n_2443),
.A2(n_2158),
.B(n_2431),
.C(n_2106),
.Y(n_2458)
);

INVxp67_ASAP7_75t_L g2459 ( 
.A(n_2437),
.Y(n_2459)
);

AOI221xp5_ASAP7_75t_L g2460 ( 
.A1(n_2449),
.A2(n_2410),
.B1(n_2435),
.B2(n_2409),
.C(n_2402),
.Y(n_2460)
);

OAI221xp5_ASAP7_75t_L g2461 ( 
.A1(n_2444),
.A2(n_2449),
.B1(n_2442),
.B2(n_2455),
.C(n_2438),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2445),
.Y(n_2462)
);

AOI221xp5_ASAP7_75t_L g2463 ( 
.A1(n_2452),
.A2(n_2410),
.B1(n_2435),
.B2(n_2413),
.C(n_2425),
.Y(n_2463)
);

AO21x1_ASAP7_75t_L g2464 ( 
.A1(n_2454),
.A2(n_2233),
.B(n_2316),
.Y(n_2464)
);

AOI222xp33_ASAP7_75t_L g2465 ( 
.A1(n_2447),
.A2(n_2425),
.B1(n_2161),
.B2(n_2428),
.C1(n_2430),
.C2(n_2401),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2436),
.Y(n_2466)
);

AOI221xp5_ASAP7_75t_L g2467 ( 
.A1(n_2453),
.A2(n_2432),
.B1(n_2412),
.B2(n_2421),
.C(n_2361),
.Y(n_2467)
);

OAI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2450),
.A2(n_2143),
.B(n_2187),
.Y(n_2468)
);

OAI211xp5_ASAP7_75t_L g2469 ( 
.A1(n_2440),
.A2(n_2106),
.B(n_2064),
.C(n_2348),
.Y(n_2469)
);

AOI22xp5_ASAP7_75t_L g2470 ( 
.A1(n_2441),
.A2(n_2382),
.B1(n_2368),
.B2(n_2384),
.Y(n_2470)
);

OAI211xp5_ASAP7_75t_L g2471 ( 
.A1(n_2446),
.A2(n_2177),
.B(n_2265),
.C(n_2241),
.Y(n_2471)
);

OAI22xp5_ASAP7_75t_L g2472 ( 
.A1(n_2448),
.A2(n_2400),
.B1(n_2404),
.B2(n_2382),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2439),
.B(n_2411),
.Y(n_2473)
);

AOI221xp5_ASAP7_75t_L g2474 ( 
.A1(n_2449),
.A2(n_2424),
.B1(n_2393),
.B2(n_2372),
.C(n_2344),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2452),
.B(n_2424),
.Y(n_2475)
);

AOI32xp33_ASAP7_75t_L g2476 ( 
.A1(n_2444),
.A2(n_2386),
.A3(n_2384),
.B1(n_2230),
.B2(n_2232),
.Y(n_2476)
);

OAI21xp33_ASAP7_75t_L g2477 ( 
.A1(n_2444),
.A2(n_2333),
.B(n_2384),
.Y(n_2477)
);

OA21x2_ASAP7_75t_L g2478 ( 
.A1(n_2443),
.A2(n_2383),
.B(n_2388),
.Y(n_2478)
);

NOR4xp25_ASAP7_75t_SL g2479 ( 
.A(n_2451),
.B(n_2016),
.C(n_1851),
.D(n_2083),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2462),
.B(n_2372),
.Y(n_2480)
);

AOI221xp5_ASAP7_75t_L g2481 ( 
.A1(n_2461),
.A2(n_2386),
.B1(n_2300),
.B2(n_2287),
.C(n_2315),
.Y(n_2481)
);

AOI222xp33_ASAP7_75t_L g2482 ( 
.A1(n_2459),
.A2(n_2062),
.B1(n_2148),
.B2(n_2302),
.C1(n_2252),
.C2(n_2247),
.Y(n_2482)
);

AO22x1_ASAP7_75t_L g2483 ( 
.A1(n_2456),
.A2(n_2148),
.B1(n_2175),
.B2(n_2174),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2463),
.B(n_2349),
.Y(n_2484)
);

OAI21xp33_ASAP7_75t_SL g2485 ( 
.A1(n_2476),
.A2(n_2293),
.B(n_2291),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_2464),
.B(n_2386),
.Y(n_2486)
);

NAND2x1_ASAP7_75t_L g2487 ( 
.A(n_2478),
.B(n_2212),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_SL g2488 ( 
.A(n_2457),
.B(n_2016),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2475),
.B(n_2277),
.Y(n_2489)
);

NOR4xp25_ASAP7_75t_L g2490 ( 
.A(n_2458),
.B(n_2123),
.C(n_2115),
.D(n_2121),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2466),
.Y(n_2491)
);

NAND4xp25_ASAP7_75t_L g2492 ( 
.A(n_2465),
.B(n_2163),
.C(n_2139),
.D(n_2137),
.Y(n_2492)
);

NOR3xp33_ASAP7_75t_SL g2493 ( 
.A(n_2469),
.B(n_2477),
.C(n_2460),
.Y(n_2493)
);

NAND4xp25_ASAP7_75t_L g2494 ( 
.A(n_2468),
.B(n_2163),
.C(n_2175),
.D(n_2174),
.Y(n_2494)
);

NAND5xp2_ASAP7_75t_L g2495 ( 
.A(n_2474),
.B(n_2051),
.C(n_2010),
.D(n_1896),
.E(n_2088),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2467),
.B(n_2277),
.Y(n_2496)
);

NOR2xp33_ASAP7_75t_L g2497 ( 
.A(n_2472),
.B(n_2051),
.Y(n_2497)
);

INVxp67_ASAP7_75t_SL g2498 ( 
.A(n_2488),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2480),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_SL g2500 ( 
.A(n_2481),
.B(n_2470),
.Y(n_2500)
);

NOR2xp67_ASAP7_75t_L g2501 ( 
.A(n_2485),
.B(n_2486),
.Y(n_2501)
);

NOR2x1_ASAP7_75t_L g2502 ( 
.A(n_2495),
.B(n_2478),
.Y(n_2502)
);

NOR3xp33_ASAP7_75t_L g2503 ( 
.A(n_2483),
.B(n_2471),
.C(n_2473),
.Y(n_2503)
);

NAND3xp33_ASAP7_75t_L g2504 ( 
.A(n_2493),
.B(n_2479),
.C(n_2119),
.Y(n_2504)
);

NOR3x1_ASAP7_75t_L g2505 ( 
.A(n_2492),
.B(n_1911),
.C(n_1977),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2489),
.B(n_2383),
.Y(n_2506)
);

AOI22xp5_ASAP7_75t_L g2507 ( 
.A1(n_2497),
.A2(n_2334),
.B1(n_2309),
.B2(n_2283),
.Y(n_2507)
);

NAND3xp33_ASAP7_75t_SL g2508 ( 
.A(n_2490),
.B(n_2482),
.C(n_2487),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2496),
.B(n_2334),
.Y(n_2509)
);

NOR2x1_ASAP7_75t_L g2510 ( 
.A(n_2494),
.B(n_2087),
.Y(n_2510)
);

NOR3xp33_ASAP7_75t_L g2511 ( 
.A(n_2484),
.B(n_2135),
.C(n_2124),
.Y(n_2511)
);

AOI211x1_ASAP7_75t_L g2512 ( 
.A1(n_2491),
.A2(n_2338),
.B(n_2342),
.C(n_2340),
.Y(n_2512)
);

AND3x2_ASAP7_75t_L g2513 ( 
.A(n_2498),
.B(n_1932),
.C(n_2260),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2511),
.B(n_2388),
.Y(n_2514)
);

NAND4xp25_ASAP7_75t_L g2515 ( 
.A(n_2505),
.B(n_2120),
.C(n_2109),
.D(n_2178),
.Y(n_2515)
);

NOR3xp33_ASAP7_75t_L g2516 ( 
.A(n_2508),
.B(n_2091),
.C(n_2109),
.Y(n_2516)
);

AND2x2_ASAP7_75t_L g2517 ( 
.A(n_2502),
.B(n_2310),
.Y(n_2517)
);

NOR3xp33_ASAP7_75t_L g2518 ( 
.A(n_2504),
.B(n_2503),
.C(n_2500),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2509),
.B(n_2310),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2501),
.B(n_1833),
.Y(n_2520)
);

NAND4xp75_ASAP7_75t_L g2521 ( 
.A(n_2510),
.B(n_1833),
.C(n_2070),
.D(n_2098),
.Y(n_2521)
);

OAI211xp5_ASAP7_75t_L g2522 ( 
.A1(n_2499),
.A2(n_2120),
.B(n_1833),
.C(n_2232),
.Y(n_2522)
);

HB1xp67_ASAP7_75t_L g2523 ( 
.A(n_2506),
.Y(n_2523)
);

NOR3x1_ASAP7_75t_L g2524 ( 
.A(n_2512),
.B(n_2090),
.C(n_2208),
.Y(n_2524)
);

NOR4xp25_ASAP7_75t_L g2525 ( 
.A(n_2507),
.B(n_1879),
.C(n_2167),
.D(n_2164),
.Y(n_2525)
);

BUFx8_ASAP7_75t_SL g2526 ( 
.A(n_2513),
.Y(n_2526)
);

NOR3xp33_ASAP7_75t_L g2527 ( 
.A(n_2520),
.B(n_2091),
.C(n_2116),
.Y(n_2527)
);

NOR2x1_ASAP7_75t_SL g2528 ( 
.A(n_2522),
.B(n_2178),
.Y(n_2528)
);

OR2x2_ASAP7_75t_L g2529 ( 
.A(n_2514),
.B(n_2332),
.Y(n_2529)
);

NAND4xp75_ASAP7_75t_L g2530 ( 
.A(n_2524),
.B(n_2098),
.C(n_2070),
.D(n_1884),
.Y(n_2530)
);

INVx2_ASAP7_75t_L g2531 ( 
.A(n_2521),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2518),
.A2(n_2186),
.B1(n_2225),
.B2(n_2206),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2523),
.B(n_2340),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2516),
.Y(n_2534)
);

OAI21xp5_ASAP7_75t_L g2535 ( 
.A1(n_2517),
.A2(n_1966),
.B(n_1958),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_2526),
.Y(n_2536)
);

XOR2x1_ASAP7_75t_L g2537 ( 
.A(n_2531),
.B(n_2519),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2533),
.Y(n_2538)
);

OAI31xp67_ASAP7_75t_L g2539 ( 
.A1(n_2530),
.A2(n_2515),
.A3(n_2525),
.B(n_2522),
.Y(n_2539)
);

OA22x2_ASAP7_75t_L g2540 ( 
.A1(n_2534),
.A2(n_2129),
.B1(n_2244),
.B2(n_2253),
.Y(n_2540)
);

OAI22xp5_ASAP7_75t_SL g2541 ( 
.A1(n_2532),
.A2(n_2186),
.B1(n_1995),
.B2(n_2253),
.Y(n_2541)
);

INVx2_ASAP7_75t_SL g2542 ( 
.A(n_2529),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2528),
.Y(n_2543)
);

AND2x2_ASAP7_75t_SL g2544 ( 
.A(n_2527),
.B(n_1953),
.Y(n_2544)
);

AO21x2_ASAP7_75t_L g2545 ( 
.A1(n_2538),
.A2(n_2543),
.B(n_2537),
.Y(n_2545)
);

XOR2x2_ASAP7_75t_L g2546 ( 
.A(n_2536),
.B(n_2542),
.Y(n_2546)
);

INVxp67_ASAP7_75t_SL g2547 ( 
.A(n_2536),
.Y(n_2547)
);

XNOR2x1_ASAP7_75t_SL g2548 ( 
.A(n_2539),
.B(n_2535),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2547),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2546),
.Y(n_2550)
);

XNOR2x1_ASAP7_75t_L g2551 ( 
.A(n_2548),
.B(n_2540),
.Y(n_2551)
);

AOI21xp33_ASAP7_75t_L g2552 ( 
.A1(n_2545),
.A2(n_2544),
.B(n_2541),
.Y(n_2552)
);

AOI21xp5_ASAP7_75t_L g2553 ( 
.A1(n_2545),
.A2(n_2535),
.B(n_1966),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2549),
.Y(n_2554)
);

AOI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2551),
.A2(n_1953),
.B(n_1930),
.Y(n_2555)
);

AOI21xp5_ASAP7_75t_L g2556 ( 
.A1(n_2552),
.A2(n_1953),
.B(n_1930),
.Y(n_2556)
);

AO21x2_ASAP7_75t_L g2557 ( 
.A1(n_2554),
.A2(n_2550),
.B(n_2553),
.Y(n_2557)
);

AO22x2_ASAP7_75t_L g2558 ( 
.A1(n_2556),
.A2(n_2555),
.B1(n_2216),
.B2(n_2116),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2554),
.B(n_1995),
.Y(n_2559)
);

OAI21x1_ASAP7_75t_L g2560 ( 
.A1(n_2559),
.A2(n_2112),
.B(n_2092),
.Y(n_2560)
);

INVxp67_ASAP7_75t_L g2561 ( 
.A(n_2560),
.Y(n_2561)
);

INVxp67_ASAP7_75t_L g2562 ( 
.A(n_2561),
.Y(n_2562)
);

AOI22xp5_ASAP7_75t_L g2563 ( 
.A1(n_2562),
.A2(n_2557),
.B1(n_2558),
.B2(n_2092),
.Y(n_2563)
);


endmodule