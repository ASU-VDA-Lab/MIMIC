module fake_netlist_6_1215_n_725 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_725);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_725;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_58),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_57),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_34),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_67),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_54),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_33),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_6),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_90),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_16),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_21),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_108),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_120),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_7),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_94),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_62),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_48),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_46),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_71),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_24),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_98),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_92),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_65),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_93),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_73),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_29),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_160),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

NAND2xp33_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_0),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_157),
.B(n_2),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_178),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_3),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

AND2x6_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_19),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_167),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_157),
.B(n_5),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_193),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

BUFx8_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_176),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_181),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_162),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_8),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_235),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_191),
.B(n_166),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

NAND2xp33_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_188),
.Y(n_249)
);

NAND2xp33_ASAP7_75t_L g250 ( 
.A(n_216),
.B(n_191),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_154),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_226),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

AND3x2_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_168),
.C(n_201),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_164),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_211),
.Y(n_263)
);

INVxp67_ASAP7_75t_R g264 ( 
.A(n_211),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_204),
.A2(n_198),
.B1(n_172),
.B2(n_185),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_221),
.B(n_156),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_L g267 ( 
.A(n_210),
.B(n_177),
.C(n_180),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_214),
.B(n_189),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_235),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_194),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_209),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_200),
.B1(n_199),
.B2(n_197),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_196),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g279 ( 
.A(n_224),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_209),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_209),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_150),
.Y(n_283)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_215),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_239),
.B(n_195),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_243),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_267),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_219),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_220),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_266),
.B(n_212),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_263),
.B(n_231),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_225),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_230),
.Y(n_300)
);

O2A1O1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_268),
.A2(n_210),
.B(n_240),
.C(n_207),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_263),
.B(n_153),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_241),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_274),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_205),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_250),
.B(n_215),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_274),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_265),
.B(n_169),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_206),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_259),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_262),
.B(n_207),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_253),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_281),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_279),
.A2(n_221),
.B1(n_237),
.B2(n_228),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_244),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_244),
.B(n_227),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_228),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_260),
.A2(n_221),
.B(n_173),
.C(n_187),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_244),
.B(n_228),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_284),
.B(n_174),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_179),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_249),
.A2(n_264),
.B1(n_279),
.B2(n_283),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_264),
.A2(n_192),
.B1(n_186),
.B2(n_184),
.Y(n_329)
);

AND2x2_ASAP7_75t_SL g330 ( 
.A(n_260),
.B(n_234),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_282),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_258),
.B(n_234),
.Y(n_332)
);

O2A1O1Ixp5_ASAP7_75t_L g333 ( 
.A1(n_247),
.A2(n_234),
.B(n_64),
.C(n_66),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_258),
.B(n_213),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_284),
.B(n_257),
.Y(n_335)
);

AND3x1_ASAP7_75t_L g336 ( 
.A(n_245),
.B(n_213),
.C(n_10),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_248),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_284),
.B(n_20),
.Y(n_340)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_245),
.B(n_9),
.C(n_10),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_308),
.A2(n_280),
.B(n_273),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_280),
.Y(n_343)
);

OA22x2_ASAP7_75t_L g344 ( 
.A1(n_327),
.A2(n_252),
.B1(n_255),
.B2(n_12),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_293),
.A2(n_273),
.B(n_248),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_273),
.B(n_248),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_292),
.B(n_278),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_302),
.B(n_9),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_320),
.A2(n_255),
.B1(n_252),
.B2(n_278),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_257),
.B1(n_273),
.B2(n_251),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_310),
.A2(n_273),
.B1(n_251),
.B2(n_247),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_11),
.Y(n_353)
);

INVx11_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_320),
.A2(n_251),
.B1(n_70),
.B2(n_72),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_303),
.Y(n_356)
);

O2A1O1Ixp33_ASAP7_75t_L g357 ( 
.A1(n_297),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_290),
.A2(n_251),
.B1(n_14),
.B2(n_15),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_303),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_297),
.A2(n_74),
.B(n_145),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_288),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_333),
.A2(n_68),
.B(n_144),
.Y(n_362)
);

OR2x6_ASAP7_75t_SL g363 ( 
.A(n_341),
.B(n_13),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_15),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_299),
.Y(n_365)
);

A2O1A1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_314),
.A2(n_301),
.B(n_307),
.C(n_312),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_22),
.Y(n_367)
);

AO21x1_ASAP7_75t_L g368 ( 
.A1(n_340),
.A2(n_16),
.B(n_17),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_329),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_307),
.B(n_23),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_290),
.A2(n_78),
.B1(n_143),
.B2(n_25),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_26),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_340),
.A2(n_317),
.B1(n_330),
.B2(n_325),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_287),
.B(n_27),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_325),
.A2(n_79),
.B(n_140),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_321),
.A2(n_76),
.B(n_138),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_316),
.B(n_28),
.Y(n_377)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_336),
.B(n_17),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_309),
.B(n_18),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_287),
.B(n_18),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_299),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_332),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_317),
.B(n_30),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_334),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_312),
.B(n_31),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_289),
.Y(n_387)
);

BUFx12f_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_296),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_389)
);

AOI21xp33_ASAP7_75t_L g390 ( 
.A1(n_295),
.A2(n_146),
.B(n_38),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_324),
.B(n_37),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_305),
.B(n_39),
.Y(n_392)
);

AO21x1_ASAP7_75t_L g393 ( 
.A1(n_328),
.A2(n_339),
.B(n_331),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_SL g394 ( 
.A(n_291),
.B(n_298),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_300),
.Y(n_395)
);

AO21x1_ASAP7_75t_L g396 ( 
.A1(n_337),
.A2(n_40),
.B(n_41),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_319),
.A2(n_43),
.B(n_44),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_326),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_399)
);

NOR2x1p5_ASAP7_75t_SL g400 ( 
.A(n_315),
.B(n_50),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_322),
.A2(n_51),
.B(n_52),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_323),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_323),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_373),
.Y(n_404)
);

CKINVDCx11_ASAP7_75t_R g405 ( 
.A(n_388),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_385),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_379),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_338),
.B1(n_294),
.B2(n_315),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_299),
.Y(n_409)
);

CKINVDCx11_ASAP7_75t_R g410 ( 
.A(n_363),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_347),
.B(n_53),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_365),
.A2(n_55),
.B(n_56),
.Y(n_412)
);

NOR2x1_ASAP7_75t_SL g413 ( 
.A(n_372),
.B(n_59),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_382),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_365),
.A2(n_60),
.B(n_63),
.Y(n_415)
);

NAND2x1_ASAP7_75t_L g416 ( 
.A(n_381),
.B(n_75),
.Y(n_416)
);

OA22x2_ASAP7_75t_L g417 ( 
.A1(n_358),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_387),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_370),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

AO31x2_ASAP7_75t_L g423 ( 
.A1(n_368),
.A2(n_84),
.A3(n_88),
.B(n_89),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_95),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_348),
.B(n_353),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_354),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_369),
.B(n_99),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_345),
.A2(n_100),
.B(n_102),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_SL g429 ( 
.A(n_358),
.B(n_105),
.C(n_106),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_359),
.B(n_107),
.Y(n_430)
);

AO21x2_ASAP7_75t_L g431 ( 
.A1(n_376),
.A2(n_135),
.B(n_111),
.Y(n_431)
);

AO31x2_ASAP7_75t_L g432 ( 
.A1(n_396),
.A2(n_110),
.A3(n_112),
.B(n_113),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_374),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_359),
.B(n_383),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_359),
.Y(n_436)
);

NAND2x1p5_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_115),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_344),
.B(n_117),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_343),
.A2(n_118),
.B(n_121),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_397),
.Y(n_440)
);

AOI211x1_ASAP7_75t_L g441 ( 
.A1(n_375),
.A2(n_122),
.B(n_124),
.C(n_125),
.Y(n_441)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_346),
.A2(n_134),
.B(n_130),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_380),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_349),
.B(n_133),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_127),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_378),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_342),
.A2(n_132),
.B(n_362),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_400),
.B(n_355),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_352),
.A2(n_360),
.B(n_350),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_398),
.A2(n_401),
.B(n_399),
.Y(n_450)
);

OAI22xp33_ASAP7_75t_L g451 ( 
.A1(n_417),
.A2(n_371),
.B1(n_390),
.B2(n_357),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_404),
.A2(n_389),
.B(n_392),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_426),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_414),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_367),
.Y(n_455)
);

OA21x2_ASAP7_75t_L g456 ( 
.A1(n_447),
.A2(n_404),
.B(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_406),
.Y(n_457)
);

A2O1A1Ixp33_ASAP7_75t_L g458 ( 
.A1(n_425),
.A2(n_443),
.B(n_421),
.C(n_449),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_446),
.Y(n_459)
);

OAI21x1_ASAP7_75t_SL g460 ( 
.A1(n_413),
.A2(n_403),
.B(n_439),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_433),
.Y(n_461)
);

AND2x4_ASAP7_75t_L g462 ( 
.A(n_418),
.B(n_436),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_422),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_421),
.B(n_403),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_409),
.Y(n_465)
);

AOI21xp33_ASAP7_75t_L g466 ( 
.A1(n_444),
.A2(n_431),
.B(n_427),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_436),
.B(n_416),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_419),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_448),
.A2(n_411),
.B(n_450),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_406),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_435),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_434),
.Y(n_473)
);

AO31x2_ASAP7_75t_L g474 ( 
.A1(n_445),
.A2(n_424),
.A3(n_430),
.B(n_412),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_407),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

OAI211xp5_ASAP7_75t_SL g477 ( 
.A1(n_407),
.A2(n_410),
.B(n_408),
.C(n_445),
.Y(n_477)
);

OAI222xp33_ASAP7_75t_L g478 ( 
.A1(n_438),
.A2(n_437),
.B1(n_429),
.B2(n_441),
.C1(n_415),
.C2(n_431),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_428),
.A2(n_442),
.B(n_423),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_446),
.Y(n_480)
);

INVx8_ASAP7_75t_L g481 ( 
.A(n_446),
.Y(n_481)
);

AO21x2_ASAP7_75t_L g482 ( 
.A1(n_432),
.A2(n_423),
.B(n_405),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_432),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_432),
.A2(n_404),
.B(n_402),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_404),
.A2(n_384),
.B1(n_373),
.B2(n_443),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_414),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_436),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_404),
.A2(n_384),
.B1(n_373),
.B2(n_443),
.Y(n_489)
);

INVx4_ASAP7_75t_SL g490 ( 
.A(n_423),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_404),
.A2(n_448),
.B(n_402),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_419),
.Y(n_492)
);

AO31x2_ASAP7_75t_L g493 ( 
.A1(n_404),
.A2(n_393),
.A3(n_448),
.B(n_421),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_405),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_470),
.Y(n_496)
);

OR2x2_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_459),
.Y(n_497)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_453),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_457),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_462),
.B(n_480),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_454),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_488),
.Y(n_503)
);

AOI221xp5_ASAP7_75t_L g504 ( 
.A1(n_485),
.A2(n_489),
.B1(n_451),
.B2(n_466),
.C(n_478),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_463),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

AO21x2_ASAP7_75t_L g507 ( 
.A1(n_469),
.A2(n_484),
.B(n_466),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_495),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_472),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_495),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_473),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_491),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_481),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_481),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

BUFx4f_ASAP7_75t_SL g518 ( 
.A(n_461),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_486),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_492),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_488),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_462),
.Y(n_523)
);

INVx4_ASAP7_75t_L g524 ( 
.A(n_481),
.Y(n_524)
);

CKINVDCx16_ASAP7_75t_R g525 ( 
.A(n_461),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_465),
.B(n_464),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_464),
.B(n_458),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_461),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_493),
.Y(n_529)
);

NAND4xp25_ASAP7_75t_L g530 ( 
.A(n_477),
.B(n_485),
.C(n_489),
.D(n_484),
.Y(n_530)
);

OR2x6_ASAP7_75t_L g531 ( 
.A(n_476),
.B(n_455),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_493),
.Y(n_532)
);

AOI221xp5_ASAP7_75t_L g533 ( 
.A1(n_451),
.A2(n_478),
.B1(n_477),
.B2(n_452),
.C(n_460),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g534 ( 
.A(n_493),
.B(n_455),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_526),
.B(n_482),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_499),
.B(n_482),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_529),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_499),
.B(n_456),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_508),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_511),
.B(n_456),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_508),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_532),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_530),
.A2(n_452),
.B1(n_476),
.B2(n_469),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_512),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_512),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_510),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_483),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_527),
.B(n_467),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_501),
.B(n_502),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_505),
.B(n_490),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_506),
.B(n_490),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_514),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_514),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_509),
.B(n_533),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_497),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_516),
.B(n_490),
.Y(n_556)
);

INVx5_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_531),
.B(n_479),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_500),
.B(n_467),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_531),
.B(n_500),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_500),
.B(n_474),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_519),
.B(n_474),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_474),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_504),
.B(n_494),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_523),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_523),
.B(n_496),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_503),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_496),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_507),
.B(n_531),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_507),
.B(n_525),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_521),
.B(n_522),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_498),
.B(n_515),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_517),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_522),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_517),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_528),
.B(n_524),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_528),
.B(n_513),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_528),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_528),
.B(n_513),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_518),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_555),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_546),
.B(n_524),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_524),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_554),
.B(n_518),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_537),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_554),
.B(n_564),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_542),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_564),
.B(n_503),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_542),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_552),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_538),
.B(n_503),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_552),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_536),
.B(n_535),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_539),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_553),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_571),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_536),
.B(n_535),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_547),
.B(n_563),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_541),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_547),
.B(n_563),
.Y(n_603)
);

NOR2x1_ASAP7_75t_L g604 ( 
.A(n_548),
.B(n_570),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_549),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_540),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_549),
.B(n_568),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_540),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_565),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_572),
.B(n_560),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_560),
.B(n_559),
.Y(n_611)
);

AND2x4_ASAP7_75t_SL g612 ( 
.A(n_560),
.B(n_567),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_560),
.B(n_565),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_586),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_595),
.B(n_569),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_595),
.B(n_570),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_588),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_561),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_573),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_609),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_600),
.B(n_569),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g623 ( 
.A(n_602),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_600),
.B(n_544),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_582),
.B(n_587),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_588),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_589),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_606),
.B(n_544),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_589),
.B(n_591),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_591),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_599),
.B(n_558),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_596),
.B(n_575),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_601),
.B(n_545),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_585),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_606),
.B(n_545),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_592),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_592),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_610),
.B(n_581),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_611),
.B(n_575),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_599),
.B(n_573),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_594),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_594),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_597),
.B(n_558),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_613),
.B(n_543),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_590),
.B(n_583),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_615),
.B(n_601),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_617),
.B(n_608),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_615),
.B(n_603),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_629),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_634),
.A2(n_604),
.B1(n_603),
.B2(n_571),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_622),
.B(n_608),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_629),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_614),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_622),
.B(n_593),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_614),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_629),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_627),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_643),
.B(n_604),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_617),
.B(n_593),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_627),
.Y(n_660)
);

AOI32xp33_ASAP7_75t_L g661 ( 
.A1(n_645),
.A2(n_584),
.A3(n_550),
.B1(n_612),
.B2(n_577),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_621),
.Y(n_662)
);

O2A1O1Ixp33_ASAP7_75t_SL g663 ( 
.A1(n_662),
.A2(n_625),
.B(n_632),
.C(n_639),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_L g664 ( 
.A1(n_658),
.A2(n_644),
.B1(n_619),
.B2(n_620),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_649),
.B(n_643),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_662),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_651),
.B(n_631),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_650),
.B(n_638),
.Y(n_668)
);

NAND3x2_ASAP7_75t_L g669 ( 
.A(n_652),
.B(n_643),
.C(n_631),
.Y(n_669)
);

OAI322xp33_ASAP7_75t_L g670 ( 
.A1(n_650),
.A2(n_628),
.A3(n_635),
.B1(n_640),
.B2(n_618),
.C1(n_616),
.C2(n_626),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_660),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_653),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_651),
.B(n_631),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_653),
.Y(n_674)
);

O2A1O1Ixp5_ASAP7_75t_L g675 ( 
.A1(n_664),
.A2(n_656),
.B(n_655),
.C(n_657),
.Y(n_675)
);

OAI211xp5_ASAP7_75t_SL g676 ( 
.A1(n_663),
.A2(n_661),
.B(n_659),
.C(n_623),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_671),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_668),
.A2(n_669),
.B(n_666),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_665),
.A2(n_612),
.B1(n_658),
.B2(n_584),
.Y(n_679)
);

NAND2x1p5_ASAP7_75t_L g680 ( 
.A(n_665),
.B(n_635),
.Y(n_680)
);

AOI222xp33_ASAP7_75t_L g681 ( 
.A1(n_666),
.A2(n_624),
.B1(n_646),
.B2(n_648),
.C1(n_633),
.C2(n_654),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_667),
.B(n_647),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_678),
.B(n_673),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_680),
.B(n_658),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_677),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_676),
.A2(n_670),
.B1(n_672),
.B2(n_674),
.C(n_657),
.Y(n_686)
);

NOR3xp33_ASAP7_75t_L g687 ( 
.A(n_675),
.B(n_567),
.C(n_577),
.Y(n_687)
);

NAND3xp33_ASAP7_75t_L g688 ( 
.A(n_681),
.B(n_641),
.C(n_637),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_687),
.B(n_679),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_685),
.B(n_682),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_683),
.A2(n_628),
.B1(n_672),
.B2(n_637),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g692 ( 
.A(n_688),
.B(n_567),
.C(n_580),
.Y(n_692)
);

NOR3xp33_ASAP7_75t_L g693 ( 
.A(n_686),
.B(n_567),
.C(n_580),
.Y(n_693)
);

NAND4xp75_ASAP7_75t_L g694 ( 
.A(n_689),
.B(n_684),
.C(n_551),
.D(n_556),
.Y(n_694)
);

NAND3xp33_ASAP7_75t_L g695 ( 
.A(n_693),
.B(n_578),
.C(n_550),
.Y(n_695)
);

XNOR2x1_ASAP7_75t_SL g696 ( 
.A(n_692),
.B(n_551),
.Y(n_696)
);

NOR2x1_ASAP7_75t_L g697 ( 
.A(n_694),
.B(n_691),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_695),
.Y(n_698)
);

NOR3xp33_ASAP7_75t_L g699 ( 
.A(n_696),
.B(n_690),
.C(n_578),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_655),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_698),
.Y(n_701)
);

AOI22x1_ASAP7_75t_L g702 ( 
.A1(n_697),
.A2(n_556),
.B1(n_558),
.B2(n_576),
.Y(n_702)
);

NOR3xp33_ASAP7_75t_L g703 ( 
.A(n_699),
.B(n_700),
.C(n_579),
.Y(n_703)
);

AND2x2_ASAP7_75t_SL g704 ( 
.A(n_699),
.B(n_558),
.Y(n_704)
);

OAI22x1_ASAP7_75t_L g705 ( 
.A1(n_697),
.A2(n_557),
.B1(n_630),
.B2(n_642),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_698),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_701),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_706),
.B(n_624),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_702),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_705),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_703),
.B(n_704),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_707),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_708),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_711),
.A2(n_557),
.B(n_574),
.Y(n_714)
);

OAI321xp33_ASAP7_75t_L g715 ( 
.A1(n_710),
.A2(n_576),
.A3(n_574),
.B1(n_597),
.B2(n_598),
.C(n_630),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_714),
.A2(n_711),
.B(n_709),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_712),
.Y(n_717)
);

XOR2xp5_ASAP7_75t_L g718 ( 
.A(n_713),
.B(n_579),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_718),
.A2(n_715),
.B1(n_579),
.B2(n_636),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_642),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_717),
.A2(n_576),
.B(n_574),
.Y(n_721)
);

XNOR2xp5_ASAP7_75t_L g722 ( 
.A(n_720),
.B(n_633),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_722),
.B(n_721),
.Y(n_723)
);

OR2x6_ASAP7_75t_L g724 ( 
.A(n_723),
.B(n_719),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_724),
.A2(n_557),
.B(n_636),
.Y(n_725)
);


endmodule