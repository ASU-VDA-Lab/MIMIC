module fake_jpeg_10942_n_390 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_0),
.B(n_1),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_7),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_SL g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_57),
.Y(n_157)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_59),
.B(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_60),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_62),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_63),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_64),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_65),
.B(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_67),
.Y(n_165)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx2_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_17),
.B(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_72),
.B(n_86),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_26),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_74),
.B(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g130 ( 
.A(n_76),
.Y(n_130)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_9),
.Y(n_81)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g136 ( 
.A(n_82),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_17),
.B(n_30),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_24),
.B(n_9),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_18),
.B(n_4),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_88),
.B(n_96),
.Y(n_152)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g142 ( 
.A(n_92),
.Y(n_142)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

OR2x2_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_6),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g144 ( 
.A(n_95),
.B(n_34),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_13),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_14),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_99),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_19),
.A2(n_15),
.B(n_2),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_104),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_25),
.B(n_2),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

CKINVDCx12_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_106),
.Y(n_125)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_112),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_111),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_25),
.B(n_2),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_39),
.B(n_53),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_124),
.C(n_151),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_60),
.A2(n_46),
.B1(n_22),
.B2(n_31),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_120),
.A2(n_164),
.B1(n_166),
.B2(n_137),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_57),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_121),
.B(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_58),
.A2(n_42),
.B1(n_46),
.B2(n_53),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_123),
.A2(n_76),
.B1(n_100),
.B2(n_175),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_39),
.C(n_22),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_95),
.A2(n_34),
.B(n_27),
.C(n_30),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_139),
.B(n_145),
.Y(n_212)
);

OR2x2_ASAP7_75t_SL g229 ( 
.A(n_144),
.B(n_95),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_36),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_101),
.A2(n_31),
.B1(n_27),
.B2(n_36),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_159),
.B1(n_175),
.B2(n_114),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_71),
.B(n_51),
.Y(n_149)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_61),
.B(n_31),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_92),
.B(n_54),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_92),
.B(n_51),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_56),
.A2(n_32),
.B1(n_33),
.B2(n_43),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_69),
.B(n_32),
.C(n_33),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_119),
.C(n_125),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_84),
.B(n_43),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g211 ( 
.A(n_163),
.B(n_168),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_66),
.A2(n_52),
.B1(n_54),
.B2(n_48),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_67),
.A2(n_52),
.B1(n_48),
.B2(n_3),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_63),
.B(n_3),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_64),
.B(n_89),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_136),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_80),
.A2(n_3),
.B1(n_70),
.B2(n_57),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_177),
.Y(n_235)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_136),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_179),
.B(n_198),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_90),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_180),
.B(n_189),
.Y(n_237)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_108),
.B1(n_93),
.B2(n_103),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_183),
.A2(n_205),
.B1(n_209),
.B2(n_193),
.Y(n_261)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_186),
.A2(n_187),
.B1(n_197),
.B2(n_180),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_123),
.A2(n_159),
.B1(n_146),
.B2(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_190),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_134),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_195),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_127),
.A2(n_120),
.B1(n_151),
.B2(n_124),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_135),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_196),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_152),
.B(n_143),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_127),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_213),
.Y(n_260)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_161),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_202),
.Y(n_231)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_150),
.B1(n_170),
.B2(n_176),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_201),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_133),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_203),
.B(n_207),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_210),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_150),
.A2(n_118),
.B1(n_147),
.B2(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_208),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_118),
.A2(n_167),
.B1(n_173),
.B2(n_156),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_230),
.B(n_211),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_131),
.B(n_171),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_116),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_216),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_128),
.A2(n_130),
.B(n_157),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_201),
.C(n_217),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_170),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_222),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_140),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_229),
.B1(n_185),
.B2(n_195),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_147),
.B(n_165),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_220),
.Y(n_265)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_128),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_167),
.A2(n_138),
.B1(n_140),
.B2(n_156),
.Y(n_221)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_205),
.B1(n_203),
.B2(n_200),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_138),
.B(n_116),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_116),
.B(n_160),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_225),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_142),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_160),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_227),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_152),
.B(n_132),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_228),
.Y(n_243)
);

NOR2x1_ASAP7_75t_L g230 ( 
.A(n_134),
.B(n_122),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_232),
.A2(n_265),
.B(n_249),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_239),
.A2(n_261),
.B1(n_255),
.B2(n_237),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_247),
.B(n_220),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_252),
.A2(n_239),
.B1(n_231),
.B2(n_245),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_254),
.B(n_258),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_194),
.B(n_207),
.C(n_189),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_267),
.C(n_248),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_213),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_184),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_259),
.B(n_262),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_261),
.A2(n_181),
.B1(n_182),
.B2(n_190),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_198),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_270),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_191),
.B(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_268),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_230),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_188),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_187),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_260),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_252),
.A2(n_271),
.B1(n_234),
.B2(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_272),
.A2(n_285),
.B1(n_301),
.B2(n_242),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_232),
.A2(n_212),
.B(n_215),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_280),
.B(n_281),
.Y(n_303)
);

OA21x2_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_229),
.B(n_212),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_275),
.C(n_276),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_SL g275 ( 
.A(n_248),
.B(n_199),
.C(n_201),
.Y(n_275)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_234),
.B(n_201),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_268),
.B(n_178),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_279),
.B(n_263),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_256),
.A2(n_186),
.B(n_226),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_216),
.B(n_214),
.Y(n_281)
);

INVx13_ASAP7_75t_L g282 ( 
.A(n_250),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_288),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_283),
.A2(n_266),
.B1(n_238),
.B2(n_257),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_284),
.A2(n_287),
.B(n_292),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_262),
.A2(n_177),
.B1(n_206),
.B2(n_208),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_286),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_218),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_290),
.C(n_300),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_218),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_258),
.B(n_265),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_302),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_233),
.Y(n_296)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

NOR2x1_ASAP7_75t_L g298 ( 
.A(n_254),
.B(n_260),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_299),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_264),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_245),
.A2(n_243),
.B(n_241),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_253),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_311),
.C(n_315),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_302),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_291),
.B(n_270),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_286),
.Y(n_312)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_243),
.C(n_259),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_240),
.C(n_238),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_316),
.B(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_317),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_240),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_321),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_257),
.C(n_244),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_236),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_324),
.B(n_280),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_272),
.A2(n_242),
.B1(n_246),
.B2(n_269),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_305),
.Y(n_327)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_328),
.A2(n_298),
.B(n_283),
.Y(n_352)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_330),
.B(n_331),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_296),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_308),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_334),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_303),
.A2(n_301),
.B(n_277),
.C(n_281),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_SL g347 ( 
.A1(n_333),
.A2(n_322),
.B(n_303),
.C(n_275),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_299),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_324),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_336),
.A2(n_339),
.B1(n_341),
.B2(n_315),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_293),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_338),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_323),
.A2(n_292),
.B1(n_287),
.B2(n_273),
.Y(n_339)
);

OAI322xp33_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_294),
.A3(n_279),
.B1(n_295),
.B2(n_274),
.C1(n_298),
.C2(n_289),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_311),
.C(n_309),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_342),
.B(n_326),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_313),
.C(n_309),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_349),
.C(n_351),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_329),
.A2(n_314),
.B1(n_320),
.B2(n_287),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_328),
.Y(n_358)
);

OAI31xp33_ASAP7_75t_L g357 ( 
.A1(n_347),
.A2(n_348),
.A3(n_333),
.B(n_339),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_313),
.C(n_307),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_290),
.C(n_322),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_352),
.A2(n_326),
.B(n_333),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_285),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_334),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_350),
.A2(n_329),
.B1(n_336),
.B2(n_341),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_355),
.Y(n_368)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_353),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_356),
.A2(n_357),
.B(n_364),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_358),
.A2(n_359),
.B(n_363),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_365),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_331),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_362),
.B(n_342),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_344),
.A2(n_332),
.B1(n_340),
.B2(n_330),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_325),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_362),
.B(n_343),
.C(n_351),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_370),
.A2(n_235),
.B(n_246),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_361),
.B(n_345),
.C(n_347),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_361),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_359),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_SL g377 ( 
.A1(n_373),
.A2(n_365),
.B(n_347),
.Y(n_377)
);

AOI322xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_355),
.A3(n_357),
.B1(n_333),
.B2(n_358),
.C1(n_347),
.C2(n_346),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_378),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_379),
.B(n_371),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_377),
.A2(n_367),
.B(n_372),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_369),
.A2(n_333),
.B1(n_325),
.B2(n_360),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_376),
.B(n_368),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_380),
.B(n_382),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_381),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_383),
.B(n_366),
.C(n_370),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_384),
.B(n_371),
.C(n_288),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_385),
.A2(n_368),
.B(n_377),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_388),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_389),
.A2(n_386),
.B(n_288),
.Y(n_390)
);


endmodule