module fake_jpeg_8160_n_83 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_48;
wire n_46;
wire n_62;
wire n_43;
wire n_82;

INVx8_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_0),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g68 ( 
.A(n_54),
.B(n_59),
.Y(n_68)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_43),
.Y(n_56)
);

AO22x1_ASAP7_75t_L g63 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_3),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_52),
.B1(n_51),
.B2(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_42),
.B1(n_40),
.B2(n_8),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_47),
.Y(n_73)
);

NOR4xp25_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_4),
.C(n_7),
.D(n_9),
.Y(n_70)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_71),
.B1(n_73),
.B2(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_69),
.B1(n_64),
.B2(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_10),
.B(n_11),
.Y(n_78)
);

AOI322xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_17),
.C2(n_18),
.Y(n_79)
);

OAI31xp33_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_21),
.A3(n_22),
.B(n_25),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_80),
.A2(n_27),
.B(n_30),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_33),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_36),
.Y(n_83)
);


endmodule