module fake_jpeg_30224_n_348 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_348);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_348;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_3),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_53),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_26),
.B(n_1),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_39),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_40),
.B1(n_26),
.B2(n_31),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_65),
.A2(n_82),
.B1(n_92),
.B2(n_35),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_67),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_76),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_77),
.B(n_85),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_53),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_43),
.B(n_36),
.Y(n_85)
);

CKINVDCx12_ASAP7_75t_R g86 ( 
.A(n_48),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_40),
.B1(n_28),
.B2(n_33),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_87),
.A2(n_95),
.B1(n_24),
.B2(n_22),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_21),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_40),
.B1(n_28),
.B2(n_22),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_39),
.B(n_20),
.C(n_38),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_20),
.Y(n_103)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_52),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_105),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_73),
.A2(n_21),
.B(n_40),
.C(n_22),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_108),
.A2(n_79),
.B(n_63),
.C(n_97),
.Y(n_165)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_75),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_116),
.Y(n_145)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_30),
.B1(n_35),
.B2(n_33),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_140),
.B1(n_91),
.B2(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_119),
.B1(n_81),
.B2(n_80),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_69),
.A2(n_35),
.B1(n_28),
.B2(n_37),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_64),
.B(n_21),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_121),
.B(n_138),
.Y(n_177)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_122),
.A2(n_123),
.B(n_137),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_123)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_21),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_132),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_21),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_79),
.Y(n_159)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_33),
.B1(n_37),
.B2(n_32),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_75),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_71),
.A2(n_33),
.B1(n_21),
.B2(n_27),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_95),
.A2(n_27),
.B1(n_6),
.B2(n_7),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_106),
.B(n_27),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_147),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_108),
.A2(n_100),
.B(n_63),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_180),
.C(n_119),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_102),
.B1(n_125),
.B2(n_132),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_100),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_156),
.B(n_158),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_168),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

BUFx8_ASAP7_75t_L g207 ( 
.A(n_160),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_96),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_162),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_144),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_170),
.B1(n_117),
.B2(n_140),
.Y(n_184)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_91),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_178),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_97),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_130),
.Y(n_172)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_5),
.B(n_6),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_7),
.Y(n_182)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_131),
.B(n_5),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_107),
.B(n_6),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_179),
.B(n_8),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_128),
.A2(n_102),
.B(n_74),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_186),
.C(n_206),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_184),
.A2(n_195),
.B1(n_214),
.B2(n_151),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_134),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_202),
.B(n_148),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_118),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_196),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_149),
.A2(n_124),
.B1(n_114),
.B2(n_143),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_194),
.A2(n_197),
.B(n_209),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_127),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_163),
.A2(n_125),
.B1(n_124),
.B2(n_111),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_114),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_201),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_145),
.B(n_112),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_111),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_205),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_144),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_158),
.B(n_8),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_10),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_135),
.C(n_81),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_146),
.C(n_174),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_212),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_165),
.A2(n_80),
.B1(n_98),
.B2(n_11),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_9),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_11),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_159),
.A2(n_149),
.B1(n_165),
.B2(n_163),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_176),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_216),
.B(n_218),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_208),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_223),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_185),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_226),
.Y(n_251)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_227),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_228),
.B(n_232),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_230),
.A2(n_234),
.B(n_211),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_190),
.B(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_171),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_191),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_198),
.B(n_175),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_186),
.B(n_12),
.Y(n_235)
);

AOI221xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_242),
.B1(n_243),
.B2(n_209),
.C(n_203),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_237),
.A2(n_183),
.B1(n_207),
.B2(n_15),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_241),
.C(n_183),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_181),
.B1(n_174),
.B2(n_166),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_146),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_196),
.B(n_15),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_182),
.A2(n_153),
.B(n_157),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_214),
.A2(n_157),
.B(n_164),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_244),
.A2(n_210),
.B(n_194),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_236),
.B(n_222),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_202),
.B1(n_229),
.B2(n_237),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_247),
.A2(n_257),
.B1(n_222),
.B2(n_225),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_248),
.B(n_261),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_192),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_253),
.C(n_259),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_184),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_202),
.B1(n_195),
.B2(n_204),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_258),
.A2(n_242),
.B1(n_226),
.B2(n_235),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_193),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_204),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_234),
.Y(n_273)
);

AOI221xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_181),
.B1(n_188),
.B2(n_153),
.C(n_164),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_239),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_223),
.B1(n_216),
.B2(n_221),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_252),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_274),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_240),
.B(n_217),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_269),
.A2(n_277),
.B(n_284),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_270),
.A2(n_259),
.B(n_225),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_275),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_246),
.A2(n_217),
.B(n_236),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_278),
.B(n_279),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_249),
.B(n_221),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_280),
.A2(n_285),
.B1(n_264),
.B2(n_253),
.Y(n_301)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_218),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_282),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_232),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_283),
.Y(n_302)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_262),
.B(n_219),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_272),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_296),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_266),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_293),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_261),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_264),
.Y(n_294)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_245),
.C(n_250),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_301),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_280),
.B1(n_270),
.B2(n_273),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_298),
.A2(n_273),
.B(n_281),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_305),
.A2(n_314),
.B(n_299),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_310),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_288),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_295),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_311),
.B(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_299),
.A2(n_277),
.B(n_269),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_276),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_318),
.Y(n_329)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_317),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_289),
.B(n_300),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_297),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_320),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_293),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_288),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_324),
.C(n_306),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

AOI21xp33_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_304),
.B(n_289),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_312),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_323),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_296),
.C(n_307),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_308),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_308),
.C(n_315),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_247),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_323),
.C(n_301),
.Y(n_337)
);

INVx11_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_254),
.C(n_257),
.Y(n_339)
);

AOI31xp67_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_329),
.A3(n_326),
.B(n_330),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_215),
.Y(n_344)
);

OAI311xp33_ASAP7_75t_L g343 ( 
.A1(n_341),
.A2(n_336),
.A3(n_334),
.B1(n_284),
.C1(n_248),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_343),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_344),
.C(n_342),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_254),
.B(n_227),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_224),
.Y(n_348)
);


endmodule