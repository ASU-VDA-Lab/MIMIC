module fake_jpeg_15700_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_19),
.B1(n_23),
.B2(n_31),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_29),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_17),
.B1(n_30),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_29),
.B1(n_18),
.B2(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_82),
.B1(n_48),
.B2(n_45),
.Y(n_94)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_61),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_36),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_0),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_76),
.B(n_0),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_37),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_45),
.B1(n_55),
.B2(n_50),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_44),
.B1(n_55),
.B2(n_50),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_23),
.B1(n_30),
.B2(n_17),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_70),
.A2(n_55),
.B1(n_56),
.B2(n_25),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_21),
.B1(n_30),
.B2(n_34),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_13),
.B1(n_12),
.B2(n_48),
.Y(n_96)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_35),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_26),
.B(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_50),
.B(n_12),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_13),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_37),
.B1(n_35),
.B2(n_26),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_32),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_40),
.B(n_12),
.C(n_13),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_86),
.B(n_93),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_105),
.Y(n_134)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_92),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_99),
.B1(n_101),
.B2(n_113),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_32),
.C(n_39),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_61),
.C(n_74),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_100),
.B1(n_114),
.B2(n_56),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

CKINVDCx12_ASAP7_75t_R g105 ( 
.A(n_59),
.Y(n_105)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

CKINVDCx9p33_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_62),
.A2(n_56),
.B1(n_25),
.B2(n_22),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_109),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_115),
.B(n_110),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_111),
.C(n_108),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_22),
.Y(n_158)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_87),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_22),
.B(n_20),
.Y(n_154)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_104),
.A2(n_63),
.B1(n_65),
.B2(n_75),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_129),
.B1(n_132),
.B2(n_135),
.Y(n_167)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_63),
.B1(n_65),
.B2(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_114),
.A2(n_77),
.B1(n_57),
.B2(n_79),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_88),
.A2(n_57),
.B1(n_77),
.B2(n_78),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_85),
.B1(n_84),
.B2(n_53),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_108),
.B1(n_97),
.B2(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_99),
.A2(n_54),
.B1(n_2),
.B2(n_3),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_86),
.A2(n_1),
.B(n_2),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_139),
.B(n_1),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_98),
.B(n_39),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_96),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_142),
.B(n_20),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_144),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_145),
.A2(n_153),
.B1(n_119),
.B2(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_120),
.B(n_93),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_146),
.B(n_156),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_150),
.C(n_162),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_107),
.B1(n_102),
.B2(n_112),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_152),
.B(n_117),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_109),
.C(n_89),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_105),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_151),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_136),
.A2(n_89),
.B(n_16),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_110),
.B1(n_102),
.B2(n_54),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_169),
.B(n_20),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_92),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_89),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_129),
.B(n_83),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_1),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_134),
.B(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_173),
.A2(n_175),
.B(n_183),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_147),
.C(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_181),
.C(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_191),
.Y(n_210)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_134),
.B(n_139),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_193),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_89),
.C(n_135),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g183 ( 
.A(n_141),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_119),
.Y(n_184)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_187),
.A2(n_197),
.B(n_199),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_167),
.B1(n_166),
.B2(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_194),
.B1(n_198),
.B2(n_22),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_145),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_137),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_166),
.A2(n_128),
.B1(n_137),
.B2(n_92),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_153),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_106),
.B1(n_66),
.B2(n_20),
.Y(n_198)
);

AOI32xp33_ASAP7_75t_L g199 ( 
.A1(n_152),
.A2(n_92),
.A3(n_16),
.B1(n_28),
.B2(n_27),
.Y(n_199)
);

XOR2x1_ASAP7_75t_L g200 ( 
.A(n_142),
.B(n_169),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_27),
.B(n_24),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_28),
.B(n_27),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_159),
.B(n_157),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_220),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_213),
.C(n_214),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_200),
.B(n_171),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_223),
.C(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_217),
.B(n_192),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_177),
.B(n_201),
.Y(n_212)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_212),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_143),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_143),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_140),
.B1(n_149),
.B2(n_155),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_215),
.A2(n_226),
.B1(n_228),
.B2(n_203),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_221),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_187),
.A2(n_140),
.B(n_155),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_25),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_218),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_28),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_186),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_222),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_106),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_224),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_185),
.B1(n_184),
.B2(n_173),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_106),
.B1(n_54),
.B2(n_4),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_24),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_172),
.Y(n_243)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_234),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_SL g234 ( 
.A1(n_217),
.A2(n_175),
.B(n_188),
.C(n_182),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_203),
.B(n_188),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_243),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_190),
.B1(n_178),
.B2(n_195),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_237),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_209),
.A2(n_178),
.B(n_179),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

NOR2x1_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_227),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_218),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_24),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_2),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_54),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_213),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_256),
.C(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_207),
.C(n_214),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_226),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_243),
.C(n_245),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_204),
.C(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_264),
.C(n_222),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_223),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_229),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_215),
.C(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_267),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_238),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_268),
.B(n_232),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_259),
.A2(n_240),
.B(n_234),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_270),
.B(n_275),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_272),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_249),
.C(n_231),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_247),
.B1(n_236),
.B2(n_232),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_280),
.B1(n_281),
.B2(n_263),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_211),
.B(n_234),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_234),
.B(n_211),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_266),
.B1(n_264),
.B2(n_253),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_256),
.B1(n_260),
.B2(n_254),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_262),
.A2(n_228),
.B1(n_3),
.B2(n_4),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_2),
.B(n_3),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_5),
.C(n_6),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_251),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_283),
.B(n_5),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_274),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_286),
.B(n_287),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_288),
.B(n_291),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_5),
.CI(n_6),
.CON(n_290),
.SN(n_290)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_292),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_5),
.C(n_6),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_277),
.C(n_282),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_272),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_269),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_298),
.C(n_303),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_284),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_269),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_271),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_293),
.C(n_275),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_285),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_307),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_281),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_311),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_293),
.B1(n_292),
.B2(n_290),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_300),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_298),
.B(n_303),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_313),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_317),
.A2(n_315),
.B(n_312),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_305),
.A3(n_306),
.B1(n_287),
.B2(n_278),
.C1(n_11),
.C2(n_10),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_7),
.B(n_8),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_7),
.C(n_8),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_11),
.C(n_8),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_10),
.Y(n_323)
);


endmodule