module fake_jpeg_11498_n_644 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_12),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_65),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_66),
.Y(n_175)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_67),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_69),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_70),
.B(n_86),
.Y(n_137)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_72),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_73),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_74),
.Y(n_214)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_76),
.Y(n_215)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_81),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_82),
.Y(n_199)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g156 ( 
.A(n_85),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_18),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_89),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_18),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_37),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_98),
.Y(n_166)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_95),
.Y(n_183)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_27),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_16),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_99),
.B(n_106),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_101),
.Y(n_202)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_56),
.B(n_14),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_35),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_50),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_54),
.B1(n_22),
.B2(n_40),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_35),
.Y(n_115)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_56),
.B(n_14),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_117),
.B(n_118),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g118 ( 
.A(n_28),
.Y(n_118)
);

CKINVDCx9p33_ASAP7_75t_R g119 ( 
.A(n_48),
.Y(n_119)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_48),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_121),
.B(n_124),
.Y(n_197)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_123),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_53),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_28),
.Y(n_125)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_39),
.Y(n_126)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_39),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g194 ( 
.A(n_127),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_54),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_128),
.B(n_31),
.Y(n_208)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_129),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_130),
.A2(n_164),
.B1(n_13),
.B2(n_11),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_62),
.B(n_22),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_139),
.B(n_151),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

CKINVDCx11_ASAP7_75t_R g158 ( 
.A(n_85),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_158),
.B(n_160),
.Y(n_243)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx11_ASAP7_75t_L g266 ( 
.A(n_159),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_62),
.B(n_24),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_61),
.B1(n_109),
.B2(n_110),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_65),
.A2(n_51),
.B1(n_39),
.B2(n_45),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_169),
.A2(n_84),
.B1(n_80),
.B2(n_41),
.Y(n_236)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

NAND2x1_ASAP7_75t_L g174 ( 
.A(n_67),
.B(n_58),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_174),
.B(n_13),
.C(n_134),
.Y(n_276)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_176),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_24),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_177),
.B(n_180),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_116),
.B(n_58),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_40),
.Y(n_180)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_68),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_198),
.Y(n_291)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_201),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_68),
.Y(n_205)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_60),
.Y(n_207)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_64),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g247 ( 
.A(n_209),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_90),
.B(n_31),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_210),
.B(n_212),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_66),
.B(n_26),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_69),
.B(n_26),
.Y(n_216)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_208),
.C(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_72),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_2),
.Y(n_250)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

INVx11_ASAP7_75t_L g220 ( 
.A(n_74),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_221),
.Y(n_297)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_227),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_147),
.A2(n_114),
.B1(n_108),
.B2(n_107),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_228),
.A2(n_232),
.B1(n_254),
.B2(n_270),
.Y(n_321)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_149),
.Y(n_229)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_229),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_45),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_231),
.B(n_239),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_130),
.A2(n_105),
.B1(n_104),
.B2(n_100),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_233),
.B(n_242),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_236),
.A2(n_237),
.B1(n_260),
.B2(n_269),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_141),
.A2(n_41),
.B1(n_34),
.B2(n_3),
.Y(n_237)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_238),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_34),
.Y(n_239)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_137),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_136),
.Y(n_244)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_244),
.Y(n_343)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

INVx6_ASAP7_75t_SL g246 ( 
.A(n_156),
.Y(n_246)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_246),
.Y(n_317)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_196),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_248),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_166),
.B(n_1),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_249),
.B(n_255),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_250),
.Y(n_349)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_252),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_179),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_253),
.A2(n_272),
.B(n_161),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_169),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_166),
.B(n_135),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_148),
.Y(n_256)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_138),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_258),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_187),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_152),
.B(n_10),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_261),
.B(n_271),
.Y(n_356)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_168),
.Y(n_262)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_262),
.Y(n_332)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_150),
.Y(n_264)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_264),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_265),
.A2(n_287),
.B1(n_184),
.B2(n_195),
.Y(n_331)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_150),
.Y(n_267)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

CKINVDCx12_ASAP7_75t_R g268 ( 
.A(n_156),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_268),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_187),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_164),
.A2(n_11),
.B1(n_13),
.B2(n_212),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_153),
.B(n_157),
.Y(n_271)
);

NAND2xp33_ASAP7_75t_SL g272 ( 
.A(n_174),
.B(n_11),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_183),
.Y(n_274)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_274),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_175),
.Y(n_275)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_275),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_288),
.Y(n_301)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_142),
.Y(n_277)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_277),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_190),
.B(n_137),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_279),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_134),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_280),
.Y(n_346)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_138),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_204),
.A2(n_173),
.B1(n_145),
.B2(n_131),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_285),
.B1(n_237),
.B2(n_260),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_190),
.B(n_216),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_286),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g285 ( 
.A1(n_146),
.A2(n_191),
.B1(n_185),
.B2(n_203),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_210),
.B(n_140),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_211),
.A2(n_162),
.B1(n_197),
.B2(n_155),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_197),
.B(n_218),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_167),
.Y(n_289)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

BUFx4f_ASAP7_75t_SL g290 ( 
.A(n_178),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_290),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_170),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_295),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_161),
.Y(n_293)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_293),
.Y(n_347)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_154),
.Y(n_294)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_132),
.B(n_133),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_186),
.B(n_202),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_298),
.Y(n_313)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_143),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_236),
.A2(n_204),
.B1(n_143),
.B2(n_193),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_302),
.A2(n_266),
.B1(n_247),
.B2(n_258),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_193),
.C(n_214),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g366 ( 
.A(n_306),
.B(n_309),
.CI(n_326),
.CON(n_366),
.SN(n_366)
);

MAJx2_ASAP7_75t_L g309 ( 
.A(n_223),
.B(n_144),
.C(n_199),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_318),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_320),
.B(n_269),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_226),
.B(n_273),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_324),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_171),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_206),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_325),
.B(n_338),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_276),
.B(n_175),
.C(n_184),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_331),
.A2(n_282),
.B1(n_294),
.B2(n_281),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_250),
.B(n_192),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_334),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_225),
.A2(n_195),
.B(n_214),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_270),
.B(n_213),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_243),
.B(n_192),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_339),
.B(n_348),
.Y(n_390)
);

OA22x2_ASAP7_75t_L g341 ( 
.A1(n_254),
.A2(n_215),
.B1(n_285),
.B2(n_266),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_341),
.B(n_267),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_224),
.B(n_215),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_351),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_263),
.B(n_234),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_291),
.B(n_259),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_350),
.B(n_290),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_253),
.B(n_235),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_251),
.B(n_297),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_357),
.B(n_252),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_359),
.A2(n_329),
.B1(n_310),
.B2(n_354),
.Y(n_441)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_361),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_362),
.A2(n_337),
.B(n_333),
.Y(n_408)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_300),
.B(n_246),
.Y(n_363)
);

AOI21xp33_ASAP7_75t_L g409 ( 
.A1(n_363),
.A2(n_396),
.B(n_334),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_291),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_364),
.B(n_380),
.Y(n_442)
);

INVx13_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_365),
.Y(n_439)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_304),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_367),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_368),
.A2(n_388),
.B1(n_400),
.B2(n_340),
.Y(n_417)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_369),
.Y(n_434)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_344),
.Y(n_370)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_357),
.Y(n_372)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_338),
.A2(n_284),
.B1(n_247),
.B2(n_299),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_374),
.A2(n_395),
.B1(n_352),
.B2(n_358),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_376),
.A2(n_342),
.B1(n_310),
.B2(n_354),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_325),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_377),
.B(n_378),
.Y(n_438)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_319),
.Y(n_379)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_308),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_345),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_384),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_324),
.A2(n_259),
.B(n_290),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_382),
.A2(n_358),
.B(n_353),
.Y(n_416)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_345),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_385),
.B(n_389),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_301),
.B(n_248),
.Y(n_386)
);

NAND2x1_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_397),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_312),
.B(n_230),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_321),
.A2(n_264),
.B1(n_244),
.B2(n_275),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_392),
.Y(n_423)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_393),
.B(n_394),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_322),
.B(n_240),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_321),
.A2(n_227),
.B1(n_238),
.B2(n_256),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_320),
.Y(n_396)
);

INVx13_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_327),
.B(n_277),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_398),
.B(n_402),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_301),
.B(n_333),
.Y(n_399)
);

OAI21xp33_ASAP7_75t_L g413 ( 
.A1(n_399),
.A2(n_401),
.B(n_336),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_331),
.A2(n_222),
.B1(n_293),
.B2(n_245),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_301),
.B(n_229),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_222),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_313),
.B(n_222),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_404),
.B(n_405),
.Y(n_431)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_335),
.Y(n_405)
);

NOR4xp25_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_349),
.C(n_309),
.D(n_351),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_SL g447 ( 
.A(n_406),
.B(n_383),
.C(n_394),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_407),
.B(n_413),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_408),
.A2(n_428),
.B(n_401),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_409),
.B(n_366),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_326),
.C(n_306),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_415),
.C(n_425),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_362),
.A2(n_349),
.B(n_352),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_420),
.B(n_360),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_386),
.C(n_401),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_416),
.A2(n_430),
.B(n_376),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_417),
.B(n_368),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_403),
.A2(n_341),
.B1(n_353),
.B2(n_328),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_418),
.A2(n_419),
.B1(n_427),
.B2(n_359),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_403),
.A2(n_341),
.B1(n_328),
.B2(n_305),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_362),
.A2(n_341),
.B(n_347),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_371),
.A2(n_305),
.B1(n_355),
.B2(n_330),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_421),
.A2(n_441),
.B1(n_400),
.B2(n_392),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_346),
.C(n_347),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_388),
.A2(n_355),
.B1(n_330),
.B2(n_343),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_382),
.A2(n_371),
.B(n_360),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_383),
.B(n_311),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_410),
.C(n_377),
.Y(n_456)
);

OAI32xp33_ASAP7_75t_L g440 ( 
.A1(n_375),
.A2(n_342),
.A3(n_311),
.B1(n_343),
.B2(n_316),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_376),
.Y(n_450)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_443),
.Y(n_445)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_445),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_446),
.A2(n_451),
.B(n_416),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_447),
.B(n_409),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_431),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_449),
.B(n_473),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_450),
.A2(n_478),
.B1(n_479),
.B2(n_426),
.Y(n_511)
);

AO21x1_ASAP7_75t_L g452 ( 
.A1(n_428),
.A2(n_360),
.B(n_375),
.Y(n_452)
);

AO22x1_ASAP7_75t_L g482 ( 
.A1(n_452),
.A2(n_406),
.B1(n_411),
.B2(n_414),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_390),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_453),
.B(n_468),
.Y(n_492)
);

BUFx8_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_454),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_455),
.A2(n_408),
.B(n_422),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_412),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_423),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_457),
.B(n_465),
.Y(n_494)
);

INVx13_ASAP7_75t_L g458 ( 
.A(n_435),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_460),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_419),
.A2(n_395),
.B1(n_370),
.B2(n_372),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_461),
.A2(n_414),
.B1(n_411),
.B2(n_441),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_462),
.A2(n_474),
.B1(n_407),
.B2(n_421),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_366),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_463),
.B(n_422),
.C(n_389),
.Y(n_507)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_464),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_423),
.Y(n_465)
);

INVx13_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_466),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_444),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_467),
.B(n_472),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_378),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_433),
.Y(n_469)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_469),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_424),
.B(n_393),
.Y(n_470)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_470),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_475),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_438),
.B(n_384),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_329),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_432),
.B(n_391),
.Y(n_475)
);

INVx13_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_476),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_424),
.B(n_381),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_434),
.Y(n_506)
);

INVx3_ASAP7_75t_SL g479 ( 
.A(n_434),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_456),
.B(n_415),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_480),
.B(n_486),
.C(n_489),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_374),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_485),
.A2(n_496),
.B1(n_478),
.B2(n_460),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_438),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_477),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_488),
.B(n_467),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_490),
.A2(n_502),
.B(n_446),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_448),
.B(n_366),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_497),
.C(n_500),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_448),
.B(n_431),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_498),
.B(n_507),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_452),
.B(n_425),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_502),
.A2(n_451),
.B(n_459),
.Y(n_525)
);

AO22x1_ASAP7_75t_L g505 ( 
.A1(n_455),
.A2(n_420),
.B1(n_436),
.B2(n_440),
.Y(n_505)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_506),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_L g508 ( 
.A1(n_450),
.A2(n_418),
.B1(n_417),
.B2(n_430),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_511),
.B1(n_461),
.B2(n_462),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_452),
.B(n_422),
.C(n_433),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_422),
.C(n_445),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_471),
.B(n_363),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_513),
.B(n_447),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_514),
.A2(n_525),
.B(n_535),
.Y(n_564)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_515),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_516),
.A2(n_541),
.B(n_482),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_518),
.A2(n_505),
.B1(n_504),
.B2(n_503),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_494),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_520),
.B(n_527),
.Y(n_549)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_483),
.Y(n_521)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_521),
.Y(n_556)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_522),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_508),
.A2(n_474),
.B1(n_459),
.B2(n_457),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_526),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_494),
.A2(n_474),
.B1(n_459),
.B2(n_465),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_492),
.B(n_495),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_532),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_533),
.Y(n_547)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_493),
.Y(n_530)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_530),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_481),
.B(n_464),
.Y(n_531)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_531),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_510),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_484),
.B(n_472),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_499),
.B(n_449),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_534),
.B(n_487),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_490),
.A2(n_470),
.B(n_426),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_SL g566 ( 
.A(n_536),
.B(n_427),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_480),
.B(n_469),
.C(n_479),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_537),
.B(n_500),
.C(n_507),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_497),
.B(n_405),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_539),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_385),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_540),
.A2(n_379),
.B1(n_476),
.B2(n_466),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_501),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_509),
.A2(n_479),
.B(n_466),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_496),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_545),
.B(n_524),
.C(n_519),
.Y(n_580)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_548),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_491),
.C(n_489),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_551),
.B(n_561),
.Y(n_571)
);

XNOR2x1_ASAP7_75t_L g579 ( 
.A(n_553),
.B(n_559),
.Y(n_579)
);

INVx5_ASAP7_75t_L g554 ( 
.A(n_516),
.Y(n_554)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_554),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_486),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_555),
.B(n_527),
.Y(n_583)
);

FAx1_ASAP7_75t_SL g557 ( 
.A(n_524),
.B(n_498),
.CI(n_513),
.CON(n_557),
.SN(n_557)
);

FAx1_ASAP7_75t_SL g585 ( 
.A(n_557),
.B(n_551),
.CI(n_545),
.CON(n_585),
.SN(n_585)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_523),
.B(n_487),
.C(n_429),
.Y(n_561)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_562),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_523),
.B(n_316),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_566),
.Y(n_568)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_567),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_544),
.A2(n_518),
.B1(n_517),
.B2(n_540),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_570),
.A2(n_552),
.B1(n_559),
.B2(n_531),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_542),
.Y(n_572)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_572),
.Y(n_589)
);

OAI22x1_ASAP7_75t_L g573 ( 
.A1(n_563),
.A2(n_526),
.B1(n_515),
.B2(n_517),
.Y(n_573)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_573),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_547),
.B(n_519),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g595 ( 
.A(n_576),
.B(n_583),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_R g577 ( 
.A(n_564),
.B(n_535),
.C(n_514),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_577),
.A2(n_560),
.B1(n_476),
.B2(n_458),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_580),
.B(n_581),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_557),
.A2(n_561),
.B(n_558),
.Y(n_581)
);

INVx13_ASAP7_75t_L g582 ( 
.A(n_562),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_582),
.B(n_549),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_546),
.B(n_543),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_584),
.B(n_550),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_585),
.B(n_586),
.Y(n_599)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_556),
.Y(n_586)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_587),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_571),
.B(n_565),
.C(n_547),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_588),
.B(n_593),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_591),
.B(n_592),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_569),
.B(n_543),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_555),
.C(n_553),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_541),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_598),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_572),
.A2(n_552),
.B1(n_557),
.B2(n_525),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_596),
.B(n_600),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_580),
.B(n_566),
.C(n_536),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_575),
.B(n_534),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_601),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_578),
.A2(n_533),
.B1(n_530),
.B2(n_521),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_602),
.A2(n_603),
.B1(n_570),
.B2(n_574),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_608),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_597),
.A2(n_585),
.B(n_577),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_SL g618 ( 
.A1(n_607),
.A2(n_612),
.B(n_596),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_588),
.B(n_593),
.C(n_600),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_595),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_609),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_590),
.B(n_585),
.C(n_579),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_611),
.B(n_613),
.Y(n_625)
);

AO21x1_ASAP7_75t_L g612 ( 
.A1(n_589),
.A2(n_573),
.B(n_579),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_576),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_610),
.B(n_602),
.Y(n_617)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_617),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_618),
.A2(n_626),
.B(n_458),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_614),
.B(n_595),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_619),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_616),
.C(n_609),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_620),
.A2(n_622),
.B(n_624),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_615),
.B(n_568),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_612),
.B(n_568),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_605),
.B(n_603),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_617),
.A2(n_604),
.B1(n_611),
.B2(n_582),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_633),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_629),
.A2(n_630),
.B(n_633),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_625),
.A2(n_621),
.B(n_623),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g633 ( 
.A(n_626),
.B(n_454),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_631),
.B(n_454),
.C(n_369),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_635),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_SL g639 ( 
.A1(n_636),
.A2(n_637),
.B(n_628),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_632),
.A2(n_454),
.B(n_369),
.Y(n_637)
);

OAI31xp33_ASAP7_75t_SL g640 ( 
.A1(n_639),
.A2(n_634),
.A3(n_365),
.B(n_361),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_640),
.B(n_361),
.C(n_365),
.Y(n_641)
);

OAI31xp33_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_638),
.A3(n_367),
.B(n_373),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_642),
.B(n_367),
.Y(n_643)
);

AO21x1_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_397),
.B(n_640),
.Y(n_644)
);


endmodule