module fake_jpeg_25712_n_228 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_15),
.B1(n_19),
.B2(n_45),
.Y(n_62)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_27),
.Y(n_45)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_60),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_18),
.B1(n_24),
.B2(n_22),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_33),
.B(n_32),
.C(n_31),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_62),
.B1(n_42),
.B2(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_64),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_18),
.B1(n_24),
.B2(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_15),
.B1(n_33),
.B2(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_63),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_43),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_64),
.A2(n_13),
.B(n_47),
.Y(n_66)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_74),
.B(n_30),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_68),
.A2(n_79),
.B1(n_82),
.B2(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_61),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_72),
.Y(n_84)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_41),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_41),
.C(n_47),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_53),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_30),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_74),
.B(n_73),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_20),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_15),
.B1(n_39),
.B2(n_25),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_39),
.B1(n_15),
.B2(n_19),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_71),
.B1(n_75),
.B2(n_81),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_77),
.C(n_81),
.Y(n_110)
);

NAND2x1_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_87),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_55),
.B1(n_54),
.B2(n_50),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_99),
.B1(n_68),
.B2(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_90),
.Y(n_102)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_94),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_69),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_59),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_19),
.B(n_1),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_98),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_59),
.B1(n_48),
.B2(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_109),
.B1(n_85),
.B2(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_67),
.B1(n_65),
.B2(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_90),
.Y(n_122)
);

NOR4xp25_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_65),
.C(n_75),
.D(n_49),
.Y(n_106)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_98),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_88),
.A2(n_75),
.B1(n_48),
.B2(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_116),
.B1(n_57),
.B2(n_19),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_117),
.C(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx6_ASAP7_75t_SL g115 ( 
.A(n_83),
.Y(n_115)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_71),
.B1(n_57),
.B2(n_19),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_40),
.C(n_57),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_86),
.B(n_95),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_132),
.B(n_13),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_87),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_135),
.B(n_20),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_117),
.C(n_101),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_121),
.C(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_134),
.B1(n_13),
.B2(n_25),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_87),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_83),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_83),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_128),
.B(n_111),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_144),
.Y(n_169)
);

AOI21x1_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_118),
.B(n_101),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_151),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_108),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_147),
.C(n_120),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_146),
.A2(n_154),
.B1(n_20),
.B2(n_25),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_115),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_150),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_129),
.B(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_13),
.B(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_119),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_14),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_148),
.A2(n_126),
.B1(n_123),
.B2(n_130),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_156),
.A2(n_166),
.B1(n_0),
.B2(n_1),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_155),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_157),
.A2(n_141),
.B(n_149),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_135),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_161),
.C(n_165),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_160),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_141),
.B(n_119),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_138),
.A2(n_134),
.B1(n_127),
.B2(n_120),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_167),
.B1(n_146),
.B2(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_127),
.C(n_40),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_14),
.B1(n_21),
.B2(n_16),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_21),
.B1(n_16),
.B2(n_14),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

OAI321xp33_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_171),
.A3(n_159),
.B1(n_158),
.B2(n_169),
.C(n_5),
.Y(n_187)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_182),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_170),
.A2(n_150),
.B1(n_144),
.B2(n_145),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_176),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_17),
.B(n_40),
.C(n_21),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_0),
.B(n_1),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_21),
.B1(n_16),
.B2(n_8),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_180),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_17),
.C(n_7),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_0),
.C(n_3),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_193),
.B(n_12),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_8),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_202),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_177),
.C(n_176),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_178),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_204),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_189),
.A2(n_183),
.B(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_196),
.A2(n_174),
.B1(n_178),
.B2(n_5),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_178),
.A3(n_3),
.B1(n_6),
.B2(n_9),
.C1(n_4),
.C2(n_11),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_213),
.Y(n_214)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_4),
.C(n_10),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_210),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_10),
.B(n_11),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_198),
.B(n_201),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_12),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_17),
.C(n_12),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_3),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_17),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

O2A1O1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_217),
.A2(n_17),
.B(n_216),
.C(n_219),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_222),
.A2(n_223),
.B(n_17),
.C(n_220),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_17),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_17),
.B(n_225),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_17),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_17),
.Y(n_228)
);


endmodule