module real_aes_8311_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_449;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g335 ( .A(n_0), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_1), .A2(n_81), .B1(n_175), .B2(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_1), .Y(n_529) );
AOI21xp33_ASAP7_75t_L g296 ( .A1(n_2), .A2(n_219), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g204 ( .A(n_3), .Y(n_204) );
AND2x6_ASAP7_75t_L g224 ( .A(n_3), .B(n_202), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_3), .B(n_520), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_4), .A2(n_218), .B(n_225), .Y(n_217) );
INVx1_ASAP7_75t_L g527 ( .A(n_4), .Y(n_527) );
INVx1_ASAP7_75t_L g302 ( .A(n_5), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_6), .B(n_283), .Y(n_282) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_7), .A2(n_21), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g216 ( .A(n_8), .Y(n_216) );
INVx1_ASAP7_75t_L g235 ( .A(n_9), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_10), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_11), .B(n_252), .Y(n_268) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_12), .A2(n_23), .B1(n_90), .B2(n_94), .Y(n_93) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_13), .B(n_219), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_14), .B(n_295), .Y(n_325) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_15), .A2(n_232), .B(n_234), .C(n_236), .Y(n_231) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_16), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_17), .B(n_267), .Y(n_336) );
INVx1_ASAP7_75t_L g314 ( .A(n_18), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g167 ( .A1(n_19), .A2(n_26), .B1(n_168), .B2(n_171), .Y(n_167) );
INVx2_ASAP7_75t_L g222 ( .A(n_20), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g106 ( .A1(n_22), .A2(n_45), .B1(n_107), .B2(n_113), .Y(n_106) );
OAI221xp5_ASAP7_75t_L g195 ( .A1(n_23), .A2(n_38), .B1(n_48), .B2(n_196), .C(n_197), .Y(n_195) );
INVxp67_ASAP7_75t_L g198 ( .A(n_23), .Y(n_198) );
OAI22xp5_ASAP7_75t_SL g187 ( .A1(n_24), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_187) );
INVxp67_ASAP7_75t_L g190 ( .A(n_24), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_25), .A2(n_224), .B(n_228), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g312 ( .A(n_27), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_28), .B(n_267), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_29), .Y(n_100) );
AOI22xp33_ASAP7_75t_L g160 ( .A1(n_30), .A2(n_51), .B1(n_161), .B2(n_164), .Y(n_160) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_31), .A2(n_55), .B1(n_180), .B2(n_181), .Y(n_179) );
INVxp67_ASAP7_75t_L g181 ( .A(n_31), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g315 ( .A(n_32), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_33), .B(n_219), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_34), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_35), .A2(n_228), .B1(n_309), .B2(n_311), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_36), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g332 ( .A(n_37), .Y(n_332) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_38), .A2(n_57), .B1(n_90), .B2(n_94), .Y(n_99) );
INVxp67_ASAP7_75t_L g199 ( .A(n_38), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_39), .A2(n_300), .B(n_301), .C(n_303), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_40), .Y(n_271) );
INVx1_ASAP7_75t_L g298 ( .A(n_41), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_42), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_43), .A2(n_58), .B1(n_152), .B2(n_156), .Y(n_151) );
INVx1_ASAP7_75t_L g202 ( .A(n_44), .Y(n_202) );
INVx1_ASAP7_75t_L g215 ( .A(n_46), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_47), .Y(n_196) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_48), .A2(n_64), .B1(n_90), .B2(n_91), .Y(n_97) );
A2O1A1Ixp33_ASAP7_75t_SL g322 ( .A1(n_49), .A2(n_252), .B(n_303), .C(n_323), .Y(n_322) );
INVxp67_ASAP7_75t_L g324 ( .A(n_50), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_52), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_53), .Y(n_317) );
INVx1_ASAP7_75t_L g262 ( .A(n_54), .Y(n_262) );
INVx1_ASAP7_75t_L g180 ( .A(n_55), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_55), .A2(n_224), .B(n_228), .C(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g189 ( .A(n_56), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_59), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g213 ( .A(n_60), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_61), .B(n_252), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_62), .A2(n_185), .B1(n_186), .B2(n_187), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_62), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_63), .A2(n_178), .B1(n_179), .B2(n_182), .Y(n_177) );
CKINVDCx14_ASAP7_75t_R g182 ( .A(n_63), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g333 ( .A1(n_63), .A2(n_224), .B(n_228), .C(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_65), .B(n_212), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_66), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g279 ( .A1(n_67), .A2(n_224), .B(n_228), .C(n_280), .Y(n_279) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_68), .Y(n_288) );
INVx1_ASAP7_75t_L g321 ( .A(n_69), .Y(n_321) );
CKINVDCx16_ASAP7_75t_R g226 ( .A(n_70), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_70), .A2(n_81), .B1(n_175), .B2(n_226), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_71), .B(n_249), .Y(n_281) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_72), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_73), .B(n_240), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_74), .A2(n_81), .B1(n_174), .B2(n_175), .Y(n_80) );
INVx2_ASAP7_75t_L g174 ( .A(n_74), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_75), .A2(n_219), .B(n_320), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_76), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_77), .Y(n_105) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_192), .B1(n_205), .B2(n_512), .C(n_515), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_176), .Y(n_79) );
INVx1_ASAP7_75t_L g175 ( .A(n_81), .Y(n_175) );
AND2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_138), .Y(n_81) );
NOR2xp33_ASAP7_75t_SL g82 ( .A(n_83), .B(n_117), .Y(n_82) );
OAI221xp5_ASAP7_75t_SL g83 ( .A1(n_84), .A2(n_100), .B1(n_101), .B2(n_105), .C(n_106), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_95), .Y(n_86) );
INVx2_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
OR2x2_ASAP7_75t_L g87 ( .A(n_88), .B(n_93), .Y(n_87) );
AND2x2_ASAP7_75t_L g104 ( .A(n_88), .B(n_93), .Y(n_104) );
AND2x2_ASAP7_75t_L g149 ( .A(n_88), .B(n_123), .Y(n_149) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g112 ( .A(n_89), .B(n_99), .Y(n_112) );
AND2x2_ASAP7_75t_L g116 ( .A(n_89), .B(n_93), .Y(n_116) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
INVx1_ASAP7_75t_L g111 ( .A(n_93), .Y(n_111) );
INVx2_ASAP7_75t_L g123 ( .A(n_93), .Y(n_123) );
INVx1_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
NAND2x1p5_ASAP7_75t_L g103 ( .A(n_96), .B(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g148 ( .A(n_96), .B(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_98), .Y(n_96) );
INVx1_ASAP7_75t_L g115 ( .A(n_97), .Y(n_115) );
INVx1_ASAP7_75t_L g122 ( .A(n_97), .Y(n_122) );
INVx1_ASAP7_75t_L g130 ( .A(n_97), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_97), .B(n_99), .Y(n_158) );
AND2x2_ASAP7_75t_L g129 ( .A(n_98), .B(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g155 ( .A(n_99), .B(n_115), .Y(n_155) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g154 ( .A(n_104), .B(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g166 ( .A(n_104), .B(n_129), .Y(n_166) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x6_ASAP7_75t_L g157 ( .A(n_111), .B(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g120 ( .A(n_112), .B(n_121), .Y(n_120) );
AND2x4_ASAP7_75t_L g135 ( .A(n_112), .B(n_136), .Y(n_135) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x6_ASAP7_75t_L g128 ( .A(n_116), .B(n_129), .Y(n_128) );
OAI222xp33_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_124), .B1(n_125), .B2(n_131), .C1(n_132), .C2(n_137), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g136 ( .A(n_122), .Y(n_136) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x6_ASAP7_75t_L g143 ( .A(n_129), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g163 ( .A(n_129), .B(n_149), .Y(n_163) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx4f_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
BUFx12f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_159), .Y(n_138) );
OAI221xp5_ASAP7_75t_SL g139 ( .A1(n_140), .A2(n_145), .B1(n_146), .B2(n_150), .C(n_151), .Y(n_139) );
INVx1_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx11_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g170 ( .A(n_149), .B(n_155), .Y(n_170) );
AND2x4_ASAP7_75t_L g172 ( .A(n_149), .B(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx8_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
NAND2xp33_ASAP7_75t_SL g159 ( .A(n_160), .B(n_167), .Y(n_159) );
BUFx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx6_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_183), .B1(n_184), .B2(n_191), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_177), .Y(n_191) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g193 ( .A(n_194), .Y(n_193) );
AND3x1_ASAP7_75t_SL g194 ( .A(n_195), .B(n_200), .C(n_203), .Y(n_194) );
INVxp67_ASAP7_75t_L g520 ( .A(n_195), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVx1_ASAP7_75t_SL g522 ( .A(n_200), .Y(n_522) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_200), .A2(n_220), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g533 ( .A(n_200), .Y(n_533) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_201), .B(n_204), .Y(n_526) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_SL g532 ( .A(n_203), .B(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_204), .Y(n_203) );
OR4x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_408), .C(n_467), .D(n_494), .Y(n_205) );
NAND3xp33_ASAP7_75t_SL g206 ( .A(n_207), .B(n_350), .C(n_375), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_273), .B(n_293), .C(n_326), .Y(n_207) );
AOI211xp5_ASAP7_75t_SL g498 ( .A1(n_208), .A2(n_499), .B(n_501), .C(n_504), .Y(n_498) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_242), .Y(n_208) );
INVx1_ASAP7_75t_L g373 ( .A(n_209), .Y(n_373) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_L g348 ( .A(n_210), .B(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g380 ( .A(n_210), .Y(n_380) );
AND2x2_ASAP7_75t_L g435 ( .A(n_210), .B(n_404), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_210), .B(n_291), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_210), .B(n_292), .Y(n_493) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g354 ( .A(n_211), .Y(n_354) );
AND2x2_ASAP7_75t_L g397 ( .A(n_211), .B(n_260), .Y(n_397) );
AND2x2_ASAP7_75t_L g415 ( .A(n_211), .B(n_292), .Y(n_415) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_217), .B(n_239), .Y(n_211) );
INVx1_ASAP7_75t_L g272 ( .A(n_212), .Y(n_272) );
INVx2_ASAP7_75t_L g277 ( .A(n_212), .Y(n_277) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g241 ( .A(n_213), .B(n_214), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_218), .Y(n_514) );
BUFx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_220), .B(n_224), .Y(n_263) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_223), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g229 ( .A(n_222), .Y(n_229) );
INVx1_ASAP7_75t_L g310 ( .A(n_222), .Y(n_310) );
INVx1_ASAP7_75t_L g230 ( .A(n_223), .Y(n_230) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
INVx3_ASAP7_75t_L g250 ( .A(n_223), .Y(n_250) );
INVx1_ASAP7_75t_L g252 ( .A(n_223), .Y(n_252) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_223), .Y(n_267) );
INVx4_ASAP7_75t_SL g238 ( .A(n_224), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_231), .C(n_238), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_227), .A2(n_238), .B(n_298), .C(n_299), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_227), .A2(n_238), .B(n_321), .C(n_322), .Y(n_320) );
INVx5_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
BUFx3_ASAP7_75t_L g237 ( .A(n_229), .Y(n_237) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_229), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_232), .B(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g311 ( .A1(n_233), .A2(n_312), .B1(n_313), .B2(n_314), .Y(n_311) );
INVx2_ASAP7_75t_L g313 ( .A(n_233), .Y(n_313) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g254 ( .A(n_237), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_238), .A2(n_263), .B1(n_308), .B2(n_315), .Y(n_307) );
INVx4_ASAP7_75t_L g259 ( .A(n_240), .Y(n_259) );
OA21x2_ASAP7_75t_L g318 ( .A1(n_240), .A2(n_319), .B(n_325), .Y(n_318) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g256 ( .A(n_241), .Y(n_256) );
INVx4_ASAP7_75t_L g347 ( .A(n_242), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g402 ( .A1(n_242), .A2(n_403), .B(n_405), .Y(n_402) );
AND2x2_ASAP7_75t_L g483 ( .A(n_242), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_260), .Y(n_242) );
INVx1_ASAP7_75t_L g290 ( .A(n_243), .Y(n_290) );
AND2x2_ASAP7_75t_L g352 ( .A(n_243), .B(n_292), .Y(n_352) );
OR2x2_ASAP7_75t_L g381 ( .A(n_243), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g395 ( .A(n_243), .Y(n_395) );
INVx3_ASAP7_75t_L g404 ( .A(n_243), .Y(n_404) );
AND2x2_ASAP7_75t_L g414 ( .A(n_243), .B(n_415), .Y(n_414) );
AND2x2_ASAP7_75t_L g447 ( .A(n_243), .B(n_353), .Y(n_447) );
AND2x2_ASAP7_75t_L g471 ( .A(n_243), .B(n_427), .Y(n_471) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_257), .Y(n_243) );
AOI21xp5_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_246), .B(n_255), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_251), .B(n_253), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_249), .A2(n_335), .B(n_336), .C(n_337), .Y(n_334) );
INVx5_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_250), .B(n_302), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_250), .B(n_324), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_253), .A2(n_266), .B(n_268), .Y(n_265) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g269 ( .A(n_255), .Y(n_269) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_256), .A2(n_307), .B(n_316), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_256), .B(n_317), .Y(n_316) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_256), .A2(n_331), .B(n_338), .Y(n_330) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx3_ASAP7_75t_L g295 ( .A(n_259), .Y(n_295) );
INVx2_ASAP7_75t_L g292 ( .A(n_260), .Y(n_292) );
AND2x2_ASAP7_75t_L g507 ( .A(n_260), .B(n_349), .Y(n_507) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_269), .B(n_270), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_264), .Y(n_261) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_263), .A2(n_332), .B(n_333), .Y(n_331) );
INVx4_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
INVx2_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_272), .B(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_272), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_289), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_275), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g427 ( .A(n_275), .B(n_415), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_275), .B(n_404), .Y(n_489) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g349 ( .A(n_276), .Y(n_349) );
AND2x2_ASAP7_75t_L g353 ( .A(n_276), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g394 ( .A(n_276), .B(n_395), .Y(n_394) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_287), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_286), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_284), .Y(n_280) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx3_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_289), .B(n_390), .Y(n_412) );
INVx1_ASAP7_75t_L g451 ( .A(n_289), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_289), .B(n_378), .Y(n_495) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g358 ( .A(n_290), .B(n_353), .Y(n_358) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_292), .B(n_349), .Y(n_382) );
INVx1_ASAP7_75t_L g461 ( .A(n_292), .Y(n_461) );
AOI322xp5_ASAP7_75t_L g485 ( .A1(n_293), .A2(n_400), .A3(n_460), .B1(n_486), .B2(n_488), .C1(n_490), .C2(n_492), .Y(n_485) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_294), .B(n_305), .Y(n_293) );
AND2x2_ASAP7_75t_L g340 ( .A(n_294), .B(n_318), .Y(n_340) );
INVx1_ASAP7_75t_SL g343 ( .A(n_294), .Y(n_343) );
AND2x2_ASAP7_75t_L g345 ( .A(n_294), .B(n_306), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_294), .B(n_362), .Y(n_368) );
INVx2_ASAP7_75t_L g387 ( .A(n_294), .Y(n_387) );
AND2x2_ASAP7_75t_L g400 ( .A(n_294), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g438 ( .A(n_294), .B(n_362), .Y(n_438) );
BUFx2_ASAP7_75t_L g455 ( .A(n_294), .Y(n_455) );
AND2x2_ASAP7_75t_L g469 ( .A(n_294), .B(n_329), .Y(n_469) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_304), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_305), .B(n_357), .Y(n_384) );
AND2x2_ASAP7_75t_L g511 ( .A(n_305), .B(n_387), .Y(n_511) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_318), .Y(n_305) );
OR2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_357), .Y(n_356) );
INVx3_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
AND2x2_ASAP7_75t_L g407 ( .A(n_306), .B(n_330), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_306), .B(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_306), .Y(n_491) );
INVx2_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g342 ( .A(n_318), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g364 ( .A(n_318), .Y(n_364) );
BUFx2_ASAP7_75t_L g370 ( .A(n_318), .Y(n_370) );
AND2x2_ASAP7_75t_L g389 ( .A(n_318), .B(n_362), .Y(n_389) );
INVx3_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
OR2x2_ASAP7_75t_L g411 ( .A(n_318), .B(n_362), .Y(n_411) );
AOI31xp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_341), .A3(n_344), .B(n_346), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_340), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_328), .B(n_363), .Y(n_374) );
OR2x2_ASAP7_75t_L g398 ( .A(n_328), .B(n_368), .Y(n_398) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_329), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g419 ( .A(n_329), .B(n_411), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_329), .B(n_401), .Y(n_429) );
AND2x2_ASAP7_75t_L g436 ( .A(n_329), .B(n_437), .Y(n_436) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_329), .B(n_400), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_329), .B(n_455), .Y(n_465) );
AND2x2_ASAP7_75t_L g477 ( .A(n_329), .B(n_362), .Y(n_477) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx3_ASAP7_75t_L g357 ( .A(n_330), .Y(n_357) );
INVx1_ASAP7_75t_L g423 ( .A(n_340), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_340), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_342), .B(n_418), .Y(n_452) );
AND2x4_ASAP7_75t_L g363 ( .A(n_343), .B(n_364), .Y(n_363) );
CKINVDCx16_ASAP7_75t_R g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx2_ASAP7_75t_L g442 ( .A(n_348), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_348), .B(n_460), .Y(n_459) );
AND2x2_ASAP7_75t_L g390 ( .A(n_349), .B(n_380), .Y(n_390) );
AND2x2_ASAP7_75t_L g484 ( .A(n_349), .B(n_354), .Y(n_484) );
INVx1_ASAP7_75t_L g509 ( .A(n_349), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_355), .B1(n_358), .B2(n_359), .C(n_365), .Y(n_350) );
CKINVDCx14_ASAP7_75t_R g371 ( .A(n_351), .Y(n_371) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_352), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_355), .B(n_406), .Y(n_425) );
INVx3_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OR2x2_ASAP7_75t_L g474 ( .A(n_356), .B(n_370), .Y(n_474) );
AND2x2_ASAP7_75t_L g388 ( .A(n_357), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g418 ( .A(n_357), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_357), .B(n_401), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g488 ( .A(n_357), .B(n_458), .C(n_489), .Y(n_488) );
AOI211xp5_ASAP7_75t_SL g421 ( .A1(n_358), .A2(n_422), .B(n_424), .C(n_432), .Y(n_421) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_360), .A2(n_411), .B1(n_412), .B2(n_413), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_361), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_361), .B(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g503 ( .A(n_363), .B(n_477), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_371), .B1(n_372), .B2(n_374), .Y(n_365) );
NOR2xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_369), .B(n_418), .Y(n_449) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_372), .A2(n_464), .B1(n_495), .B2(n_502), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_383), .B1(n_385), .B2(n_390), .C(n_391), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_381), .A2(n_392), .B1(n_398), .B2(n_399), .C(n_402), .Y(n_391) );
INVx1_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g406 ( .A(n_387), .Y(n_406) );
OR2x2_ASAP7_75t_L g479 ( .A(n_387), .B(n_411), .Y(n_479) );
AND2x2_ASAP7_75t_L g481 ( .A(n_387), .B(n_389), .Y(n_481) );
INVx1_ASAP7_75t_L g420 ( .A(n_390), .Y(n_420) );
OR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_396), .Y(n_392) );
AOI21xp33_ASAP7_75t_SL g450 ( .A1(n_393), .A2(n_451), .B(n_452), .Y(n_450) );
OR2x2_ASAP7_75t_L g457 ( .A(n_393), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g431 ( .A(n_394), .B(n_415), .Y(n_431) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp33_ASAP7_75t_SL g448 ( .A(n_399), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_400), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_401), .B(n_437), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g416 ( .A1(n_404), .A2(n_417), .B(n_419), .C(n_420), .Y(n_416) );
NAND2x1_ASAP7_75t_SL g441 ( .A(n_404), .B(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_405), .A2(n_454), .B1(n_456), .B2(n_459), .Y(n_453) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_407), .B(n_497), .Y(n_496) );
NAND5xp2_ASAP7_75t_L g408 ( .A(n_409), .B(n_421), .C(n_439), .D(n_453), .E(n_462), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g466 ( .A(n_412), .Y(n_466) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_414), .A2(n_433), .B1(n_473), .B2(n_475), .C(n_478), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_415), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_418), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_418), .B(n_484), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_428), .B2(n_430), .Y(n_424) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
AND2x2_ASAP7_75t_L g506 ( .A(n_435), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_443), .B1(n_447), .B2(n_448), .C(n_450), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g490 ( .A(n_445), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g497 ( .A(n_455), .Y(n_497) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI21xp5_ASAP7_75t_SL g462 ( .A1(n_463), .A2(n_465), .B(n_466), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI211xp5_ASAP7_75t_SL g467 ( .A1(n_468), .A2(n_470), .B(n_472), .C(n_485), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_470), .A2(n_495), .B(n_496), .C(n_498), .Y(n_494) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_474), .B(n_476), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B(n_482), .Y(n_478) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_508), .B(n_510), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_513), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
OAI322xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .A3(n_521), .B1(n_523), .B2(n_527), .C1(n_528), .C2(n_530), .Y(n_515) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
endmodule