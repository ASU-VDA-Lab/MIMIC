module fake_jpeg_17230_n_355 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_355);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_53),
.Y(n_66)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_55),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_77),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_20),
.C(n_39),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_32),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_38),
.B(n_39),
.C(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_37),
.Y(n_104)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_87),
.Y(n_136)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_58),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_90),
.B(n_24),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_59),
.A2(n_37),
.B1(n_22),
.B2(n_25),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_96),
.B1(n_112),
.B2(n_113),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_37),
.B1(n_22),
.B2(n_25),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_76),
.Y(n_100)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_64),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_105),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_83),
.A2(n_44),
.B1(n_29),
.B2(n_27),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_29),
.B1(n_32),
.B2(n_28),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_51),
.B1(n_36),
.B2(n_28),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_36),
.B1(n_24),
.B2(n_102),
.Y(n_142)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_73),
.Y(n_116)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_75),
.B1(n_68),
.B2(n_62),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_138),
.B1(n_102),
.B2(n_107),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_121),
.B(n_123),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_63),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_61),
.B(n_85),
.C(n_66),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_103),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_79),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_147),
.C(n_40),
.Y(n_165)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_140),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_115),
.A2(n_68),
.B1(n_62),
.B2(n_61),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

AOI32xp33_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_72),
.A3(n_78),
.B1(n_21),
.B2(n_34),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_72),
.B1(n_21),
.B2(n_40),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_145),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_65),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_146),
.B(n_34),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_21),
.B(n_40),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_145),
.Y(n_151)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_100),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_152),
.A2(n_164),
.B(n_40),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_159),
.B1(n_169),
.B2(n_136),
.Y(n_180)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_168),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_116),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_172),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_122),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_167),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_87),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_35),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_0),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_172),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_117),
.B(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_170),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_128),
.Y(n_167)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_109),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_129),
.A2(n_103),
.B1(n_35),
.B2(n_21),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_136),
.C(n_130),
.Y(n_172)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_132),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_150),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_125),
.B(n_21),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_197),
.B(n_169),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_152),
.A2(n_171),
.B1(n_159),
.B2(n_149),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_178),
.A2(n_182),
.B1(n_189),
.B2(n_190),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_151),
.B1(n_167),
.B2(n_161),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_138),
.A3(n_35),
.B1(n_40),
.B2(n_126),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_153),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_172),
.A2(n_141),
.B1(n_118),
.B2(n_124),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_183),
.B(n_185),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_2),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_186),
.C(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_192),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_143),
.B1(n_119),
.B2(n_131),
.Y(n_189)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_98),
.B(n_119),
.C(n_143),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_166),
.Y(n_205)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_195),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_165),
.A2(n_19),
.B(n_3),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_198),
.B(n_200),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_194),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_187),
.Y(n_200)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_205),
.Y(n_242)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_209),
.Y(n_231)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_213),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_162),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.Y(n_232)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_192),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_215),
.Y(n_227)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_223),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_218),
.B1(n_219),
.B2(n_191),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_188),
.A2(n_156),
.B1(n_150),
.B2(n_163),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_221),
.Y(n_238)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

INVx4_ASAP7_75t_SL g222 ( 
.A(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_191),
.B1(n_190),
.B2(n_160),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_158),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_156),
.B(n_158),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_224),
.B(n_184),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_181),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_202),
.Y(n_253)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_226),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_219),
.B(n_186),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_230),
.A2(n_247),
.B(n_249),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_243),
.C(n_203),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_160),
.Y(n_236)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_222),
.B1(n_212),
.B2(n_204),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_190),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_240),
.B(n_244),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_207),
.A2(n_190),
.B1(n_194),
.B2(n_160),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_246),
.B1(n_222),
.B2(n_214),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_224),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_2),
.Y(n_244)
);

NOR4xp25_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_173),
.C(n_168),
.D(n_155),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_245),
.A2(n_173),
.B(n_98),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_216),
.A2(n_220),
.B1(n_221),
.B2(n_217),
.Y(n_246)
);

NAND2x1_ASAP7_75t_L g247 ( 
.A(n_201),
.B(n_168),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_200),
.B(n_198),
.Y(n_248)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_213),
.B(n_155),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_256),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_261),
.B1(n_269),
.B2(n_249),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_223),
.C(n_204),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_239),
.C(n_227),
.Y(n_282)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_209),
.Y(n_259)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_232),
.B(n_157),
.Y(n_260)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_260),
.Y(n_290)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_262),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_271),
.Y(n_272)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_249),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_132),
.B1(n_4),
.B2(n_5),
.Y(n_269)
);

AO21x1_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_19),
.B(n_4),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_279),
.B1(n_226),
.B2(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_243),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_278),
.C(n_256),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_230),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_265),
.A2(n_230),
.B1(n_238),
.B2(n_241),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_270),
.B(n_244),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_281),
.B(n_284),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_157),
.Y(n_304)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_254),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_266),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_242),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_267),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_294),
.Y(n_311)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_272),
.A2(n_238),
.B(n_268),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_295),
.B(n_296),
.Y(n_308)
);

OAI322xp33_ASAP7_75t_L g294 ( 
.A1(n_275),
.A2(n_225),
.A3(n_227),
.B1(n_257),
.B2(n_258),
.C1(n_253),
.C2(n_263),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_282),
.A2(n_268),
.B(n_250),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_273),
.B(n_250),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_246),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_300),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_280),
.A2(n_269),
.B(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_242),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_302),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_264),
.B(n_271),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_6),
.B(n_7),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_278),
.C(n_276),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_288),
.A2(n_106),
.B(n_91),
.C(n_157),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_18),
.B(n_7),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_290),
.B1(n_285),
.B2(n_283),
.Y(n_309)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_277),
.C(n_19),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_277),
.C(n_19),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_3),
.C(n_5),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_317),
.C(n_8),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_3),
.C(n_5),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_6),
.B(n_8),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_8),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_305),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_321),
.B(n_322),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_306),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_323),
.B(n_328),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_325),
.B(n_327),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_306),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_326),
.B(n_329),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_306),
.C(n_9),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_316),
.B(n_10),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_10),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_SL g335 ( 
.A1(n_326),
.A2(n_315),
.B(n_308),
.C(n_311),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_335),
.A2(n_332),
.B(n_340),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_331),
.A2(n_313),
.B(n_312),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_336),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_324),
.A2(n_330),
.B(n_12),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_337),
.B(n_13),
.Y(n_345)
);

AOI31xp67_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_11),
.A3(n_13),
.B(n_14),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_339),
.B(n_11),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_334),
.B(n_11),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_343),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_332),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g343 ( 
.A(n_338),
.B(n_18),
.CI(n_13),
.CON(n_343),
.SN(n_343)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_344),
.B(n_345),
.Y(n_349)
);

OAI21xp33_ASAP7_75t_SL g350 ( 
.A1(n_348),
.A2(n_346),
.B(n_342),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_333),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_347),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_352),
.B(n_349),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_14),
.C(n_17),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_17),
.Y(n_355)
);


endmodule