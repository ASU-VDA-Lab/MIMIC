module fake_jpeg_3999_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OR2x2_ASAP7_75t_SL g28 ( 
.A(n_6),
.B(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_43),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_26),
.B1(n_16),
.B2(n_19),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_63),
.B1(n_27),
.B2(n_32),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_19),
.B1(n_16),
.B2(n_25),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_26),
.C(n_29),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_30),
.C(n_29),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_34),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_17),
.B1(n_28),
.B2(n_24),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_64),
.Y(n_83)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_69),
.Y(n_86)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_71),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_20),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_67),
.B(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_20),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_77),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_70),
.B1(n_40),
.B2(n_18),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_28),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_48),
.A2(n_52),
.B(n_55),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_38),
.C(n_36),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_20),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_32),
.Y(n_85)
);

NAND2xp67_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_32),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_93),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_30),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_38),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_22),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_47),
.A2(n_37),
.B1(n_39),
.B2(n_69),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_107)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_115),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_51),
.B1(n_47),
.B2(n_65),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_62),
.B1(n_51),
.B2(n_46),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_105),
.B1(n_112),
.B2(n_85),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_113),
.B1(n_125),
.B2(n_93),
.Y(n_128)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_46),
.B1(n_39),
.B2(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_59),
.B1(n_45),
.B2(n_38),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_121),
.C(n_124),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_13),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_15),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_36),
.C(n_45),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_82),
.A2(n_59),
.B1(n_18),
.B2(n_31),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_128),
.A2(n_97),
.B1(n_106),
.B2(n_2),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_77),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_SL g171 ( 
.A(n_129),
.B(n_131),
.C(n_153),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_124),
.B(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_101),
.B(n_77),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_137),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_92),
.B(n_78),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_142),
.B(n_147),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_144),
.B1(n_145),
.B2(n_75),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_73),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_143),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_76),
.B1(n_93),
.B2(n_95),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_151),
.B1(n_104),
.B2(n_112),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_79),
.B(n_93),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_95),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_105),
.A2(n_115),
.B1(n_104),
.B2(n_116),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_75),
.B1(n_94),
.B2(n_81),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_122),
.B(n_83),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_83),
.C(n_80),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_106),
.C(n_15),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_113),
.A2(n_75),
.B1(n_94),
.B2(n_81),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_90),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_22),
.B(n_18),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_154),
.B(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_159),
.B1(n_178),
.B2(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_161),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_99),
.B(n_98),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_163),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_107),
.B1(n_125),
.B2(n_94),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_136),
.B(n_108),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_168),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_81),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_175),
.B1(n_179),
.B2(n_142),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_165),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_166),
.A2(n_167),
.B(n_127),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_131),
.A2(n_22),
.B(n_33),
.C(n_31),
.D(n_21),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_151),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_173),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_22),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_176),
.C(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_139),
.A2(n_97),
.B1(n_109),
.B2(n_31),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_174),
.A2(n_132),
.B1(n_148),
.B2(n_127),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_15),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_141),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_138),
.A2(n_14),
.B1(n_13),
.B2(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_184),
.A2(n_203),
.B1(n_155),
.B2(n_169),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_185),
.A2(n_195),
.B1(n_201),
.B2(n_189),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_165),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_201),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_192),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_198),
.CI(n_144),
.CON(n_219),
.SN(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_195),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_164),
.Y(n_195)
);

AND2x4_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_166),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_147),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_149),
.C(n_153),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_149),
.C(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_160),
.B1(n_159),
.B2(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_204),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_163),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_221),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_220),
.C(n_223),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_219),
.B(n_182),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_177),
.C(n_129),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_129),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_191),
.B(n_129),
.C(n_152),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_224),
.A2(n_232),
.B1(n_194),
.B2(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_126),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_202),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_126),
.C(n_134),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_230),
.C(n_233),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_190),
.C(n_187),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_136),
.B1(n_134),
.B2(n_137),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_193),
.C(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_185),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_237),
.C(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_239),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_186),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_240),
.B(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_186),
.Y(n_241)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_244),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_222),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_206),
.C(n_184),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_218),
.B1(n_224),
.B2(n_232),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_208),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_0),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_202),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_251),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_233),
.Y(n_252)
);

XNOR2x1_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_221),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_0),
.C(n_1),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_223),
.C(n_229),
.Y(n_258)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_264),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_262),
.C(n_267),
.Y(n_277)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

INVx11_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_265),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_219),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_236),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_209),
.C(n_1),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_0),
.C(n_3),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_270),
.C(n_235),
.Y(n_278)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_269),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_235),
.C(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_245),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_275),
.A2(n_284),
.B(n_268),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_283),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_274),
.B(n_251),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_286),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_257),
.A2(n_252),
.B1(n_234),
.B2(n_246),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_253),
.B1(n_4),
.B2(n_5),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_274),
.A2(n_3),
.B(n_4),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_290),
.B(n_5),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_265),
.A2(n_5),
.B(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_271),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_294),
.B(n_296),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_267),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_272),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_256),
.B(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_302),
.C(n_276),
.Y(n_313)
);

NOR3xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_299),
.C(n_14),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_259),
.B1(n_258),
.B2(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_260),
.B(n_263),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_301),
.A2(n_289),
.B(n_284),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_287),
.C(n_281),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_287),
.B(n_7),
.CI(n_8),
.CON(n_304),
.SN(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_291),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_311),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_279),
.B(n_290),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_313),
.C(n_315),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_298),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_314),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_293),
.A2(n_9),
.B(n_10),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_312),
.B(n_302),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_295),
.C(n_8),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_321),
.B(n_323),
.Y(n_327)
);

AOI21x1_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_304),
.B(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_308),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_325),
.B(n_326),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_317),
.A2(n_293),
.B(n_304),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_318),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_320),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_330),
.C(n_327),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_319),
.B(n_13),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_8),
.B(n_104),
.Y(n_334)
);


endmodule