module fake_jpeg_4488_n_307 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_41),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_8),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_8),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_19),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_46),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_51),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_35),
.A2(n_18),
.B(n_31),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_48),
.A2(n_49),
.B(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_18),
.B1(n_31),
.B2(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_38),
.A2(n_18),
.B1(n_31),
.B2(n_25),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_61),
.B1(n_28),
.B2(n_29),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_19),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_34),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_27),
.B1(n_32),
.B2(n_17),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_39),
.C(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_32),
.B1(n_25),
.B2(n_17),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_32),
.B1(n_34),
.B2(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_34),
.B1(n_21),
.B2(n_29),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_42),
.B1(n_30),
.B2(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_69),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_70),
.B(n_72),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

INVx5_ASAP7_75t_SL g103 ( 
.A(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_45),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_28),
.B1(n_21),
.B2(n_24),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_75),
.A2(n_86),
.B1(n_64),
.B2(n_47),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_76),
.A2(n_46),
.B(n_65),
.Y(n_95)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_85),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_39),
.B1(n_40),
.B2(n_30),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_91),
.A2(n_92),
.B1(n_63),
.B2(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_94),
.A2(n_109),
.B1(n_93),
.B2(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_91),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_83),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_48),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_54),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_113),
.Y(n_125)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_96),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_89),
.A2(n_49),
.B1(n_42),
.B2(n_53),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_107),
.A2(n_77),
.B1(n_76),
.B2(n_79),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_66),
.B(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_44),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_43),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_43),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_0),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_43),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_43),
.B(n_23),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_104),
.B(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_105),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_72),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_134),
.B1(n_139),
.B2(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_80),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_141),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_105),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_81),
.B1(n_77),
.B2(n_83),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_142),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_69),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_71),
.B1(n_78),
.B2(n_40),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_145),
.B(n_142),
.Y(n_178)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_78),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_109),
.B1(n_99),
.B2(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_82),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_103),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_99),
.A2(n_92),
.B1(n_70),
.B2(n_71),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_103),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_107),
.A2(n_40),
.B1(n_59),
.B2(n_52),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_109),
.A2(n_40),
.B1(n_60),
.B2(n_87),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_160),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_119),
.B1(n_113),
.B2(n_102),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_152),
.A2(n_163),
.B1(n_169),
.B2(n_179),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_113),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_154),
.B(n_162),
.C(n_180),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_171),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_159),
.A2(n_168),
.B1(n_133),
.B2(n_121),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_104),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_129),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_117),
.C(n_101),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_149),
.A2(n_94),
.B1(n_95),
.B2(n_115),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_165),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_112),
.B(n_115),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_177),
.B(n_178),
.Y(n_191)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_170),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_59),
.B1(n_103),
.B2(n_108),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_95),
.B1(n_117),
.B2(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_97),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_114),
.Y(n_175)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_175),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_120),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_141),
.A2(n_110),
.B1(n_116),
.B2(n_87),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_43),
.C(n_59),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_182),
.B1(n_190),
.B2(n_204),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_139),
.B(n_134),
.C(n_147),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_192),
.Y(n_230)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_194),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_159),
.B1(n_150),
.B2(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_163),
.A2(n_135),
.B1(n_121),
.B2(n_144),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_198),
.A2(n_26),
.B1(n_23),
.B2(n_22),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_132),
.B(n_128),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_26),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_137),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g205 ( 
.A(n_158),
.B(n_131),
.C(n_126),
.Y(n_205)
);

NOR3xp33_ASAP7_75t_SL g218 ( 
.A(n_205),
.B(n_177),
.C(n_174),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_130),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_206),
.B(n_171),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_170),
.B1(n_151),
.B2(n_153),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_208),
.B(n_226),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_169),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_154),
.C(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_166),
.C(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_152),
.C(n_177),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_221),
.B1(n_187),
.B2(n_199),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_153),
.C(n_173),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_224),
.C(n_188),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_131),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_43),
.C(n_60),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_228),
.Y(n_245)
);

OA21x2_ASAP7_75t_SL g226 ( 
.A1(n_205),
.A2(n_26),
.B(n_43),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_227),
.A2(n_231),
.B1(n_184),
.B2(n_186),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_198),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_60),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_192),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_194),
.A2(n_23),
.B1(n_26),
.B2(n_22),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_9),
.Y(n_263)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_235),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_221),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_246),
.C(n_22),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_222),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_240),
.B(n_241),
.Y(n_265)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_182),
.B1(n_200),
.B2(n_189),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_243),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_213),
.A2(n_182),
.B1(n_185),
.B2(n_183),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_244),
.A2(n_250),
.B1(n_9),
.B2(n_16),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_193),
.C(n_186),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_247),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_22),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_219),
.A2(n_204),
.B1(n_11),
.B2(n_12),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_218),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_253),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_247),
.A2(n_216),
.B1(n_214),
.B2(n_212),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_255),
.A2(n_256),
.B1(n_236),
.B2(n_249),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_229),
.B1(n_228),
.B2(n_223),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_60),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_262),
.C(n_237),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_114),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g259 ( 
.A(n_239),
.B(n_220),
.CI(n_23),
.CON(n_259),
.SN(n_259)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_10),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_268),
.C(n_274),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_237),
.C(n_234),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_269),
.A2(n_271),
.B1(n_263),
.B2(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_245),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_82),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_272),
.B(n_260),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_8),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_0),
.C(n_1),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_252),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_255),
.C(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_286),
.C(n_274),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_0),
.C(n_2),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_7),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_5),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_7),
.B(n_15),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_288),
.A2(n_278),
.B(n_7),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_282),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_11),
.B(n_14),
.Y(n_293)
);

AOI31xp67_ASAP7_75t_SL g298 ( 
.A1(n_294),
.A2(n_296),
.A3(n_13),
.B(n_16),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_3),
.Y(n_296)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_286),
.A3(n_281),
.B1(n_284),
.B2(n_6),
.C1(n_12),
.C2(n_13),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_301),
.B(n_294),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g301 ( 
.A1(n_290),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_16),
.C1(n_292),
.C2(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_300),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_302),
.A2(n_303),
.B(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_304),
.B(n_4),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_4),
.Y(n_307)
);


endmodule