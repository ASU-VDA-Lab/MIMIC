module fake_jpeg_23040_n_180 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_38),
.Y(n_44)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_36),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_35),
.B1(n_2),
.B2(n_7),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_30),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_53),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_22),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_60),
.B(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_19),
.B1(n_39),
.B2(n_41),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_64),
.A2(n_73),
.B1(n_45),
.B2(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_24),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_21),
.B1(n_33),
.B2(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_69),
.B1(n_71),
.B2(n_80),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_58),
.A2(n_47),
.B1(n_46),
.B2(n_59),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_25),
.B1(n_26),
.B2(n_22),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_43),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_20),
.B1(n_26),
.B2(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_20),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_35),
.B(n_23),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

OAI22x1_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_58),
.B1(n_43),
.B2(n_45),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_60),
.B1(n_70),
.B2(n_79),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_2),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_99),
.B(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_5),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_5),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_96),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_75),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_110),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_105),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_101),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_113),
.Y(n_131)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_114),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_75),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_119),
.A2(n_97),
.B1(n_87),
.B2(n_62),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_95),
.B(n_96),
.Y(n_123)
);

HAxp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_89),
.CON(n_143),
.SN(n_143)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_122),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_111),
.B1(n_63),
.B2(n_117),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_113),
.A2(n_112),
.B1(n_108),
.B2(n_116),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_129),
.B1(n_83),
.B2(n_107),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_87),
.B1(n_84),
.B2(n_73),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_132),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_76),
.C(n_88),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_76),
.C(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_134),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_119),
.C(n_94),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_140),
.B(n_142),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_121),
.B1(n_122),
.B2(n_135),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_148),
.B(n_134),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_107),
.C(n_10),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_7),
.C(n_11),
.Y(n_148)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_123),
.B(n_133),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_156),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_124),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_161),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_128),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_136),
.C(n_152),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_153),
.Y(n_168)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_148),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_150),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_162),
.B(n_151),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_140),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_146),
.C(n_129),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_171),
.A2(n_173),
.B(n_12),
.Y(n_176)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_169),
.B1(n_167),
.B2(n_139),
.Y(n_174)
);

NAND4xp25_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_159),
.C(n_120),
.D(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_SL g178 ( 
.A1(n_176),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_14),
.B(n_172),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);


endmodule