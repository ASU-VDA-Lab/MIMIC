module real_jpeg_9492_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_1),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_10),
.B(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_2),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_2),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_2),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_28),
.B1(n_31),
.B2(n_45),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_8),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_9),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_9),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_9),
.A2(n_35),
.B1(n_86),
.B2(n_111),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_10),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_10),
.B(n_23),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_10),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_84),
.B1(n_86),
.B2(n_111),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_10),
.A2(n_31),
.B(n_59),
.C(n_67),
.D(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_10),
.B(n_31),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_10),
.B(n_27),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_10),
.A2(n_46),
.B(n_137),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_23),
.B(n_36),
.C(n_72),
.D(n_167),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_11),
.A2(n_28),
.B1(n_31),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_11),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_65),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_65),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_91),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_12),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_25),
.B1(n_41),
.B2(n_42),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_117),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_115),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_18),
.B(n_79),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_57),
.C(n_70),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_19),
.B(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_38),
.B2(n_56),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_50),
.C(n_54),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_32),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_22),
.A2(n_26),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_27),
.B(n_29),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_26),
.B(n_34),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_28),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_28),
.B(n_30),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_31),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_42),
.B1(n_60),
.B2(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_41),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_41),
.B(n_156),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_42),
.A2(n_62),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_46),
.A2(n_136),
.B(n_137),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_46),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_47),
.A2(n_143),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_47),
.B(n_84),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_51),
.B(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_53),
.B(n_86),
.C(n_109),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_53),
.B(n_86),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_57),
.B(n_70),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_64),
.B(n_66),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_58),
.A2(n_64),
.B1(n_68),
.B2(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_68),
.A2(n_99),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_68),
.B(n_84),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_69),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_75),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_71),
.B(n_75),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_77),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_95),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_81),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_106),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_105),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_97),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_173),
.B(n_177),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_160),
.B(n_172),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_139),
.B(n_159),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_121),
.B(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_124),
.B1(n_125),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_133),
.C(n_135),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_136),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_148),
.B(n_158),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_146),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_153),
.B(n_157),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_150),
.B(n_151),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_162),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_170),
.B2(n_171),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_165),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_166),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_170),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_174),
.B(n_175),
.Y(n_177)
);


endmodule