module fake_jpeg_5106_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_0),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_15),
.B(n_18),
.Y(n_24)
);

OR2x2_ASAP7_75t_SL g16 ( 
.A(n_7),
.B(n_11),
.Y(n_16)
);

XNOR2x1_ASAP7_75t_SL g25 ( 
.A(n_16),
.B(n_21),
.Y(n_25)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_20),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_4),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_22),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_4),
.B1(n_8),
.B2(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_6),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_23),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_21),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_28),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_32),
.B(n_29),
.C(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_20),
.Y(n_39)
);

OAI33xp33_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_33),
.A3(n_34),
.B1(n_28),
.B2(n_16),
.B3(n_10),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

OAI21x1_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_34),
.B(n_10),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_8),
.Y(n_42)
);


endmodule