module fake_jpeg_13946_n_593 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_593);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_593;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_575;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_14),
.B(n_5),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_9),
.C(n_2),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_59),
.B(n_64),
.Y(n_146)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_9),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_65),
.Y(n_130)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_66),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_53),
.B(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_71),
.B(n_74),
.Y(n_163)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_73),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_23),
.B(n_10),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_29),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_23),
.B(n_10),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_32),
.Y(n_135)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_86),
.Y(n_167)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_29),
.Y(n_88)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_33),
.B(n_10),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_99),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_22),
.B(n_27),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_107),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_72),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_125),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_65),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_109),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_135),
.B(n_36),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_57),
.A2(n_21),
.B1(n_22),
.B2(n_48),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_41),
.B1(n_28),
.B2(n_36),
.Y(n_182)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_64),
.A2(n_97),
.B1(n_74),
.B2(n_82),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_156),
.A2(n_162),
.B1(n_34),
.B2(n_37),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_61),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_21),
.B1(n_48),
.B2(n_41),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_56),
.A2(n_32),
.B1(n_43),
.B2(n_38),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_42),
.B(n_37),
.Y(n_207)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_92),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_63),
.B(n_27),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_28),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_176),
.B(n_185),
.Y(n_253)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_177),
.Y(n_283)
);

INVx3_ASAP7_75t_SL g178 ( 
.A(n_116),
.Y(n_178)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_178),
.Y(n_270)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_120),
.Y(n_180)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_183),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_182),
.A2(n_222),
.B1(n_46),
.B2(n_38),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_121),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_184),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_126),
.B(n_42),
.Y(n_185)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g293 ( 
.A(n_186),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_187),
.B(n_196),
.Y(n_291)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_194),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_50),
.B1(n_100),
.B2(n_86),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_195),
.A2(n_224),
.B1(n_227),
.B2(n_229),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_197),
.Y(n_255)
);

AO22x2_ASAP7_75t_L g198 ( 
.A1(n_144),
.A2(n_104),
.B1(n_108),
.B2(n_84),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_198),
.B(n_230),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_164),
.A2(n_81),
.B1(n_98),
.B2(n_91),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_199),
.A2(n_228),
.B1(n_239),
.B2(n_151),
.Y(n_276)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_202),
.B(n_208),
.Y(n_259)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_204),
.Y(n_264)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_50),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_206),
.A2(n_138),
.B(n_112),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_163),
.B(n_40),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_209),
.Y(n_262)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_129),
.Y(n_210)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_210),
.Y(n_280)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_150),
.Y(n_211)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_211),
.Y(n_281)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_212),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_213),
.B(n_220),
.Y(n_261)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_131),
.Y(n_214)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx11_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_157),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_130),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_163),
.B(n_44),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_130),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_221),
.Y(n_246)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_115),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_174),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_134),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_225),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_153),
.A2(n_67),
.B1(n_85),
.B2(n_78),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_160),
.B1(n_159),
.B2(n_154),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_128),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_146),
.A2(n_44),
.B1(n_40),
.B2(n_52),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_137),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_146),
.B(n_52),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_231),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_117),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_232),
.Y(n_287)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_233),
.Y(n_292)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_119),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_174),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_236),
.B(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_111),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_140),
.A2(n_38),
.B1(n_80),
.B2(n_109),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_176),
.A2(n_161),
.B(n_127),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_241),
.A2(n_268),
.B(n_1),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_162),
.C(n_50),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_242),
.B(n_12),
.C(n_5),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_244),
.B(n_276),
.Y(n_314)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_46),
.B(n_114),
.C(n_141),
.Y(n_248)
);

AO22x1_ASAP7_75t_L g302 ( 
.A1(n_248),
.A2(n_256),
.B1(n_257),
.B2(n_218),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_277),
.B1(n_215),
.B2(n_224),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_123),
.B(n_80),
.C(n_143),
.Y(n_256)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_198),
.A2(n_142),
.B(n_124),
.C(n_140),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_258),
.A2(n_266),
.B1(n_184),
.B2(n_193),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_198),
.A2(n_160),
.B1(n_159),
.B2(n_154),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_182),
.A2(n_198),
.B1(n_199),
.B2(n_191),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_195),
.A2(n_38),
.B(n_2),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_179),
.B(n_137),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_274),
.B(n_178),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_182),
.A2(n_151),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_201),
.A2(n_10),
.B(n_3),
.C(n_4),
.Y(n_278)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_278),
.A2(n_253),
.A3(n_243),
.B1(n_248),
.B2(n_251),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_226),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_286),
.A2(n_295),
.B1(n_1),
.B2(n_19),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_188),
.A2(n_192),
.B1(n_231),
.B2(n_180),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_238),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_297),
.B(n_305),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_186),
.B1(n_229),
.B2(n_227),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_298),
.A2(n_304),
.B1(n_326),
.B2(n_331),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_299),
.B(n_318),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_300),
.A2(n_330),
.B1(n_272),
.B2(n_287),
.Y(n_372)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g370 ( 
.A(n_302),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_260),
.A2(n_232),
.B1(n_234),
.B2(n_216),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_259),
.B(n_189),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_253),
.B(n_259),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_313),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_266),
.A2(n_194),
.B1(n_196),
.B2(n_5),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_308),
.Y(n_353)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_247),
.Y(n_311)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_312),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_315),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_243),
.B(n_11),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_316),
.B(n_347),
.C(n_325),
.Y(n_391)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_317),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_261),
.B(n_12),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_283),
.A2(n_12),
.B1(n_3),
.B2(n_5),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_319),
.A2(n_256),
.B(n_245),
.Y(n_352)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_248),
.A2(n_256),
.B(n_252),
.Y(n_322)
);

BUFx12f_ASAP7_75t_SL g360 ( 
.A(n_322),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_246),
.B(n_279),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_324),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_296),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_246),
.B(n_1),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_329),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_15),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_328),
.Y(n_375)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_290),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_257),
.A2(n_15),
.B1(n_6),
.B2(n_7),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_276),
.A2(n_1),
.B1(n_6),
.B2(n_8),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_250),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_332),
.B(n_333),
.Y(n_381)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_262),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_280),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_337),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_6),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_335),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_336),
.A2(n_302),
.B(n_327),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_295),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_280),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_338),
.B(n_341),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_244),
.A2(n_8),
.B1(n_16),
.B2(n_17),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_345),
.B1(n_346),
.B2(n_245),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_275),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_265),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_342),
.Y(n_368)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_343),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_16),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_344),
.B(n_296),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_268),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_257),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_241),
.B(n_18),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_348),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_340),
.A2(n_286),
.B1(n_285),
.B2(n_242),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_354),
.B1(n_356),
.B2(n_372),
.Y(n_396)
);

AOI21xp33_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_389),
.B(n_376),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_340),
.A2(n_242),
.B1(n_258),
.B2(n_293),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_300),
.A2(n_293),
.B1(n_282),
.B2(n_263),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_366),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_336),
.A2(n_278),
.B(n_273),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_385),
.B(n_390),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_314),
.A2(n_273),
.B(n_287),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_365),
.A2(n_302),
.B(n_341),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_314),
.A2(n_293),
.B1(n_283),
.B2(n_292),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_298),
.B1(n_337),
.B2(n_323),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_377),
.B(n_316),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_301),
.A2(n_272),
.B1(n_283),
.B2(n_289),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_382),
.A2(n_388),
.B1(n_392),
.B2(n_356),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_314),
.A2(n_292),
.B(n_284),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_308),
.A2(n_272),
.B1(n_289),
.B2(n_249),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_347),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_309),
.A2(n_288),
.B1(n_284),
.B2(n_281),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_394),
.A2(n_407),
.B(n_412),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_397),
.B(n_393),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_350),
.B(n_310),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_405),
.C(n_411),
.Y(n_434)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_371),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_401),
.A2(n_372),
.B1(n_353),
.B2(n_369),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_425),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_306),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_403),
.B(n_404),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_386),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_386),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_406),
.B(n_418),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_349),
.A2(n_331),
.B1(n_326),
.B2(n_345),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_408),
.A2(n_420),
.B1(n_358),
.B2(n_361),
.Y(n_439)
);

A2O1A1O1Ixp25_ASAP7_75t_L g409 ( 
.A1(n_350),
.A2(n_339),
.B(n_344),
.C(n_312),
.D(n_311),
.Y(n_409)
);

OAI31xp33_ASAP7_75t_L g457 ( 
.A1(n_409),
.A2(n_413),
.A3(n_415),
.B(n_379),
.Y(n_457)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_333),
.C(n_338),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_370),
.A2(n_334),
.B(n_321),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_370),
.A2(n_343),
.B(n_329),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_366),
.B(n_369),
.C(n_351),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_414),
.B(n_417),
.C(n_419),
.Y(n_450)
);

AO22x2_ASAP7_75t_SL g415 ( 
.A1(n_360),
.A2(n_330),
.B1(n_315),
.B2(n_317),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_416),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_288),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_381),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_366),
.B(n_240),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_354),
.A2(n_332),
.B1(n_320),
.B2(n_324),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_421),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_249),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_422),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_362),
.B(n_255),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_423),
.Y(n_451)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_387),
.Y(n_424)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_368),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_429),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_381),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_427),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_351),
.B(n_240),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_412),
.C(n_374),
.Y(n_455)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_387),
.Y(n_430)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_431),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_365),
.Y(n_432)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_432),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_435),
.A2(n_446),
.B1(n_424),
.B2(n_380),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_353),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_437),
.B(n_444),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_415),
.A2(n_360),
.B1(n_390),
.B2(n_364),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_438),
.A2(n_358),
.B1(n_429),
.B2(n_425),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_439),
.A2(n_401),
.B1(n_415),
.B2(n_413),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_398),
.B(n_405),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_SL g484 ( 
.A(n_441),
.B(n_408),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_453),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_357),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_410),
.A2(n_352),
.B1(n_388),
.B2(n_382),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_357),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_452),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_414),
.B(n_393),
.Y(n_452)
);

XOR2x2_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_360),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_462),
.C(n_422),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_428),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_409),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_457),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_395),
.B(n_416),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_461),
.B(n_464),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_399),
.B(n_363),
.C(n_367),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_399),
.B(n_363),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_473),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_465),
.B(n_359),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_469),
.B(n_483),
.Y(n_509)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_466),
.Y(n_470)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_470),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_471),
.A2(n_487),
.B1(n_438),
.B2(n_433),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_396),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_450),
.B(n_422),
.C(n_396),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_486),
.C(n_492),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_475),
.B(n_476),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_368),
.Y(n_477)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_477),
.Y(n_505)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_482),
.Y(n_522)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_443),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_484),
.B(n_496),
.Y(n_503)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_485),
.B(n_489),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_434),
.B(n_407),
.C(n_420),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_439),
.A2(n_415),
.B1(n_426),
.B2(n_402),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_497),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_380),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_446),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_490),
.A2(n_493),
.B1(n_458),
.B2(n_459),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_434),
.B(n_392),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_495),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_441),
.B(n_431),
.C(n_379),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_463),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_448),
.B(n_359),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_444),
.B(n_383),
.Y(n_497)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_473),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_500),
.B(n_375),
.Y(n_524)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_506),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_480),
.A2(n_457),
.B(n_460),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_507),
.A2(n_513),
.B(n_451),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_437),
.C(n_455),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_510),
.B(n_511),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_468),
.B(n_497),
.C(n_479),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_480),
.A2(n_460),
.B(n_436),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_479),
.B(n_452),
.C(n_462),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_514),
.B(n_476),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_472),
.B(n_453),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_515),
.B(n_519),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_490),
.A2(n_433),
.B1(n_436),
.B2(n_440),
.Y(n_517)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

FAx1_ASAP7_75t_SL g518 ( 
.A(n_492),
.B(n_464),
.CI(n_461),
.CON(n_518),
.SN(n_518)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_518),
.B(n_510),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_472),
.B(n_442),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_459),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_487),
.Y(n_538)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_521),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_507),
.A2(n_474),
.B(n_471),
.Y(n_523)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_524),
.B(n_525),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_498),
.B(n_481),
.C(n_494),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_498),
.B(n_481),
.C(n_494),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_526),
.B(n_530),
.C(n_536),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_484),
.C(n_496),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_516),
.Y(n_531)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_531),
.Y(n_545)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_508),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_540),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_514),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_535),
.B(n_539),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_504),
.B(n_520),
.C(n_511),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_505),
.B(n_517),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_537),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_538),
.B(n_502),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_509),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_513),
.A2(n_375),
.B1(n_355),
.B2(n_383),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_542),
.A2(n_378),
.B1(n_348),
.B2(n_342),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_559),
.Y(n_565)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_546),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_538),
.B(n_515),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_530),
.Y(n_566)
);

OAI31xp67_ASAP7_75t_L g549 ( 
.A1(n_537),
.A2(n_512),
.A3(n_518),
.B(n_506),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_549),
.B(n_552),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_529),
.A2(n_499),
.B1(n_501),
.B2(n_502),
.Y(n_551)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_551),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_529),
.A2(n_522),
.B1(n_518),
.B2(n_355),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_531),
.B(n_501),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_553),
.B(n_539),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_536),
.B(n_519),
.C(n_503),
.Y(n_554)
);

NOR2xp67_ASAP7_75t_SL g560 ( 
.A(n_554),
.B(n_533),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_555),
.B(n_542),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_541),
.B(n_503),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_560),
.A2(n_564),
.B(n_569),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_535),
.C(n_525),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_563),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_526),
.C(n_523),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_527),
.C(n_528),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_566),
.B(n_571),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_568),
.B(n_557),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_544),
.B(n_527),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_561),
.A2(n_558),
.B(n_544),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g581 ( 
.A1(n_573),
.A2(n_576),
.B(n_557),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_567),
.A2(n_545),
.B1(n_564),
.B2(n_570),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_574),
.B(n_575),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_565),
.A2(n_558),
.B(n_554),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_565),
.A2(n_545),
.B1(n_548),
.B2(n_551),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_578),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_581),
.B(n_582),
.Y(n_586)
);

OAI321xp33_ASAP7_75t_L g582 ( 
.A1(n_579),
.A2(n_548),
.A3(n_528),
.B1(n_532),
.B2(n_568),
.C(n_555),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_577),
.B(n_543),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_584),
.B(n_579),
.Y(n_585)
);

AOI21x1_ASAP7_75t_SL g588 ( 
.A1(n_585),
.A2(n_572),
.B(n_583),
.Y(n_588)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_580),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_587),
.B(n_547),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_588),
.A2(n_589),
.B(n_586),
.Y(n_590)
);

AOI321xp33_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_378),
.A3(n_559),
.B1(n_541),
.B2(n_324),
.C(n_281),
.Y(n_591)
);

OAI211xp5_ASAP7_75t_SL g592 ( 
.A1(n_591),
.A2(n_255),
.B(n_264),
.C(n_275),
.Y(n_592)
);

OAI321xp33_ASAP7_75t_L g593 ( 
.A1(n_592),
.A2(n_264),
.A3(n_271),
.B1(n_294),
.B2(n_586),
.C(n_477),
.Y(n_593)
);


endmodule