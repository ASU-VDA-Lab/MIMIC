module fake_netlist_6_1040_n_3858 (n_52, n_591, n_435, n_1, n_91, n_793, n_326, n_801, n_256, n_440, n_587, n_695, n_507, n_580, n_762, n_209, n_367, n_465, n_680, n_741, n_760, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_726, n_316, n_419, n_28, n_304, n_212, n_700, n_50, n_694, n_7, n_740, n_578, n_703, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_783, n_106, n_725, n_358, n_160, n_751, n_449, n_131, n_749, n_798, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_677, n_805, n_396, n_495, n_815, n_350, n_78, n_84, n_585, n_732, n_568, n_392, n_442, n_480, n_142, n_724, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_698, n_255, n_807, n_739, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_768, n_38, n_471, n_289, n_421, n_781, n_424, n_789, n_615, n_59, n_181, n_182, n_238, n_573, n_769, n_202, n_320, n_108, n_639, n_676, n_327, n_794, n_727, n_369, n_597, n_685, n_280, n_287, n_353, n_610, n_555, n_389, n_814, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_718, n_747, n_667, n_71, n_74, n_229, n_542, n_644, n_682, n_621, n_305, n_72, n_721, n_750, n_532, n_742, n_173, n_535, n_691, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_791, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_704, n_748, n_506, n_56, n_763, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_710, n_387, n_452, n_616, n_658, n_744, n_39, n_344, n_73, n_581, n_428, n_761, n_785, n_746, n_609, n_765, n_432, n_641, n_693, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_720, n_525, n_758, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_772, n_96, n_8, n_797, n_666, n_371, n_795, n_770, n_567, n_189, n_738, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_705, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_684, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_752, n_112, n_172, n_713, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_782, n_490, n_803, n_290, n_220, n_809, n_118, n_224, n_48, n_25, n_93, n_80, n_734, n_708, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_779, n_9, n_800, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_709, n_366, n_777, n_407, n_450, n_103, n_808, n_272, n_526, n_185, n_712, n_348, n_711, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_717, n_46, n_330, n_771, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_699, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_686, n_796, n_252, n_757, n_228, n_565, n_594, n_719, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_813, n_592, n_745, n_654, n_323, n_606, n_393, n_411, n_503, n_716, n_152, n_623, n_92, n_599, n_513, n_776, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_731, n_406, n_483, n_735, n_102, n_204, n_482, n_755, n_474, n_527, n_261, n_608, n_620, n_420, n_683, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_792, n_476, n_714, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_788, n_325, n_767, n_804, n_329, n_464, n_600, n_802, n_561, n_33, n_477, n_549, n_533, n_408, n_806, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_707, n_345, n_409, n_231, n_354, n_689, n_40, n_799, n_505, n_240, n_756, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_810, n_635, n_95, n_787, n_311, n_10, n_403, n_723, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_764, n_556, n_159, n_157, n_162, n_692, n_733, n_754, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_753, n_642, n_276, n_569, n_441, n_221, n_811, n_444, n_586, n_423, n_146, n_737, n_318, n_303, n_511, n_715, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_790, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_775, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_679, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_759, n_355, n_426, n_317, n_149, n_632, n_702, n_431, n_90, n_347, n_812, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_780, n_773, n_675, n_85, n_99, n_257, n_730, n_655, n_13, n_706, n_786, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_690, n_29, n_75, n_401, n_324, n_743, n_766, n_816, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_728, n_681, n_729, n_110, n_151, n_774, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_784, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_696, n_688, n_722, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_687, n_697, n_364, n_637, n_295, n_385, n_701, n_817, n_629, n_388, n_190, n_262, n_484, n_613, n_736, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_778, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_678, n_192, n_57, n_169, n_51, n_649, n_283, n_3858);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_793;
input n_326;
input n_801;
input n_256;
input n_440;
input n_587;
input n_695;
input n_507;
input n_580;
input n_762;
input n_209;
input n_367;
input n_465;
input n_680;
input n_741;
input n_760;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_726;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_700;
input n_50;
input n_694;
input n_7;
input n_740;
input n_578;
input n_703;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_783;
input n_106;
input n_725;
input n_358;
input n_160;
input n_751;
input n_449;
input n_131;
input n_749;
input n_798;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_677;
input n_805;
input n_396;
input n_495;
input n_815;
input n_350;
input n_78;
input n_84;
input n_585;
input n_732;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_724;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_698;
input n_255;
input n_807;
input n_739;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_768;
input n_38;
input n_471;
input n_289;
input n_421;
input n_781;
input n_424;
input n_789;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_769;
input n_202;
input n_320;
input n_108;
input n_639;
input n_676;
input n_327;
input n_794;
input n_727;
input n_369;
input n_597;
input n_685;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_814;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_718;
input n_747;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_682;
input n_621;
input n_305;
input n_72;
input n_721;
input n_750;
input n_532;
input n_742;
input n_173;
input n_535;
input n_691;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_791;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_704;
input n_748;
input n_506;
input n_56;
input n_763;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_710;
input n_387;
input n_452;
input n_616;
input n_658;
input n_744;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_761;
input n_785;
input n_746;
input n_609;
input n_765;
input n_432;
input n_641;
input n_693;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_720;
input n_525;
input n_758;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_772;
input n_96;
input n_8;
input n_797;
input n_666;
input n_371;
input n_795;
input n_770;
input n_567;
input n_189;
input n_738;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_705;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_684;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_752;
input n_112;
input n_172;
input n_713;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_782;
input n_490;
input n_803;
input n_290;
input n_220;
input n_809;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_734;
input n_708;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_779;
input n_9;
input n_800;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_709;
input n_366;
input n_777;
input n_407;
input n_450;
input n_103;
input n_808;
input n_272;
input n_526;
input n_185;
input n_712;
input n_348;
input n_711;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_717;
input n_46;
input n_330;
input n_771;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_699;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_686;
input n_796;
input n_252;
input n_757;
input n_228;
input n_565;
input n_594;
input n_719;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_813;
input n_592;
input n_745;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_716;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_776;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_731;
input n_406;
input n_483;
input n_735;
input n_102;
input n_204;
input n_482;
input n_755;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_683;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_792;
input n_476;
input n_714;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_788;
input n_325;
input n_767;
input n_804;
input n_329;
input n_464;
input n_600;
input n_802;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_806;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_707;
input n_345;
input n_409;
input n_231;
input n_354;
input n_689;
input n_40;
input n_799;
input n_505;
input n_240;
input n_756;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_810;
input n_635;
input n_95;
input n_787;
input n_311;
input n_10;
input n_403;
input n_723;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_764;
input n_556;
input n_159;
input n_157;
input n_162;
input n_692;
input n_733;
input n_754;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_753;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_811;
input n_444;
input n_586;
input n_423;
input n_146;
input n_737;
input n_318;
input n_303;
input n_511;
input n_715;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_790;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_775;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_679;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_759;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_702;
input n_431;
input n_90;
input n_347;
input n_812;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_780;
input n_773;
input n_675;
input n_85;
input n_99;
input n_257;
input n_730;
input n_655;
input n_13;
input n_706;
input n_786;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_690;
input n_29;
input n_75;
input n_401;
input n_324;
input n_743;
input n_766;
input n_816;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_728;
input n_681;
input n_729;
input n_110;
input n_151;
input n_774;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_784;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_696;
input n_688;
input n_722;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_687;
input n_697;
input n_364;
input n_637;
input n_295;
input n_385;
input n_701;
input n_817;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_736;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_778;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_678;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_3858;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1674;
wire n_1199;
wire n_3392;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_1189;
wire n_3152;
wire n_3579;
wire n_1212;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3773;
wire n_3783;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_1357;
wire n_1853;
wire n_3741;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_2324;
wire n_1854;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_1708;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_3465;
wire n_1975;
wire n_1743;
wire n_1930;
wire n_1009;
wire n_2405;
wire n_3706;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_1264;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_1371;
wire n_873;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_1985;
wire n_2989;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_2247;
wire n_1711;
wire n_1078;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_3345;
wire n_2074;
wire n_2447;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_2356;
wire n_1143;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_2480;
wire n_1300;
wire n_2739;
wire n_3023;
wire n_822;
wire n_3232;
wire n_2791;
wire n_1313;
wire n_3750;
wire n_3607;
wire n_3251;
wire n_1056;
wire n_3316;
wire n_2212;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_940;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_3765;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_1467;
wire n_3297;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_1088;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3368;
wire n_917;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_1446;
wire n_2591;
wire n_3507;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_913;
wire n_1658;
wire n_2593;
wire n_867;
wire n_3506;
wire n_3568;
wire n_3269;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_1967;
wire n_1193;
wire n_1054;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_1986;
wire n_2397;
wire n_824;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_2907;
wire n_3438;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1599;
wire n_1068;
wire n_3732;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_3446;
wire n_3317;
wire n_3857;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_3716;
wire n_1873;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_3842;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1605;
wire n_1330;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_2355;
wire n_966;
wire n_2908;
wire n_3168;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_3403;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_1233;
wire n_2714;
wire n_1289;
wire n_2245;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_1014;
wire n_3734;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_1265;
wire n_2711;
wire n_3490;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_2878;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_3247;
wire n_871;
wire n_3069;
wire n_922;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1722;
wire n_1664;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_1801;
wire n_835;
wire n_928;
wire n_2347;
wire n_850;
wire n_1214;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3428;
wire n_3153;
wire n_3410;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_1588;
wire n_3785;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_1624;
wire n_1124;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_3434;
wire n_1515;
wire n_961;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_890;
wire n_2377;
wire n_3271;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_3545;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_1767;
wire n_3253;
wire n_1779;
wire n_1465;
wire n_3337;
wire n_3431;
wire n_3209;
wire n_3450;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_2493;
wire n_1128;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1565;
wire n_1067;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_3616;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_2693;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_963;
wire n_2767;
wire n_3793;
wire n_894;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1714;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3171;
wire n_1913;
wire n_3608;
wire n_837;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_3491;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_1432;
wire n_2208;
wire n_843;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_2134;
wire n_1176;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_2539;
wire n_2698;
wire n_2667;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_947;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1448;
wire n_1087;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_1049;
wire n_3223;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_1717;
wire n_1817;
wire n_926;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_1299;
wire n_2896;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_998;
wire n_3200;
wire n_1665;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_3390;
wire n_3656;
wire n_1178;
wire n_2127;
wire n_2338;
wire n_1424;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_1073;
wire n_1000;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_1507;
wire n_2482;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_1398;
wire n_2354;
wire n_884;
wire n_1048;
wire n_2682;
wire n_1201;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_1021;
wire n_931;
wire n_3393;
wire n_2442;
wire n_1207;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3480;
wire n_3451;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_3591;
wire n_3641;
wire n_1314;
wire n_1837;
wire n_831;
wire n_964;
wire n_2218;
wire n_2788;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2860;
wire n_2292;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_3481;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_2990;
wire n_3847;
wire n_1775;
wire n_1773;
wire n_1286;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3226;
wire n_3323;
wire n_3364;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_3425;
wire n_2384;
wire n_1745;
wire n_914;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_2920;
wire n_3547;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_1617;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_1470;
wire n_2550;
wire n_3093;
wire n_3175;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_2249;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_1390;
wire n_906;
wire n_2289;
wire n_1733;
wire n_2315;
wire n_1077;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_2627;
wire n_3234;
wire n_956;
wire n_960;
wire n_2276;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_1129;
wire n_2829;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_3751;
wire n_1869;
wire n_3625;
wire n_2911;
wire n_3804;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_3338;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_2984;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3276;
wire n_3250;
wire n_1934;
wire n_3194;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_845;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_1510;
wire n_892;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_1667;
wire n_1206;
wire n_3230;
wire n_1397;
wire n_1037;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_1499;
wire n_901;
wire n_3592;
wire n_2755;
wire n_3141;
wire n_923;
wire n_1409;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_3195;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_2439;
wire n_1818;
wire n_1108;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_2740;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1943;
wire n_1216;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_3784;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_3594;
wire n_1043;
wire n_3819;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_3485;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_3501;
wire n_1840;
wire n_1152;
wire n_1705;
wire n_3262;
wire n_3544;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_3790;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_3320;
wire n_2541;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_1637;
wire n_934;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_2871;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_2390;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_2986;
wire n_1900;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_2962;
wire n_2727;
wire n_2154;
wire n_3377;
wire n_2939;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_1706;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_3156;
wire n_2083;
wire n_1931;
wire n_1269;
wire n_2834;
wire n_3207;
wire n_2668;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_2128;
wire n_1650;
wire n_1794;
wire n_1962;
wire n_1045;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_3818;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1002;
wire n_1325;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_3524;
wire n_2671;
wire n_2761;
wire n_2885;
wire n_2793;
wire n_2715;
wire n_2888;
wire n_1804;
wire n_2923;
wire n_3711;
wire n_3776;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_3511;
wire n_2054;
wire n_876;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1600;
wire n_1113;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_2261;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_1476;
wire n_841;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_3808;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1882;
wire n_1023;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1929;
wire n_1007;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_3806;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_2400;
wire n_1716;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_3565;
wire n_1953;
wire n_933;
wire n_3343;
wire n_3303;
wire n_978;
wire n_2752;
wire n_3135;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_1074;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_1554;
wire n_3231;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_2380;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_2290;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_3541;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_1461;
wire n_3432;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_1598;
wire n_3493;
wire n_2935;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_2385;
wire n_1283;
wire n_918;
wire n_1785;
wire n_1848;
wire n_1114;
wire n_1147;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_1994;
wire n_957;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_971;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_2769;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3336;
wire n_844;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_3553;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_2465;
wire n_1112;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_3584;
wire n_3486;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_3556;
wire n_2034;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_2444;
wire n_2437;
wire n_1215;
wire n_839;
wire n_2743;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_990;
wire n_1500;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_2312;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_1509;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_2609;
wire n_1161;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_1584;
wire n_2425;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_3680;
wire n_2318;
wire n_3286;
wire n_2408;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1362;
wire n_1156;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_859;
wire n_3086;
wire n_2033;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_3285;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_3478;
wire n_1349;
wire n_2071;
wire n_1144;
wire n_3669;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_3344;
wire n_2334;
wire n_3295;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_1133;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_2367;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_3187;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_2968;
wire n_1629;
wire n_2221;
wire n_1170;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_2553;
wire n_1040;
wire n_915;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_3815;
wire n_2774;
wire n_3039;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3274;
wire n_3333;
wire n_3186;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_2579;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3387;
wire n_2027;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_3504;
wire n_1449;
wire n_827;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_191),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_283),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_371),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_61),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_794),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_318),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_277),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_716),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_256),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_495),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_194),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_600),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_506),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_811),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_97),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_506),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_83),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_756),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_422),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_429),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_384),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_100),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_737),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_417),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_752),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_724),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_430),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_16),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_167),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_230),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_148),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_566),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_440),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_377),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_632),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_760),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_792),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_765),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_595),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_60),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_390),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_698),
.Y(n_859)
);

CKINVDCx14_ASAP7_75t_R g860 ( 
.A(n_774),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_537),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_304),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_398),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_800),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_665),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_677),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_557),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_631),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_646),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_646),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_536),
.Y(n_871)
);

BUFx5_ASAP7_75t_L g872 ( 
.A(n_723),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_164),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_24),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_747),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_393),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_685),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_325),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_719),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_745),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_775),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_734),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_451),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_138),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_445),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_815),
.Y(n_886)
);

BUFx10_ASAP7_75t_L g887 ( 
.A(n_207),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_753),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_421),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_492),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_451),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_394),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_753),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_485),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_457),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_298),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_284),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_227),
.Y(n_898)
);

CKINVDCx16_ASAP7_75t_R g899 ( 
.A(n_736),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_699),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_513),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_432),
.Y(n_902)
);

CKINVDCx14_ASAP7_75t_R g903 ( 
.A(n_341),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_807),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_91),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_720),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_232),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_124),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_462),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_78),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_66),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_699),
.Y(n_912)
);

CKINVDCx20_ASAP7_75t_R g913 ( 
.A(n_722),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_633),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_686),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_38),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_66),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_767),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_770),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_369),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_161),
.Y(n_921)
);

BUFx5_ASAP7_75t_L g922 ( 
.A(n_210),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_763),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_444),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_695),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_435),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_784),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_710),
.Y(n_928)
);

BUFx3_ASAP7_75t_L g929 ( 
.A(n_53),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_137),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_675),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_746),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_113),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_334),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_361),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_228),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_13),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_188),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_32),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_817),
.Y(n_940)
);

BUFx10_ASAP7_75t_L g941 ( 
.A(n_85),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_679),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_669),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_494),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_458),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_133),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_407),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_213),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_593),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_742),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_445),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_809),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_594),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_490),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_369),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_300),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_468),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_597),
.Y(n_958)
);

BUFx2_ASAP7_75t_SL g959 ( 
.A(n_628),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_713),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_731),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_223),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_226),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_341),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_635),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_84),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_127),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_89),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_375),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_331),
.Y(n_970)
);

CKINVDCx16_ASAP7_75t_R g971 ( 
.A(n_197),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_145),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_510),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_18),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_19),
.Y(n_975)
);

CKINVDCx11_ASAP7_75t_R g976 ( 
.A(n_127),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_477),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_567),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_515),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_517),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_697),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_524),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_377),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_101),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_393),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_580),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_80),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_540),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_412),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_755),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_689),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_751),
.Y(n_992)
);

BUFx2_ASAP7_75t_SL g993 ( 
.A(n_739),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_117),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_266),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_762),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_408),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_801),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_185),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_21),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_213),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_744),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_356),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_669),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_189),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_406),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_523),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_123),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_346),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_743),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_740),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_726),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_327),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_375),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_707),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_554),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_557),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_165),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_730),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_115),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_804),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_630),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_675),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_119),
.Y(n_1024)
);

CKINVDCx14_ASAP7_75t_R g1025 ( 
.A(n_298),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_609),
.Y(n_1026)
);

BUFx10_ASAP7_75t_L g1027 ( 
.A(n_159),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_319),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_791),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_782),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_25),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_759),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_648),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_771),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_616),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_339),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_333),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_785),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_567),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_120),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_814),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_812),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_SL g1043 ( 
.A(n_106),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_137),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_767),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_511),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_746),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_96),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_155),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_563),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_772),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_780),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_325),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_520),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_751),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_411),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_722),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_229),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_614),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_354),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_657),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_706),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_714),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_108),
.Y(n_1064)
);

BUFx10_ASAP7_75t_L g1065 ( 
.A(n_715),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_16),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_269),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_219),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_209),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_143),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_601),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_765),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_43),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_587),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_476),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_132),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_769),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_766),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_49),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_589),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_424),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_303),
.Y(n_1082)
);

BUFx10_ASAP7_75t_L g1083 ( 
.A(n_386),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_59),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_135),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_647),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_718),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_490),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_631),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_240),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_790),
.Y(n_1091)
);

BUFx3_ASAP7_75t_L g1092 ( 
.A(n_709),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_584),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_233),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_243),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_768),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_540),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_175),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_790),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_719),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_521),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_518),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_600),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_773),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_431),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_229),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_418),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_729),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_563),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_542),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_517),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_615),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_710),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_49),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_172),
.Y(n_1115)
);

CKINVDCx16_ASAP7_75t_R g1116 ( 
.A(n_209),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_165),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_593),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_725),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_394),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_35),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_378),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_314),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_331),
.Y(n_1124)
);

CKINVDCx14_ASAP7_75t_R g1125 ( 
.A(n_56),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_374),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_507),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_381),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_735),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_74),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_511),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_706),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_526),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_327),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_440),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_712),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_579),
.Y(n_1137)
);

INVx1_ASAP7_75t_SL g1138 ( 
.A(n_771),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_176),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_439),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_448),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_456),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_748),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_522),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_744),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_750),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_266),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_573),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_749),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_113),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_8),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_317),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_153),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_337),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_214),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_575),
.Y(n_1156)
);

BUFx3_ASAP7_75t_L g1157 ( 
.A(n_55),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_426),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_285),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_741),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_499),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_518),
.Y(n_1162)
);

CKINVDCx16_ASAP7_75t_R g1163 ( 
.A(n_606),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_373),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_212),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_816),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_475),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_462),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_677),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_115),
.Y(n_1170)
);

CKINVDCx12_ASAP7_75t_R g1171 ( 
.A(n_539),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_648),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_756),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_520),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_768),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_90),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_577),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_808),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_147),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_336),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_123),
.Y(n_1181)
);

BUFx5_ASAP7_75t_L g1182 ( 
.A(n_491),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_78),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_776),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_92),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_181),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_140),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_207),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_592),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_204),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_141),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_398),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_234),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_48),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_688),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_455),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_482),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_778),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_653),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_378),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_438),
.Y(n_1201)
);

BUFx5_ASAP7_75t_L g1202 ( 
.A(n_566),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_592),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_120),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_296),
.Y(n_1205)
);

BUFx10_ASAP7_75t_L g1206 ( 
.A(n_736),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_596),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_795),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_758),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_466),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_470),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_264),
.Y(n_1212)
);

BUFx10_ASAP7_75t_L g1213 ( 
.A(n_288),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_426),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_32),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_732),
.Y(n_1216)
);

BUFx10_ASAP7_75t_L g1217 ( 
.A(n_57),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_702),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_573),
.Y(n_1219)
);

INVx1_ASAP7_75t_SL g1220 ( 
.A(n_621),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_537),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_343),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_673),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_747),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_430),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_574),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_721),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_734),
.Y(n_1228)
);

BUFx10_ASAP7_75t_L g1229 ( 
.A(n_764),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_174),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_743),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_615),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_68),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_627),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_247),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_524),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_272),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_217),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_489),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_190),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_386),
.Y(n_1241)
);

BUFx2_ASAP7_75t_SL g1242 ( 
.A(n_246),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_485),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_114),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_376),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_576),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_791),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_118),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_725),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_366),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_277),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_217),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_502),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_105),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_659),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_268),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_397),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_528),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_89),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_145),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_203),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_754),
.Y(n_1262)
);

CKINVDCx16_ASAP7_75t_R g1263 ( 
.A(n_190),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_152),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_212),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_218),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_423),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_326),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_616),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_333),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_638),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_783),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_531),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_544),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_636),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_138),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_740),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_22),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_255),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_301),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_387),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_29),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_738),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_806),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_770),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_569),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_456),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_272),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_733),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_625),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_536),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_187),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_561),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_680),
.Y(n_1294)
);

CKINVDCx16_ASAP7_75t_R g1295 ( 
.A(n_314),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_612),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_111),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_531),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_361),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_72),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_813),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_17),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_417),
.Y(n_1303)
);

CKINVDCx20_ASAP7_75t_R g1304 ( 
.A(n_263),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_47),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_608),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_561),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_200),
.Y(n_1308)
);

CKINVDCx16_ASAP7_75t_R g1309 ( 
.A(n_432),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_465),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_810),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_264),
.Y(n_1312)
);

CKINVDCx16_ASAP7_75t_R g1313 ( 
.A(n_727),
.Y(n_1313)
);

BUFx6f_ASAP7_75t_L g1314 ( 
.A(n_488),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_533),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_643),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_559),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_406),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_726),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_779),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_708),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_43),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_711),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_554),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_795),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_763),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_460),
.Y(n_1327)
);

INVxp67_ASAP7_75t_L g1328 ( 
.A(n_569),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_141),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_352),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_348),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_460),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_709),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_728),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_238),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_647),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_175),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_303),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_59),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_623),
.Y(n_1340)
);

CKINVDCx20_ASAP7_75t_R g1341 ( 
.A(n_688),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_781),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_332),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_25),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_122),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_366),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_708),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_160),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_757),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_103),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_104),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_415),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_761),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_446),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_717),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_441),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_777),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_847),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_872),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_860),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_903),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1025),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_976),
.Y(n_1363)
);

INVxp33_ASAP7_75t_L g1364 ( 
.A(n_1063),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_872),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_872),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_872),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_831),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_872),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_872),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_872),
.Y(n_1371)
);

NOR2xp67_ASAP7_75t_L g1372 ( 
.A(n_1222),
.B(n_0),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_952),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_922),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_922),
.Y(n_1375)
);

INVxp33_ASAP7_75t_SL g1376 ( 
.A(n_1069),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1222),
.B(n_0),
.Y(n_1377)
);

INVxp33_ASAP7_75t_SL g1378 ( 
.A(n_1260),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_922),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_922),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1301),
.Y(n_1381)
);

INVxp33_ASAP7_75t_SL g1382 ( 
.A(n_821),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_847),
.Y(n_1383)
);

INVxp67_ASAP7_75t_L g1384 ( 
.A(n_992),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_922),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_922),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_922),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1182),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1182),
.Y(n_1389)
);

CKINVDCx16_ASAP7_75t_R g1390 ( 
.A(n_838),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1182),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1182),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1182),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1110),
.Y(n_1394)
);

INVxp33_ASAP7_75t_SL g1395 ( 
.A(n_1349),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1182),
.Y(n_1396)
);

INVx3_ASAP7_75t_L g1397 ( 
.A(n_834),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1182),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1125),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1222),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1202),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1021),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_865),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1202),
.Y(n_1404)
);

INVxp33_ASAP7_75t_L g1405 ( 
.A(n_1203),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_818),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1202),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1202),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_865),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1202),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1166),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1232),
.Y(n_1412)
);

INVxp33_ASAP7_75t_SL g1413 ( 
.A(n_1353),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1202),
.Y(n_1414)
);

INVxp33_ASAP7_75t_L g1415 ( 
.A(n_1043),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1202),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1232),
.B(n_1),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1232),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_867),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1073),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_867),
.Y(n_1421)
);

CKINVDCx16_ASAP7_75t_R g1422 ( 
.A(n_899),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_929),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_929),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_932),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1178),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_834),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_932),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_L g1429 ( 
.A(n_897),
.B(n_1),
.Y(n_1429)
);

CKINVDCx16_ASAP7_75t_R g1430 ( 
.A(n_971),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_965),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_965),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_968),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_968),
.Y(n_1434)
);

CKINVDCx16_ASAP7_75t_R g1435 ( 
.A(n_1116),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1033),
.Y(n_1436)
);

CKINVDCx16_ASAP7_75t_R g1437 ( 
.A(n_1142),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1033),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1073),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_818),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1092),
.Y(n_1441)
);

INVxp33_ASAP7_75t_L g1442 ( 
.A(n_840),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1092),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_859),
.Y(n_1444)
);

INVxp67_ASAP7_75t_SL g1445 ( 
.A(n_834),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_834),
.B(n_2),
.Y(n_1446)
);

INVxp33_ASAP7_75t_SL g1447 ( 
.A(n_821),
.Y(n_1447)
);

INVxp33_ASAP7_75t_SL g1448 ( 
.A(n_822),
.Y(n_1448)
);

CKINVDCx16_ASAP7_75t_R g1449 ( 
.A(n_1163),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1126),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1126),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1134),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_834),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1284),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1134),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1157),
.Y(n_1456)
);

CKINVDCx16_ASAP7_75t_R g1457 ( 
.A(n_1263),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1157),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1164),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1285),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1164),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1219),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1219),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1231),
.Y(n_1464)
);

INVxp33_ASAP7_75t_L g1465 ( 
.A(n_840),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_904),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1231),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_864),
.Y(n_1468)
);

INVxp67_ASAP7_75t_SL g1469 ( 
.A(n_939),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_859),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1234),
.Y(n_1471)
);

CKINVDCx16_ASAP7_75t_R g1472 ( 
.A(n_1295),
.Y(n_1472)
);

CKINVDCx16_ASAP7_75t_R g1473 ( 
.A(n_1309),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1234),
.Y(n_1474)
);

CKINVDCx16_ASAP7_75t_R g1475 ( 
.A(n_1313),
.Y(n_1475)
);

INVxp67_ASAP7_75t_SL g1476 ( 
.A(n_939),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_939),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1274),
.Y(n_1478)
);

CKINVDCx16_ASAP7_75t_R g1479 ( 
.A(n_859),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_824),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_939),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1274),
.Y(n_1482)
);

CKINVDCx16_ASAP7_75t_R g1483 ( 
.A(n_887),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_939),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1004),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1004),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1004),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1004),
.Y(n_1488)
);

CKINVDCx14_ASAP7_75t_R g1489 ( 
.A(n_864),
.Y(n_1489)
);

INVxp67_ASAP7_75t_SL g1490 ( 
.A(n_1004),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1053),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1053),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1053),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_940),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_825),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1053),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1359),
.A2(n_1042),
.B(n_1041),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1406),
.A2(n_827),
.B1(n_853),
.B2(n_832),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1427),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1445),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1460),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1453),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1397),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1381),
.B(n_1311),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1477),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1477),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_SL g1507 ( 
.A(n_1360),
.B(n_827),
.Y(n_1507)
);

CKINVDCx20_ASAP7_75t_R g1508 ( 
.A(n_1411),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1481),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1376),
.A2(n_1070),
.B1(n_826),
.B2(n_829),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1397),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_1381),
.B(n_1140),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1481),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1469),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1484),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1485),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1486),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1487),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1476),
.Y(n_1519)
);

INVx5_ASAP7_75t_L g1520 ( 
.A(n_1458),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1378),
.A2(n_828),
.B1(n_839),
.B2(n_836),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1368),
.B(n_886),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1488),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_1373),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1454),
.Y(n_1526)
);

AND2x6_ASAP7_75t_L g1527 ( 
.A(n_1365),
.B(n_998),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_SL g1528 ( 
.A(n_1361),
.B(n_832),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1496),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1400),
.B(n_1140),
.Y(n_1530)
);

BUFx6f_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1492),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1412),
.B(n_1160),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1493),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1466),
.Y(n_1535)
);

AND2x2_ASAP7_75t_SL g1536 ( 
.A(n_1390),
.B(n_1053),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1466),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1366),
.A2(n_868),
.B(n_845),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1419),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1415),
.B(n_887),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_SL g1541 ( 
.A1(n_1406),
.A2(n_854),
.B1(n_862),
.B2(n_853),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1362),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1418),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1384),
.B(n_1160),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1388),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1394),
.B(n_1272),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1402),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1388),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1421),
.Y(n_1549)
);

INVx5_ASAP7_75t_L g1550 ( 
.A(n_1479),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1423),
.B(n_1272),
.Y(n_1551)
);

AND2x6_ASAP7_75t_L g1552 ( 
.A(n_1367),
.B(n_998),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1369),
.Y(n_1553)
);

AND2x2_ASAP7_75t_SL g1554 ( 
.A(n_1422),
.B(n_1154),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1424),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1494),
.Y(n_1556)
);

BUFx6f_ASAP7_75t_L g1557 ( 
.A(n_1494),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1480),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1425),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1363),
.Y(n_1560)
);

BUFx8_ASAP7_75t_SL g1561 ( 
.A(n_1440),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1370),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1428),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1371),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1374),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1431),
.B(n_1343),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1495),
.Y(n_1567)
);

AOI22x1_ASAP7_75t_SL g1568 ( 
.A1(n_1440),
.A2(n_862),
.B1(n_879),
.B2(n_854),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1375),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1426),
.B(n_886),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1358),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1399),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1430),
.A2(n_842),
.B1(n_844),
.B2(n_843),
.Y(n_1573)
);

BUFx12f_ASAP7_75t_L g1574 ( 
.A(n_1435),
.Y(n_1574)
);

OAI22xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1415),
.A2(n_896),
.B1(n_913),
.B2(n_879),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_SL g1576 ( 
.A1(n_1468),
.A2(n_913),
.B1(n_918),
.B2(n_896),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_1379),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1437),
.B(n_1154),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1444),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1380),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1489),
.B(n_887),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1385),
.Y(n_1582)
);

CKINVDCx8_ASAP7_75t_R g1583 ( 
.A(n_1449),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1432),
.B(n_1343),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1433),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1489),
.B(n_941),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1434),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1405),
.A2(n_1328),
.B1(n_1266),
.B2(n_848),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1382),
.B(n_1154),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1386),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1387),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1436),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1389),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1358),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1457),
.Y(n_1595)
);

BUFx8_ASAP7_75t_L g1596 ( 
.A(n_1438),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1483),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1441),
.B(n_1154),
.Y(n_1598)
);

INVx4_ASAP7_75t_SL g1599 ( 
.A(n_1443),
.Y(n_1599)
);

BUFx3_ASAP7_75t_L g1600 ( 
.A(n_1450),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_SL g1601 ( 
.A(n_1472),
.B(n_1154),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1451),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_1391),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1482),
.Y(n_1604)
);

INVx4_ASAP7_75t_L g1605 ( 
.A(n_1392),
.Y(n_1605)
);

BUFx6f_ASAP7_75t_L g1606 ( 
.A(n_1393),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1396),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1452),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1455),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1456),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1459),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1470),
.Y(n_1612)
);

BUFx2_ASAP7_75t_L g1613 ( 
.A(n_1383),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1461),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1462),
.B(n_1314),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1405),
.A2(n_1364),
.B1(n_1413),
.B2(n_1395),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1398),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1401),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1478),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1463),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1383),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1549),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1553),
.B(n_1404),
.Y(n_1623)
);

AOI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1588),
.A2(n_918),
.B1(n_935),
.B2(n_927),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_SL g1625 ( 
.A(n_1536),
.B(n_1473),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1555),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1509),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1559),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1509),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1509),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1540),
.B(n_1475),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1564),
.B(n_1407),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1516),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1516),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1613),
.B(n_1442),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1554),
.A2(n_935),
.B1(n_960),
.B2(n_927),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1516),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1517),
.Y(n_1639)
);

OA21x2_ASAP7_75t_L g1640 ( 
.A1(n_1565),
.A2(n_1607),
.B(n_1582),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1587),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1592),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1604),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1614),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1517),
.Y(n_1645)
);

BUFx8_ASAP7_75t_L g1646 ( 
.A(n_1574),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1619),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_1556),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_R g1649 ( 
.A1(n_1568),
.A2(n_1318),
.B1(n_1233),
.B2(n_925),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1497),
.A2(n_1410),
.B(n_1408),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1599),
.B(n_1464),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1556),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1613),
.B(n_1442),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1517),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1620),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1535),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1518),
.Y(n_1657)
);

BUFx8_ASAP7_75t_L g1658 ( 
.A(n_1560),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1499),
.B(n_1447),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1465),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1498),
.A2(n_972),
.B1(n_986),
.B2(n_960),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1621),
.B(n_1465),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1595),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1571),
.B(n_1364),
.Y(n_1664)
);

BUFx6f_ASAP7_75t_L g1665 ( 
.A(n_1556),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1518),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1557),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1522),
.B(n_1448),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1594),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1599),
.B(n_1467),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1524),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1512),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1562),
.Y(n_1673)
);

BUFx3_ASAP7_75t_L g1674 ( 
.A(n_1535),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1562),
.Y(n_1675)
);

INVx3_ASAP7_75t_L g1676 ( 
.A(n_1518),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1531),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1562),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1531),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1569),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1557),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1569),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1531),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1581),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1532),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1520),
.B(n_1586),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1569),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1537),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1577),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1577),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1532),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1497),
.A2(n_1416),
.B(n_1414),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1532),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1577),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1617),
.B(n_1377),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1580),
.Y(n_1696)
);

AOI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1510),
.A2(n_986),
.B1(n_1059),
.B2(n_972),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1545),
.B(n_1377),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1538),
.A2(n_1417),
.B(n_1372),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1505),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1580),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1512),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1579),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1580),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1557),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1537),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1506),
.Y(n_1707)
);

INVx6_ASAP7_75t_L g1708 ( 
.A(n_1520),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1520),
.B(n_1403),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1590),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1548),
.B(n_1446),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1590),
.Y(n_1712)
);

INVx5_ASAP7_75t_L g1713 ( 
.A(n_1527),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1590),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1550),
.B(n_1429),
.Y(n_1715)
);

BUFx6f_ASAP7_75t_L g1716 ( 
.A(n_1591),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1550),
.B(n_941),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1570),
.B(n_1471),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1591),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1591),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1547),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1579),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1593),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1503),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1500),
.B(n_1474),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1605),
.B(n_1446),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1539),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1593),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1513),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1511),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1593),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1603),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1600),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1515),
.Y(n_1734)
);

BUFx2_ASAP7_75t_L g1735 ( 
.A(n_1572),
.Y(n_1735)
);

AND2x4_ASAP7_75t_L g1736 ( 
.A(n_1598),
.B(n_819),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1608),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1603),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1603),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1523),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1605),
.B(n_998),
.Y(n_1741)
);

HB1xp67_ASAP7_75t_L g1742 ( 
.A(n_1598),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1612),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1606),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1606),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1538),
.B(n_1326),
.C(n_1314),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1606),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1534),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_SL g1749 ( 
.A(n_1550),
.B(n_941),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1618),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1618),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1618),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1543),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1615),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1502),
.Y(n_1755)
);

AND2x6_ASAP7_75t_L g1756 ( 
.A(n_1589),
.B(n_998),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1706),
.B(n_1567),
.Y(n_1757)
);

AO22x2_ASAP7_75t_L g1758 ( 
.A1(n_1703),
.A2(n_1568),
.B1(n_1616),
.B2(n_1546),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1636),
.Y(n_1759)
);

INVx2_ASAP7_75t_SL g1760 ( 
.A(n_1653),
.Y(n_1760)
);

INVx4_ASAP7_75t_L g1761 ( 
.A(n_1648),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1668),
.A2(n_1514),
.B1(n_1525),
.B2(n_1519),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1718),
.B(n_1726),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1648),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1640),
.Y(n_1765)
);

NOR2x1p5_ASAP7_75t_L g1766 ( 
.A(n_1671),
.B(n_1597),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1640),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1700),
.Y(n_1768)
);

OR2x6_ASAP7_75t_L g1769 ( 
.A(n_1735),
.B(n_1526),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1660),
.Y(n_1770)
);

BUFx6f_ASAP7_75t_L g1771 ( 
.A(n_1706),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1697),
.B(n_1528),
.C(n_1507),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1662),
.B(n_1530),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1707),
.Y(n_1774)
);

INVx1_ASAP7_75t_SL g1775 ( 
.A(n_1703),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1722),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1709),
.B(n_1612),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1726),
.B(n_1695),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1743),
.B(n_1558),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1742),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1695),
.A2(n_1533),
.B1(n_1530),
.B2(n_1529),
.Y(n_1782)
);

NAND2xp33_ASAP7_75t_L g1783 ( 
.A(n_1756),
.B(n_1713),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1754),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1664),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1684),
.B(n_1533),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1729),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1711),
.B(n_1504),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1659),
.B(n_1702),
.C(n_1672),
.Y(n_1789)
);

INVx5_ASAP7_75t_L g1790 ( 
.A(n_1708),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1754),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1672),
.B(n_1702),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1734),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1711),
.B(n_1504),
.Y(n_1794)
);

BUFx3_ASAP7_75t_L g1795 ( 
.A(n_1706),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1740),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1753),
.Y(n_1797)
);

INVx4_ASAP7_75t_L g1798 ( 
.A(n_1648),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1748),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1656),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1724),
.Y(n_1801)
);

INVx2_ASAP7_75t_SL g1802 ( 
.A(n_1727),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1721),
.Y(n_1803)
);

AND3x2_ASAP7_75t_L g1804 ( 
.A(n_1743),
.B(n_1501),
.C(n_1409),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1622),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1724),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1674),
.B(n_1688),
.Y(n_1807)
);

OAI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1637),
.A2(n_1521),
.B1(n_1573),
.B2(n_1578),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1722),
.B(n_1544),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1727),
.Y(n_1810)
);

BUFx3_ASAP7_75t_L g1811 ( 
.A(n_1652),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_SL g1812 ( 
.A(n_1631),
.B(n_1597),
.Y(n_1812)
);

NOR2x1p5_ASAP7_75t_L g1813 ( 
.A(n_1730),
.B(n_822),
.Y(n_1813)
);

BUFx10_ASAP7_75t_L g1814 ( 
.A(n_1659),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1650),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1626),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1628),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1634),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1641),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1642),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1643),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1692),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1623),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1646),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1623),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1669),
.B(n_1542),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1698),
.B(n_1601),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1644),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1647),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1730),
.Y(n_1830)
);

AND2x6_ASAP7_75t_L g1831 ( 
.A(n_1698),
.B(n_998),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1669),
.B(n_1544),
.Y(n_1832)
);

INVx4_ASAP7_75t_L g1833 ( 
.A(n_1652),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1646),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1658),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1627),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1755),
.A2(n_1546),
.B1(n_1615),
.B2(n_993),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1655),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1733),
.Y(n_1839)
);

INVx5_ASAP7_75t_L g1840 ( 
.A(n_1708),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1673),
.B(n_1738),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1733),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1627),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1737),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1652),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1630),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1737),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1630),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1725),
.B(n_1566),
.C(n_1551),
.Y(n_1849)
);

NAND2xp33_ASAP7_75t_L g1850 ( 
.A(n_1756),
.B(n_1527),
.Y(n_1850)
);

INVx3_ASAP7_75t_L g1851 ( 
.A(n_1629),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1725),
.B(n_1563),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1675),
.B(n_1527),
.Y(n_1853)
);

BUFx6f_ASAP7_75t_L g1854 ( 
.A(n_1665),
.Y(n_1854)
);

INVx4_ASAP7_75t_L g1855 ( 
.A(n_1665),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1665),
.B(n_1583),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1625),
.B(n_1508),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1678),
.B(n_1739),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1680),
.A2(n_1566),
.B1(n_1584),
.B2(n_1551),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1744),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1663),
.Y(n_1861)
);

AND2x2_ASAP7_75t_SL g1862 ( 
.A(n_1637),
.B(n_1403),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1682),
.B(n_1552),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1667),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1632),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1687),
.B(n_1552),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1689),
.B(n_1552),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1632),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1690),
.B(n_1602),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1744),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1694),
.B(n_1609),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_1658),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1696),
.B(n_1747),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_SL g1874 ( 
.A1(n_1661),
.A2(n_1245),
.B1(n_1255),
.B2(n_1059),
.Y(n_1874)
);

OR2x6_ASAP7_75t_L g1875 ( 
.A(n_1661),
.B(n_1575),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1635),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1746),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1667),
.B(n_1610),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1697),
.B(n_1624),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1746),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1736),
.B(n_1611),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_SL g1882 ( 
.A(n_1651),
.B(n_1245),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1699),
.Y(n_1883)
);

BUFx8_ASAP7_75t_SL g1884 ( 
.A(n_1667),
.Y(n_1884)
);

INVx4_ASAP7_75t_L g1885 ( 
.A(n_1681),
.Y(n_1885)
);

BUFx10_ASAP7_75t_L g1886 ( 
.A(n_1736),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1741),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1681),
.B(n_1584),
.Y(n_1888)
);

BUFx10_ASAP7_75t_L g1889 ( 
.A(n_1651),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1681),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1670),
.B(n_1409),
.Y(n_1891)
);

BUFx10_ASAP7_75t_L g1892 ( 
.A(n_1670),
.Y(n_1892)
);

INVx4_ASAP7_75t_L g1893 ( 
.A(n_1705),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1741),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1751),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1716),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1705),
.B(n_1596),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1716),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1752),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1633),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1701),
.B(n_1420),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1635),
.Y(n_1902)
);

CKINVDCx5p33_ASAP7_75t_R g1903 ( 
.A(n_1705),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_SL g1904 ( 
.A(n_1716),
.B(n_1719),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1654),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1638),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1639),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1719),
.B(n_1596),
.Y(n_1908)
);

AND2x2_ASAP7_75t_SL g1909 ( 
.A(n_1624),
.B(n_1420),
.Y(n_1909)
);

BUFx6f_ASAP7_75t_L g1910 ( 
.A(n_1719),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1745),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1756),
.A2(n_1242),
.B1(n_959),
.B2(n_1314),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1745),
.B(n_1314),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1645),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1654),
.Y(n_1915)
);

NOR2xp33_ASAP7_75t_L g1916 ( 
.A(n_1763),
.B(n_1576),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1779),
.B(n_1713),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1865),
.A2(n_1756),
.B1(n_1710),
.B2(n_1712),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1768),
.Y(n_1919)
);

AOI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1827),
.A2(n_1704),
.B1(n_1720),
.B2(n_1714),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1868),
.B(n_1723),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1765),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1809),
.B(n_1802),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1775),
.B(n_1541),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1776),
.Y(n_1925)
);

BUFx6f_ASAP7_75t_L g1926 ( 
.A(n_1771),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1832),
.B(n_1686),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1777),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1774),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1823),
.B(n_1728),
.Y(n_1930)
);

CKINVDCx14_ASAP7_75t_R g1931 ( 
.A(n_1803),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1781),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1823),
.B(n_1731),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1825),
.B(n_1732),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1784),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1825),
.B(n_1745),
.Y(n_1936)
);

AOI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1788),
.A2(n_1794),
.B1(n_1808),
.B2(n_1773),
.Y(n_1937)
);

AND2x4_ASAP7_75t_SL g1938 ( 
.A(n_1889),
.B(n_1750),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1852),
.B(n_1750),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1759),
.A2(n_1657),
.B1(n_1679),
.B2(n_1677),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1887),
.B(n_1750),
.Y(n_1941)
);

INVxp67_ASAP7_75t_SL g1942 ( 
.A(n_1910),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1887),
.B(n_1666),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1780),
.B(n_1561),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1787),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1894),
.B(n_1666),
.Y(n_1946)
);

A2O1A1Ixp33_ASAP7_75t_L g1947 ( 
.A1(n_1849),
.A2(n_1717),
.B(n_1749),
.C(n_1715),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1782),
.B(n_1676),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1816),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1861),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1884),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1810),
.B(n_1713),
.Y(n_1952)
);

BUFx4_ASAP7_75t_L g1953 ( 
.A(n_1839),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1778),
.B(n_1439),
.Y(n_1954)
);

AOI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1909),
.A2(n_1691),
.B1(n_1685),
.B2(n_1683),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1760),
.B(n_1713),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1791),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1770),
.B(n_1439),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1814),
.B(n_1255),
.Y(n_1959)
);

CKINVDCx5p33_ASAP7_75t_R g1960 ( 
.A(n_1769),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1814),
.B(n_1277),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1877),
.B(n_1676),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1765),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1785),
.B(n_1683),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1862),
.A2(n_1693),
.B1(n_1326),
.B2(n_1314),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1817),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1891),
.B(n_1011),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1877),
.B(n_1693),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1789),
.B(n_1277),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1842),
.B(n_1011),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1880),
.B(n_1326),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1826),
.B(n_1286),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1818),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1844),
.B(n_1011),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1880),
.B(n_1326),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1847),
.B(n_1027),
.Y(n_1976)
);

INVxp67_ASAP7_75t_L g1977 ( 
.A(n_1882),
.Y(n_1977)
);

OAI22xp33_ASAP7_75t_L g1978 ( 
.A1(n_1879),
.A2(n_1303),
.B1(n_1304),
.B2(n_1286),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1786),
.B(n_1027),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1819),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1797),
.B(n_1326),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1807),
.B(n_820),
.Y(n_1982)
);

OAI22xp33_ASAP7_75t_R g1983 ( 
.A1(n_1874),
.A2(n_966),
.B1(n_1013),
.B2(n_895),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1807),
.B(n_823),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1771),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1805),
.B(n_846),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1828),
.B(n_1829),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1772),
.B(n_1792),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1857),
.B(n_1303),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1859),
.A2(n_1334),
.B1(n_1335),
.B2(n_1304),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1801),
.B(n_900),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_L g1992 ( 
.A(n_1812),
.B(n_1334),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1767),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1820),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1903),
.B(n_1335),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1881),
.B(n_1901),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1801),
.B(n_1806),
.Y(n_1997)
);

INVx2_ASAP7_75t_L g1998 ( 
.A(n_1821),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1838),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1793),
.Y(n_2000)
);

BUFx6f_ASAP7_75t_L g2001 ( 
.A(n_1771),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1796),
.A2(n_1649),
.B1(n_1341),
.B2(n_1344),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1799),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1914),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1806),
.B(n_1340),
.Y(n_2005)
);

INVxp67_ASAP7_75t_L g2006 ( 
.A(n_1800),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1914),
.Y(n_2007)
);

INVx2_ASAP7_75t_SL g2008 ( 
.A(n_1813),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1836),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1830),
.B(n_1762),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1767),
.Y(n_2011)
);

NAND3xp33_ASAP7_75t_L g2012 ( 
.A(n_1837),
.B(n_1875),
.C(n_1888),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1830),
.B(n_901),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1836),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1831),
.B(n_909),
.Y(n_2015)
);

AO221x1_ASAP7_75t_L g2016 ( 
.A1(n_1758),
.A2(n_835),
.B1(n_837),
.B2(n_833),
.C(n_830),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1883),
.Y(n_2017)
);

NOR2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1835),
.B(n_1340),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1831),
.A2(n_1344),
.B1(n_1341),
.B2(n_845),
.Y(n_2019)
);

OAI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_1883),
.A2(n_1103),
.B1(n_1138),
.B2(n_1082),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1831),
.B(n_910),
.Y(n_2021)
);

OR2x2_ASAP7_75t_L g2022 ( 
.A(n_1769),
.B(n_1149),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1851),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1831),
.B(n_911),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1896),
.B(n_915),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1886),
.B(n_917),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1851),
.Y(n_2027)
);

OR2x2_ASAP7_75t_L g2028 ( 
.A(n_1856),
.B(n_1220),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1890),
.B(n_1795),
.Y(n_2029)
);

OR2x2_ASAP7_75t_L g2030 ( 
.A(n_1757),
.B(n_1225),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1886),
.B(n_1027),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1843),
.Y(n_2032)
);

INVx8_ASAP7_75t_L g2033 ( 
.A(n_1790),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1896),
.B(n_920),
.Y(n_2034)
);

NOR2xp33_ASAP7_75t_L g2035 ( 
.A(n_1804),
.B(n_1246),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1898),
.B(n_928),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1846),
.Y(n_2037)
);

INVxp67_ASAP7_75t_L g2038 ( 
.A(n_1758),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1841),
.Y(n_2039)
);

AO22x2_ASAP7_75t_L g2040 ( 
.A1(n_1875),
.A2(n_1338),
.B1(n_1346),
.B2(n_1264),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1910),
.B(n_931),
.Y(n_2041)
);

INVx2_ASAP7_75t_SL g2042 ( 
.A(n_1790),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1848),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1858),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1869),
.B(n_848),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1873),
.Y(n_2046)
);

BUFx3_ASAP7_75t_L g2047 ( 
.A(n_1790),
.Y(n_2047)
);

AND2x2_ASAP7_75t_SL g2048 ( 
.A(n_1912),
.B(n_868),
.Y(n_2048)
);

O2A1O1Ixp5_ASAP7_75t_L g2049 ( 
.A1(n_1853),
.A2(n_1866),
.B(n_1867),
.C(n_1863),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1898),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1895),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1811),
.B(n_933),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1915),
.B(n_934),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1899),
.A2(n_906),
.B1(n_921),
.B2(n_898),
.Y(n_2054)
);

AOI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_1900),
.A2(n_937),
.B1(n_938),
.B2(n_936),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1783),
.A2(n_849),
.B(n_841),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1860),
.B(n_943),
.Y(n_2057)
);

OR2x6_ASAP7_75t_L g2058 ( 
.A(n_1908),
.B(n_898),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1870),
.B(n_944),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1876),
.B(n_946),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1910),
.B(n_947),
.Y(n_2061)
);

NAND3xp33_ASAP7_75t_L g2062 ( 
.A(n_1871),
.B(n_949),
.C(n_948),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1845),
.B(n_950),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1902),
.Y(n_2064)
);

INVx3_ASAP7_75t_L g2065 ( 
.A(n_1845),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1905),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1864),
.B(n_1906),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1889),
.B(n_1065),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1907),
.A2(n_921),
.B1(n_962),
.B2(n_906),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1815),
.A2(n_855),
.B(n_851),
.Y(n_2070)
);

OAI221xp5_ASAP7_75t_L g2071 ( 
.A1(n_1878),
.A2(n_870),
.B1(n_875),
.B2(n_866),
.C(n_863),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1911),
.B(n_953),
.Y(n_2072)
);

BUFx12f_ASAP7_75t_L g2073 ( 
.A(n_1824),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1840),
.B(n_1766),
.Y(n_2074)
);

OAI22xp5_ASAP7_75t_L g2075 ( 
.A1(n_1815),
.A2(n_955),
.B1(n_956),
.B2(n_954),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1822),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1845),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1822),
.Y(n_2078)
);

AND2x4_ASAP7_75t_L g2079 ( 
.A(n_1840),
.B(n_878),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1911),
.B(n_961),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1761),
.B(n_964),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1854),
.B(n_967),
.Y(n_2082)
);

INVx8_ASAP7_75t_L g2083 ( 
.A(n_1840),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1761),
.B(n_970),
.Y(n_2084)
);

OR2x6_ASAP7_75t_L g2085 ( 
.A(n_1897),
.B(n_962),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_1904),
.B(n_850),
.Y(n_2086)
);

INVx8_ASAP7_75t_L g2087 ( 
.A(n_1854),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1916),
.A2(n_1913),
.B1(n_1854),
.B2(n_1893),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_1922),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1937),
.B(n_1892),
.Y(n_2090)
);

BUFx2_ASAP7_75t_L g2091 ( 
.A(n_1928),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1922),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2039),
.B(n_1764),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2004),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2007),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_2011),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1963),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2044),
.B(n_1764),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1919),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1939),
.A2(n_1850),
.B(n_1833),
.Y(n_2100)
);

OAI21xp33_ASAP7_75t_L g2101 ( 
.A1(n_1989),
.A2(n_852),
.B(n_850),
.Y(n_2101)
);

INVx2_ASAP7_75t_SL g2102 ( 
.A(n_1950),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_1954),
.B(n_1798),
.Y(n_2103)
);

NOR2xp33_ASAP7_75t_L g2104 ( 
.A(n_1959),
.B(n_1961),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1929),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2008),
.B(n_1927),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2046),
.B(n_1798),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_1982),
.Y(n_2108)
);

INVxp67_ASAP7_75t_L g2109 ( 
.A(n_1958),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_2033),
.Y(n_2110)
);

AOI22xp33_ASAP7_75t_L g2111 ( 
.A1(n_1988),
.A2(n_1855),
.B1(n_1885),
.B2(n_1833),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1963),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1945),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2010),
.B(n_1855),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_1972),
.B(n_1885),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_1996),
.B(n_1893),
.Y(n_2116)
);

AND2x4_ASAP7_75t_L g2117 ( 
.A(n_2074),
.B(n_1892),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1987),
.B(n_1872),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2003),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1993),
.Y(n_2120)
);

OR2x6_ASAP7_75t_L g2121 ( 
.A(n_2033),
.B(n_1834),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1993),
.Y(n_2122)
);

AOI22xp5_ASAP7_75t_L g2123 ( 
.A1(n_2012),
.A2(n_974),
.B1(n_975),
.B2(n_973),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_SL g2124 ( 
.A1(n_1924),
.A2(n_1171),
.B1(n_877),
.B2(n_889),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1930),
.B(n_977),
.Y(n_2125)
);

AOI21xp5_ASAP7_75t_L g2126 ( 
.A1(n_1941),
.A2(n_894),
.B(n_893),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1925),
.Y(n_2127)
);

BUFx3_ASAP7_75t_L g2128 ( 
.A(n_2083),
.Y(n_2128)
);

NOR3xp33_ASAP7_75t_SL g2129 ( 
.A(n_1978),
.B(n_856),
.C(n_852),
.Y(n_2129)
);

BUFx4f_ASAP7_75t_L g2130 ( 
.A(n_2083),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1933),
.B(n_981),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1926),
.Y(n_2132)
);

AND2x6_ASAP7_75t_SL g2133 ( 
.A(n_1944),
.B(n_902),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_2005),
.B(n_1977),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_SL g2135 ( 
.A(n_1926),
.B(n_1985),
.Y(n_2135)
);

HB1xp67_ASAP7_75t_L g2136 ( 
.A(n_1982),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_2047),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_1953),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_SL g2139 ( 
.A(n_1926),
.B(n_982),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_SL g2140 ( 
.A(n_1985),
.B(n_984),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1949),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_1934),
.B(n_985),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1966),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1985),
.B(n_988),
.Y(n_2144)
);

INVxp67_ASAP7_75t_SL g2145 ( 
.A(n_2001),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_1951),
.Y(n_2146)
);

NAND3xp33_ASAP7_75t_L g2147 ( 
.A(n_2019),
.B(n_990),
.C(n_989),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1973),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1932),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_1992),
.B(n_991),
.Y(n_2150)
);

INVxp67_ASAP7_75t_L g2151 ( 
.A(n_2028),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1935),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_SL g2153 ( 
.A(n_2002),
.B(n_857),
.C(n_856),
.Y(n_2153)
);

CKINVDCx5p33_ASAP7_75t_R g2154 ( 
.A(n_1931),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1957),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1921),
.B(n_994),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_2001),
.B(n_997),
.Y(n_2157)
);

AOI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_1923),
.A2(n_1002),
.B1(n_1003),
.B2(n_999),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1980),
.Y(n_2159)
);

O2A1O1Ixp33_ASAP7_75t_L g2160 ( 
.A1(n_2038),
.A2(n_907),
.B(n_908),
.C(n_905),
.Y(n_2160)
);

INVx2_ASAP7_75t_SL g2161 ( 
.A(n_1984),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_SL g2162 ( 
.A(n_2001),
.B(n_1005),
.Y(n_2162)
);

BUFx6f_ASAP7_75t_L g2163 ( 
.A(n_2087),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_2072),
.B(n_1006),
.Y(n_2164)
);

INVx1_ASAP7_75t_SL g2165 ( 
.A(n_2022),
.Y(n_2165)
);

OAI22xp5_ASAP7_75t_SL g2166 ( 
.A1(n_2058),
.A2(n_881),
.B1(n_891),
.B2(n_861),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_1967),
.B(n_1065),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_1962),
.Y(n_2168)
);

INVx3_ASAP7_75t_SL g2169 ( 
.A(n_1960),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_1984),
.Y(n_2170)
);

BUFx6f_ASAP7_75t_L g2171 ( 
.A(n_2087),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_2080),
.B(n_1010),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1968),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2017),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_2074),
.B(n_912),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2017),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1999),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_2079),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1936),
.B(n_1014),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1979),
.B(n_1065),
.Y(n_2180)
);

NOR2x1p5_ASAP7_75t_L g2181 ( 
.A(n_2073),
.B(n_857),
.Y(n_2181)
);

INVx4_ASAP7_75t_L g2182 ( 
.A(n_1938),
.Y(n_2182)
);

CKINVDCx20_ASAP7_75t_R g2183 ( 
.A(n_1995),
.Y(n_2183)
);

NAND3xp33_ASAP7_75t_SL g2184 ( 
.A(n_2018),
.B(n_861),
.C(n_858),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2051),
.Y(n_2185)
);

NOR2xp33_ASAP7_75t_R g2186 ( 
.A(n_2042),
.B(n_858),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1994),
.Y(n_2187)
);

O2A1O1Ixp33_ASAP7_75t_L g2188 ( 
.A1(n_1947),
.A2(n_916),
.B(n_919),
.C(n_914),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_2065),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2000),
.Y(n_2190)
);

CKINVDCx20_ASAP7_75t_R g2191 ( 
.A(n_2006),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_2030),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1998),
.B(n_1016),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_2064),
.Y(n_2194)
);

AOI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_2048),
.A2(n_1015),
.B1(n_1040),
.B2(n_969),
.Y(n_2195)
);

INVxp67_ASAP7_75t_L g2196 ( 
.A(n_2052),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_2029),
.Y(n_2197)
);

HB1xp67_ASAP7_75t_L g2198 ( 
.A(n_2077),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1943),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_1964),
.B(n_923),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_2065),
.Y(n_2201)
);

BUFx6f_ASAP7_75t_L g2202 ( 
.A(n_2014),
.Y(n_2202)
);

CKINVDCx5p33_ASAP7_75t_R g2203 ( 
.A(n_2058),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2064),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2032),
.B(n_924),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1946),
.B(n_1019),
.Y(n_2206)
);

INVx5_ASAP7_75t_L g2207 ( 
.A(n_2085),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2081),
.B(n_1020),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2037),
.B(n_926),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1965),
.B(n_1022),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1981),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2023),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2076),
.Y(n_2213)
);

INVx2_ASAP7_75t_L g2214 ( 
.A(n_2027),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2076),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2078),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2078),
.Y(n_2217)
);

AOI22xp33_ASAP7_75t_L g2218 ( 
.A1(n_2016),
.A2(n_1015),
.B1(n_1040),
.B2(n_969),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_2043),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_SL g2220 ( 
.A(n_1990),
.B(n_871),
.C(n_869),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_2079),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2067),
.B(n_1023),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_2066),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_1970),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1991),
.B(n_2013),
.Y(n_2225)
);

AND2x6_ASAP7_75t_L g2226 ( 
.A(n_1948),
.B(n_1072),
.Y(n_2226)
);

AOI22xp33_ASAP7_75t_L g2227 ( 
.A1(n_1969),
.A2(n_1104),
.B1(n_1108),
.B2(n_1072),
.Y(n_2227)
);

INVx2_ASAP7_75t_SL g2228 ( 
.A(n_2031),
.Y(n_2228)
);

NOR2xp33_ASAP7_75t_L g2229 ( 
.A(n_2045),
.B(n_1024),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1974),
.B(n_1083),
.Y(n_2230)
);

NOR2x1p5_ASAP7_75t_L g2231 ( 
.A(n_1986),
.B(n_869),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2084),
.B(n_1026),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2050),
.Y(n_2233)
);

INVx5_ASAP7_75t_L g2234 ( 
.A(n_2085),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1997),
.B(n_1030),
.Y(n_2235)
);

INVxp67_ASAP7_75t_L g2236 ( 
.A(n_1976),
.Y(n_2236)
);

INVx4_ASAP7_75t_L g2237 ( 
.A(n_2068),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_2009),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1955),
.B(n_1032),
.Y(n_2239)
);

NAND2xp33_ASAP7_75t_SL g2240 ( 
.A(n_2163),
.B(n_1952),
.Y(n_2240)
);

NAND2xp33_ASAP7_75t_SL g2241 ( 
.A(n_2163),
.B(n_2041),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2196),
.B(n_2035),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2150),
.B(n_2025),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_2106),
.B(n_1942),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_SL g2245 ( 
.A(n_2104),
.B(n_2055),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_2103),
.B(n_2020),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_2106),
.B(n_1940),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_2197),
.B(n_2034),
.Y(n_2248)
);

NAND2xp33_ASAP7_75t_SL g2249 ( 
.A(n_2163),
.B(n_2061),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_SL g2250 ( 
.A(n_2224),
.B(n_2036),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2117),
.B(n_2063),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2168),
.B(n_2075),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2192),
.B(n_2062),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2207),
.B(n_2086),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2173),
.B(n_2114),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_SL g2256 ( 
.A(n_2207),
.B(n_2053),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2207),
.B(n_2057),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2234),
.B(n_2059),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2234),
.B(n_2151),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_2234),
.B(n_2060),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_2091),
.B(n_1920),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_2102),
.B(n_2026),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_SL g2263 ( 
.A(n_2109),
.B(n_2082),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_SL g2264 ( 
.A(n_2228),
.B(n_2015),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_2237),
.B(n_2021),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_2236),
.B(n_2116),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2115),
.B(n_2024),
.Y(n_2267)
);

NAND2xp33_ASAP7_75t_SL g2268 ( 
.A(n_2171),
.B(n_1956),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2165),
.B(n_1918),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_SL g2270 ( 
.A(n_2134),
.B(n_2070),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_SL g2271 ( 
.A(n_2232),
.B(n_1917),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_2222),
.B(n_2054),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2183),
.B(n_2069),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2180),
.B(n_2056),
.Y(n_2274)
);

NAND2xp33_ASAP7_75t_SL g2275 ( 
.A(n_2171),
.B(n_1971),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_SL g2276 ( 
.A(n_2093),
.B(n_1975),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2098),
.B(n_2049),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2125),
.B(n_2040),
.Y(n_2278)
);

NAND2xp33_ASAP7_75t_SL g2279 ( 
.A(n_2171),
.B(n_1983),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_SL g2280 ( 
.A(n_2107),
.B(n_871),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2225),
.B(n_873),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_SL g2282 ( 
.A(n_2203),
.B(n_873),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_SL g2283 ( 
.A(n_2161),
.B(n_874),
.Y(n_2283)
);

XNOR2x2_ASAP7_75t_L g2284 ( 
.A(n_2147),
.B(n_2040),
.Y(n_2284)
);

NAND2xp33_ASAP7_75t_SL g2285 ( 
.A(n_2220),
.B(n_874),
.Y(n_2285)
);

NAND2xp33_ASAP7_75t_SL g2286 ( 
.A(n_2129),
.B(n_876),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_SL g2287 ( 
.A(n_2178),
.B(n_876),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2221),
.B(n_877),
.Y(n_2288)
);

NAND2xp33_ASAP7_75t_SL g2289 ( 
.A(n_2231),
.B(n_2182),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_2229),
.B(n_880),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_SL g2291 ( 
.A(n_2108),
.B(n_880),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_SL g2292 ( 
.A(n_2136),
.B(n_881),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_SL g2293 ( 
.A(n_2170),
.B(n_882),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_SL g2294 ( 
.A(n_2167),
.B(n_882),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_SL g2295 ( 
.A(n_2230),
.B(n_883),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_SL g2296 ( 
.A(n_2127),
.B(n_883),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_2149),
.B(n_884),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2131),
.B(n_2071),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_SL g2299 ( 
.A(n_2152),
.B(n_884),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_SL g2300 ( 
.A(n_2155),
.B(n_885),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_2156),
.B(n_885),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2142),
.B(n_930),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_SL g2303 ( 
.A(n_2118),
.B(n_2094),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_SL g2304 ( 
.A(n_2095),
.B(n_2130),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_2117),
.B(n_888),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_SL g2306 ( 
.A(n_2238),
.B(n_888),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_SL g2307 ( 
.A(n_2238),
.B(n_889),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2238),
.B(n_890),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_SL g2309 ( 
.A(n_2090),
.B(n_890),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_SL g2310 ( 
.A(n_2185),
.B(n_891),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2141),
.B(n_892),
.Y(n_2311)
);

NAND2xp33_ASAP7_75t_SL g2312 ( 
.A(n_2154),
.B(n_892),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2153),
.B(n_1034),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2143),
.B(n_1106),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_SL g2315 ( 
.A(n_2148),
.B(n_1106),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_SL g2316 ( 
.A(n_2159),
.B(n_1141),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_SL g2317 ( 
.A(n_2110),
.B(n_1141),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2199),
.B(n_942),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2179),
.B(n_945),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_SL g2320 ( 
.A(n_2187),
.B(n_1329),
.Y(n_2320)
);

NAND2xp5_ASAP7_75t_L g2321 ( 
.A(n_2206),
.B(n_951),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2202),
.B(n_1329),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2200),
.B(n_1083),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_SL g2324 ( 
.A(n_2202),
.B(n_1330),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_SL g2325 ( 
.A(n_2202),
.B(n_2177),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_2200),
.B(n_1083),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2235),
.B(n_2190),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_SL g2328 ( 
.A(n_2132),
.B(n_1330),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_2175),
.B(n_1331),
.Y(n_2329)
);

NAND2xp33_ASAP7_75t_SL g2330 ( 
.A(n_2132),
.B(n_1331),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_2175),
.B(n_1332),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2101),
.B(n_1204),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_SL g2333 ( 
.A(n_2099),
.B(n_1332),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2105),
.B(n_1333),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2205),
.B(n_957),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2113),
.B(n_2119),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2111),
.B(n_1333),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2205),
.B(n_958),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_2239),
.B(n_1036),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2128),
.B(n_963),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2194),
.B(n_1336),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2204),
.B(n_1336),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2209),
.B(n_978),
.Y(n_2343)
);

NAND2xp33_ASAP7_75t_SL g2344 ( 
.A(n_2132),
.B(n_1337),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_SL g2345 ( 
.A(n_2219),
.B(n_1337),
.Y(n_2345)
);

NAND2xp33_ASAP7_75t_SL g2346 ( 
.A(n_2191),
.B(n_1339),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2209),
.B(n_979),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2223),
.B(n_2088),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2186),
.B(n_1339),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_SL g2350 ( 
.A(n_2212),
.B(n_1342),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_SL g2351 ( 
.A(n_2214),
.B(n_1342),
.Y(n_2351)
);

NAND2xp33_ASAP7_75t_SL g2352 ( 
.A(n_2169),
.B(n_1349),
.Y(n_2352)
);

NAND2xp33_ASAP7_75t_SL g2353 ( 
.A(n_2189),
.B(n_1350),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_SL g2354 ( 
.A(n_2158),
.B(n_1350),
.Y(n_2354)
);

NAND2xp33_ASAP7_75t_SL g2355 ( 
.A(n_2189),
.B(n_1351),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2123),
.B(n_1351),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_SL g2357 ( 
.A(n_2189),
.B(n_1352),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2201),
.B(n_1352),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2201),
.B(n_1353),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_SL g2360 ( 
.A(n_2201),
.B(n_1356),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_SL g2361 ( 
.A(n_2233),
.B(n_1356),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_SL g2362 ( 
.A(n_2193),
.B(n_1204),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_SL g2363 ( 
.A(n_2198),
.B(n_2124),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2210),
.B(n_2166),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_SL g2365 ( 
.A(n_2164),
.B(n_1204),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2227),
.B(n_1206),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2195),
.B(n_1206),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_SL g2368 ( 
.A(n_2172),
.B(n_2208),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2096),
.B(n_1206),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2160),
.B(n_1213),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_SL g2371 ( 
.A(n_2137),
.B(n_1213),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2139),
.B(n_2157),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2140),
.B(n_1213),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2144),
.B(n_1217),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_2162),
.B(n_1217),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2211),
.B(n_980),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_SL g2377 ( 
.A(n_2138),
.B(n_1217),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_SL g2378 ( 
.A(n_2089),
.B(n_1229),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_SL g2379 ( 
.A(n_2092),
.B(n_1229),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_SL g2380 ( 
.A(n_2097),
.B(n_1229),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2218),
.B(n_1037),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_2112),
.B(n_1038),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_SL g2383 ( 
.A(n_2120),
.B(n_1039),
.Y(n_2383)
);

NAND2xp33_ASAP7_75t_SL g2384 ( 
.A(n_2122),
.B(n_1104),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_SL g2385 ( 
.A(n_2146),
.B(n_1045),
.Y(n_2385)
);

NAND2xp33_ASAP7_75t_SL g2386 ( 
.A(n_2135),
.B(n_1108),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2126),
.B(n_2226),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2188),
.B(n_1047),
.Y(n_2388)
);

NAND2xp33_ASAP7_75t_SL g2389 ( 
.A(n_2174),
.B(n_1199),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2226),
.B(n_983),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_SL g2391 ( 
.A(n_2176),
.B(n_1049),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_2213),
.B(n_2215),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2243),
.B(n_2184),
.Y(n_2393)
);

BUFx2_ASAP7_75t_L g2394 ( 
.A(n_2244),
.Y(n_2394)
);

INVxp67_ASAP7_75t_L g2395 ( 
.A(n_2242),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2245),
.A2(n_2226),
.B1(n_1054),
.B2(n_1055),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2244),
.B(n_2145),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2392),
.Y(n_2398)
);

A2O1A1Ixp33_ASAP7_75t_L g2399 ( 
.A1(n_2339),
.A2(n_2100),
.B(n_2217),
.C(n_2216),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2255),
.B(n_2226),
.Y(n_2400)
);

INVx5_ASAP7_75t_L g2401 ( 
.A(n_2251),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_2251),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2327),
.B(n_2133),
.Y(n_2403)
);

NOR2x1_ASAP7_75t_L g2404 ( 
.A(n_2271),
.B(n_2121),
.Y(n_2404)
);

AOI22x1_ASAP7_75t_L g2405 ( 
.A1(n_2332),
.A2(n_2367),
.B1(n_2381),
.B2(n_2366),
.Y(n_2405)
);

HB1xp67_ASAP7_75t_L g2406 ( 
.A(n_2247),
.Y(n_2406)
);

BUFx2_ASAP7_75t_L g2407 ( 
.A(n_2247),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2339),
.B(n_2252),
.Y(n_2408)
);

OAI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2278),
.A2(n_1211),
.B1(n_1236),
.B2(n_1199),
.Y(n_2409)
);

AOI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2313),
.A2(n_2364),
.B1(n_2290),
.B2(n_2284),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2336),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2376),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2325),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2318),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2323),
.B(n_2181),
.Y(n_2415)
);

BUFx6f_ASAP7_75t_L g2416 ( 
.A(n_2304),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2326),
.B(n_2273),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2279),
.Y(n_2418)
);

CKINVDCx5p33_ASAP7_75t_R g2419 ( 
.A(n_2346),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2348),
.Y(n_2420)
);

AND3x1_ASAP7_75t_SL g2421 ( 
.A(n_2363),
.B(n_995),
.C(n_987),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_2340),
.Y(n_2422)
);

INVx4_ASAP7_75t_L g2423 ( 
.A(n_2340),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2335),
.B(n_2338),
.Y(n_2424)
);

BUFx4f_ASAP7_75t_L g2425 ( 
.A(n_2289),
.Y(n_2425)
);

BUFx3_ASAP7_75t_L g2426 ( 
.A(n_2343),
.Y(n_2426)
);

CKINVDCx20_ASAP7_75t_R g2427 ( 
.A(n_2312),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2352),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2390),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2298),
.B(n_1051),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2353),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2266),
.Y(n_2432)
);

AND2x2_ASAP7_75t_L g2433 ( 
.A(n_2347),
.B(n_2121),
.Y(n_2433)
);

NAND3xp33_ASAP7_75t_SL g2434 ( 
.A(n_2370),
.B(n_1061),
.C(n_1057),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2303),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2302),
.B(n_2321),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2264),
.Y(n_2437)
);

OR2x2_ASAP7_75t_L g2438 ( 
.A(n_2319),
.B(n_996),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_SL g2439 ( 
.A(n_2254),
.B(n_1324),
.Y(n_2439)
);

BUFx2_ASAP7_75t_L g2440 ( 
.A(n_2355),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2246),
.B(n_1056),
.Y(n_2441)
);

AND3x1_ASAP7_75t_SL g2442 ( 
.A(n_2285),
.B(n_1001),
.C(n_1000),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2356),
.B(n_1007),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2270),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2276),
.B(n_1008),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2248),
.B(n_1062),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2309),
.B(n_1064),
.Y(n_2447)
);

CKINVDCx5p33_ASAP7_75t_R g2448 ( 
.A(n_2385),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2267),
.Y(n_2449)
);

AND3x1_ASAP7_75t_SL g2450 ( 
.A(n_2286),
.B(n_1012),
.C(n_1009),
.Y(n_2450)
);

NAND2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2259),
.B(n_1017),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2384),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2256),
.B(n_1321),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2281),
.B(n_1068),
.Y(n_2454)
);

BUFx12f_ASAP7_75t_L g2455 ( 
.A(n_2328),
.Y(n_2455)
);

INVxp67_ASAP7_75t_L g2456 ( 
.A(n_2253),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2257),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_2301),
.B(n_1075),
.Y(n_2458)
);

AND2x2_ASAP7_75t_L g2459 ( 
.A(n_2295),
.B(n_1018),
.Y(n_2459)
);

OR2x2_ASAP7_75t_L g2460 ( 
.A(n_2261),
.B(n_1028),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2294),
.B(n_1029),
.Y(n_2461)
);

BUFx6f_ASAP7_75t_L g2462 ( 
.A(n_2258),
.Y(n_2462)
);

CKINVDCx20_ASAP7_75t_R g2463 ( 
.A(n_2241),
.Y(n_2463)
);

AND2x2_ASAP7_75t_SL g2464 ( 
.A(n_2387),
.B(n_1211),
.Y(n_2464)
);

CKINVDCx5p33_ASAP7_75t_R g2465 ( 
.A(n_2282),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_2260),
.Y(n_2466)
);

HB1xp67_ASAP7_75t_L g2467 ( 
.A(n_2306),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2362),
.B(n_1076),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2277),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2354),
.A2(n_1035),
.B1(n_1044),
.B2(n_1031),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2389),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2280),
.B(n_1078),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_2250),
.B(n_1080),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_2269),
.B(n_1084),
.Y(n_2474)
);

NAND2x1p5_ASAP7_75t_L g2475 ( 
.A(n_2265),
.B(n_1046),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2296),
.B(n_1048),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_L g2477 ( 
.A(n_2329),
.B(n_1085),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2382),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2383),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2297),
.B(n_2299),
.Y(n_2480)
);

BUFx2_ASAP7_75t_L g2481 ( 
.A(n_2249),
.Y(n_2481)
);

CKINVDCx5p33_ASAP7_75t_R g2482 ( 
.A(n_2262),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2274),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_SL g2484 ( 
.A(n_2307),
.B(n_1322),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2331),
.B(n_2368),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2391),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2308),
.B(n_1086),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2300),
.B(n_1087),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2310),
.B(n_1088),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2341),
.B(n_1050),
.Y(n_2490)
);

AND2x2_ASAP7_75t_L g2491 ( 
.A(n_2342),
.B(n_1052),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2263),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2372),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2378),
.B(n_1090),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2322),
.B(n_1058),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2379),
.B(n_1093),
.Y(n_2496)
);

OR2x2_ASAP7_75t_L g2497 ( 
.A(n_2324),
.B(n_1060),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2380),
.B(n_1096),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2386),
.Y(n_2499)
);

INVx3_ASAP7_75t_L g2500 ( 
.A(n_2275),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_L g2501 ( 
.A(n_2305),
.B(n_2291),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2311),
.B(n_1066),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2314),
.B(n_1067),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2315),
.B(n_1071),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2292),
.B(n_1098),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2377),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2350),
.Y(n_2507)
);

AOI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2369),
.A2(n_1100),
.B1(n_1101),
.B2(n_1099),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2351),
.Y(n_2509)
);

A2O1A1Ixp33_ASAP7_75t_L g2510 ( 
.A1(n_2272),
.A2(n_1271),
.B(n_1282),
.C(n_1236),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2316),
.B(n_1074),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2361),
.Y(n_2512)
);

BUFx3_ASAP7_75t_L g2513 ( 
.A(n_2240),
.Y(n_2513)
);

OAI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_2373),
.A2(n_1282),
.B1(n_1316),
.B2(n_1271),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2320),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2333),
.Y(n_2516)
);

INVx3_ASAP7_75t_L g2517 ( 
.A(n_2268),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2365),
.B(n_1325),
.Y(n_2518)
);

NAND2xp33_ASAP7_75t_SL g2519 ( 
.A(n_2371),
.B(n_1109),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2293),
.B(n_1111),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2388),
.B(n_1077),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2334),
.Y(n_2522)
);

CKINVDCx8_ASAP7_75t_R g2523 ( 
.A(n_2330),
.Y(n_2523)
);

INVx4_ASAP7_75t_L g2524 ( 
.A(n_2344),
.Y(n_2524)
);

CKINVDCx11_ASAP7_75t_R g2525 ( 
.A(n_2317),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2345),
.B(n_1079),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2357),
.B(n_1081),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2358),
.Y(n_2528)
);

AND2x2_ASAP7_75t_L g2529 ( 
.A(n_2359),
.B(n_1089),
.Y(n_2529)
);

AND2x2_ASAP7_75t_L g2530 ( 
.A(n_2360),
.B(n_1091),
.Y(n_2530)
);

INVx3_ASAP7_75t_L g2531 ( 
.A(n_2287),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2288),
.B(n_1094),
.Y(n_2532)
);

AOI22xp33_ASAP7_75t_L g2533 ( 
.A1(n_2337),
.A2(n_2375),
.B1(n_2374),
.B2(n_2349),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2283),
.Y(n_2534)
);

BUFx6f_ASAP7_75t_L g2535 ( 
.A(n_2416),
.Y(n_2535)
);

AO21x2_ASAP7_75t_L g2536 ( 
.A1(n_2469),
.A2(n_1097),
.B(n_1095),
.Y(n_2536)
);

INVx1_ASAP7_75t_SL g2537 ( 
.A(n_2482),
.Y(n_2537)
);

OAI21x1_ASAP7_75t_L g2538 ( 
.A1(n_2483),
.A2(n_2444),
.B(n_2400),
.Y(n_2538)
);

NAND2x1p5_ASAP7_75t_L g2539 ( 
.A(n_2517),
.B(n_2513),
.Y(n_2539)
);

OAI21x1_ASAP7_75t_L g2540 ( 
.A1(n_2400),
.A2(n_2500),
.B(n_2420),
.Y(n_2540)
);

BUFx2_ASAP7_75t_R g2541 ( 
.A(n_2418),
.Y(n_2541)
);

OA21x2_ASAP7_75t_L g2542 ( 
.A1(n_2399),
.A2(n_1105),
.B(n_1102),
.Y(n_2542)
);

CKINVDCx20_ASAP7_75t_R g2543 ( 
.A(n_2427),
.Y(n_2543)
);

OAI21x1_ASAP7_75t_L g2544 ( 
.A1(n_2500),
.A2(n_1348),
.B(n_1319),
.Y(n_2544)
);

OAI21x1_ASAP7_75t_L g2545 ( 
.A1(n_2405),
.A2(n_1348),
.B(n_1319),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2398),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2407),
.B(n_1107),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2435),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_2411),
.Y(n_2549)
);

BUFx4f_ASAP7_75t_L g2550 ( 
.A(n_2416),
.Y(n_2550)
);

INVx5_ASAP7_75t_L g2551 ( 
.A(n_2517),
.Y(n_2551)
);

OAI21xp5_ASAP7_75t_L g2552 ( 
.A1(n_2393),
.A2(n_1209),
.B(n_1133),
.Y(n_2552)
);

INVxp67_ASAP7_75t_SL g2553 ( 
.A(n_2432),
.Y(n_2553)
);

OAI21x1_ASAP7_75t_L g2554 ( 
.A1(n_2449),
.A2(n_1355),
.B(n_1316),
.Y(n_2554)
);

OAI21xp5_ASAP7_75t_L g2555 ( 
.A1(n_2408),
.A2(n_1251),
.B(n_1226),
.Y(n_2555)
);

INVx2_ASAP7_75t_SL g2556 ( 
.A(n_2416),
.Y(n_2556)
);

AOI22x1_ASAP7_75t_L g2557 ( 
.A1(n_2452),
.A2(n_2471),
.B1(n_2412),
.B2(n_2414),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2406),
.B(n_1354),
.Y(n_2558)
);

OAI21x1_ASAP7_75t_L g2559 ( 
.A1(n_2404),
.A2(n_1355),
.B(n_1124),
.Y(n_2559)
);

AND2x4_ASAP7_75t_L g2560 ( 
.A(n_2401),
.B(n_797),
.Y(n_2560)
);

OR2x6_ASAP7_75t_L g2561 ( 
.A(n_2423),
.B(n_1308),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2413),
.Y(n_2562)
);

OAI21x1_ASAP7_75t_L g2563 ( 
.A1(n_2404),
.A2(n_1130),
.B(n_1118),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2429),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_L g2565 ( 
.A(n_2425),
.Y(n_2565)
);

BUFx3_ASAP7_75t_L g2566 ( 
.A(n_2433),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_2425),
.Y(n_2567)
);

INVx1_ASAP7_75t_SL g2568 ( 
.A(n_2394),
.Y(n_2568)
);

INVx4_ASAP7_75t_L g2569 ( 
.A(n_2423),
.Y(n_2569)
);

OAI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2436),
.A2(n_1294),
.B(n_1152),
.Y(n_2570)
);

AO21x2_ASAP7_75t_L g2571 ( 
.A1(n_2510),
.A2(n_1137),
.B(n_1131),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2437),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2492),
.Y(n_2573)
);

INVx5_ASAP7_75t_L g2574 ( 
.A(n_2524),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2445),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2493),
.Y(n_2576)
);

AOI22x1_ASAP7_75t_L g2577 ( 
.A1(n_2475),
.A2(n_2481),
.B1(n_2499),
.B2(n_2456),
.Y(n_2577)
);

INVx3_ASAP7_75t_L g2578 ( 
.A(n_2402),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2397),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2424),
.Y(n_2580)
);

BUFx6f_ASAP7_75t_L g2581 ( 
.A(n_2457),
.Y(n_2581)
);

CKINVDCx20_ASAP7_75t_R g2582 ( 
.A(n_2463),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_2410),
.B(n_1315),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2426),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2401),
.Y(n_2585)
);

OAI21x1_ASAP7_75t_L g2586 ( 
.A1(n_2445),
.A2(n_1174),
.B(n_1144),
.Y(n_2586)
);

OAI21x1_ASAP7_75t_L g2587 ( 
.A1(n_2409),
.A2(n_1195),
.B(n_1184),
.Y(n_2587)
);

OR2x6_ASAP7_75t_L g2588 ( 
.A(n_2402),
.B(n_1345),
.Y(n_2588)
);

INVx1_ASAP7_75t_SL g2589 ( 
.A(n_2465),
.Y(n_2589)
);

INVx6_ASAP7_75t_L g2590 ( 
.A(n_2401),
.Y(n_2590)
);

INVx6_ASAP7_75t_L g2591 ( 
.A(n_2457),
.Y(n_2591)
);

CKINVDCx8_ASAP7_75t_R g2592 ( 
.A(n_2419),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2448),
.Y(n_2593)
);

AO21x2_ASAP7_75t_L g2594 ( 
.A1(n_2434),
.A2(n_1214),
.B(n_1207),
.Y(n_2594)
);

OAI21x1_ASAP7_75t_L g2595 ( 
.A1(n_2409),
.A2(n_1216),
.B(n_1215),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2521),
.Y(n_2596)
);

OAI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_2468),
.A2(n_1250),
.B(n_1247),
.Y(n_2597)
);

BUFx12f_ASAP7_75t_L g2598 ( 
.A(n_2525),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2521),
.A2(n_1267),
.B(n_1259),
.Y(n_2599)
);

INVx2_ASAP7_75t_SL g2600 ( 
.A(n_2457),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2516),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2462),
.Y(n_2602)
);

OAI21x1_ASAP7_75t_L g2603 ( 
.A1(n_2514),
.A2(n_1296),
.B(n_1292),
.Y(n_2603)
);

AO21x2_ASAP7_75t_L g2604 ( 
.A1(n_2441),
.A2(n_1298),
.B(n_1297),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2462),
.Y(n_2605)
);

OAI21x1_ASAP7_75t_SL g2606 ( 
.A1(n_2485),
.A2(n_1317),
.B(n_1312),
.Y(n_2606)
);

INVx5_ASAP7_75t_L g2607 ( 
.A(n_2524),
.Y(n_2607)
);

OAI21x1_ASAP7_75t_L g2608 ( 
.A1(n_2514),
.A2(n_1323),
.B(n_1320),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_L g2609 ( 
.A(n_2403),
.B(n_1112),
.Y(n_2609)
);

AND2x2_ASAP7_75t_L g2610 ( 
.A(n_2417),
.B(n_1327),
.Y(n_2610)
);

AOI22x1_ASAP7_75t_L g2611 ( 
.A1(n_2478),
.A2(n_1357),
.B1(n_1347),
.B2(n_1114),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2464),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2395),
.B(n_1113),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2462),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2466),
.Y(n_2615)
);

INVx8_ASAP7_75t_L g2616 ( 
.A(n_2455),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2466),
.Y(n_2617)
);

OAI21x1_ASAP7_75t_L g2618 ( 
.A1(n_2453),
.A2(n_799),
.B(n_798),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2466),
.Y(n_2619)
);

CKINVDCx11_ASAP7_75t_R g2620 ( 
.A(n_2523),
.Y(n_2620)
);

OAI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_2430),
.A2(n_1117),
.B(n_1115),
.Y(n_2621)
);

BUFx6f_ASAP7_75t_L g2622 ( 
.A(n_2422),
.Y(n_2622)
);

BUFx3_ASAP7_75t_L g2623 ( 
.A(n_2422),
.Y(n_2623)
);

OAI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2396),
.A2(n_1120),
.B(n_1119),
.Y(n_2624)
);

OAI21x1_ASAP7_75t_L g2625 ( 
.A1(n_2479),
.A2(n_2486),
.B(n_2474),
.Y(n_2625)
);

OAI21x1_ASAP7_75t_L g2626 ( 
.A1(n_2460),
.A2(n_803),
.B(n_802),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2506),
.B(n_1121),
.Y(n_2627)
);

BUFx2_ASAP7_75t_L g2628 ( 
.A(n_2467),
.Y(n_2628)
);

AOI22x1_ASAP7_75t_L g2629 ( 
.A1(n_2438),
.A2(n_1123),
.B1(n_1127),
.B2(n_1122),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2507),
.Y(n_2630)
);

BUFx8_ASAP7_75t_L g2631 ( 
.A(n_2431),
.Y(n_2631)
);

NAND2x1p5_ASAP7_75t_L g2632 ( 
.A(n_2531),
.B(n_805),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2533),
.B(n_1128),
.Y(n_2633)
);

OAI21xp5_ASAP7_75t_L g2634 ( 
.A1(n_2396),
.A2(n_1132),
.B(n_1129),
.Y(n_2634)
);

BUFx6f_ASAP7_75t_L g2635 ( 
.A(n_2440),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_L g2636 ( 
.A(n_2509),
.B(n_1288),
.Y(n_2636)
);

INVx3_ASAP7_75t_SL g2637 ( 
.A(n_2428),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2512),
.Y(n_2638)
);

INVx6_ASAP7_75t_L g2639 ( 
.A(n_2415),
.Y(n_2639)
);

AND2x2_ASAP7_75t_L g2640 ( 
.A(n_2579),
.B(n_2531),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2546),
.Y(n_2641)
);

INVx6_ASAP7_75t_L g2642 ( 
.A(n_2565),
.Y(n_2642)
);

AOI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2555),
.A2(n_2552),
.B1(n_2583),
.B2(n_2570),
.Y(n_2643)
);

AOI22xp33_ASAP7_75t_L g2644 ( 
.A1(n_2597),
.A2(n_2519),
.B1(n_2443),
.B2(n_2528),
.Y(n_2644)
);

INVx1_ASAP7_75t_SL g2645 ( 
.A(n_2584),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2580),
.B(n_2480),
.Y(n_2646)
);

CKINVDCx11_ASAP7_75t_R g2647 ( 
.A(n_2592),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2566),
.B(n_2628),
.Y(n_2648)
);

CKINVDCx11_ASAP7_75t_R g2649 ( 
.A(n_2582),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2572),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2576),
.Y(n_2651)
);

INVx4_ASAP7_75t_L g2652 ( 
.A(n_2574),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2573),
.Y(n_2653)
);

INVx4_ASAP7_75t_SL g2654 ( 
.A(n_2637),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2548),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2553),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2549),
.Y(n_2657)
);

INVx2_ASAP7_75t_L g2658 ( 
.A(n_2564),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_L g2659 ( 
.A1(n_2612),
.A2(n_2518),
.B1(n_2534),
.B2(n_2439),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_L g2660 ( 
.A(n_2596),
.B(n_2515),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2638),
.Y(n_2661)
);

INVx2_ASAP7_75t_L g2662 ( 
.A(n_2630),
.Y(n_2662)
);

AOI22xp33_ASAP7_75t_L g2663 ( 
.A1(n_2612),
.A2(n_2522),
.B1(n_2461),
.B2(n_2459),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2540),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_L g2665 ( 
.A1(n_2611),
.A2(n_2484),
.B1(n_2495),
.B2(n_2527),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2562),
.Y(n_2666)
);

INVx6_ASAP7_75t_L g2667 ( 
.A(n_2565),
.Y(n_2667)
);

INVx4_ASAP7_75t_SL g2668 ( 
.A(n_2598),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2628),
.Y(n_2669)
);

AOI22xp5_ASAP7_75t_L g2670 ( 
.A1(n_2604),
.A2(n_2421),
.B1(n_2450),
.B2(n_2442),
.Y(n_2670)
);

INVx1_ASAP7_75t_SL g2671 ( 
.A(n_2537),
.Y(n_2671)
);

CKINVDCx11_ASAP7_75t_R g2672 ( 
.A(n_2620),
.Y(n_2672)
);

INVx3_ASAP7_75t_L g2673 ( 
.A(n_2581),
.Y(n_2673)
);

CKINVDCx5p33_ASAP7_75t_R g2674 ( 
.A(n_2593),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2601),
.Y(n_2675)
);

INVx6_ASAP7_75t_L g2676 ( 
.A(n_2565),
.Y(n_2676)
);

INVx4_ASAP7_75t_L g2677 ( 
.A(n_2574),
.Y(n_2677)
);

AOI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2594),
.A2(n_2501),
.B1(n_2530),
.B2(n_2529),
.Y(n_2678)
);

INVx2_ASAP7_75t_SL g2679 ( 
.A(n_2639),
.Y(n_2679)
);

CKINVDCx20_ASAP7_75t_R g2680 ( 
.A(n_2543),
.Y(n_2680)
);

AOI22xp33_ASAP7_75t_L g2681 ( 
.A1(n_2611),
.A2(n_2532),
.B1(n_2476),
.B2(n_2491),
.Y(n_2681)
);

INVx6_ASAP7_75t_L g2682 ( 
.A(n_2567),
.Y(n_2682)
);

BUFx3_ASAP7_75t_L g2683 ( 
.A(n_2639),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_2633),
.A2(n_2490),
.B1(n_2503),
.B2(n_2502),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2538),
.Y(n_2685)
);

OAI21xp5_ASAP7_75t_SL g2686 ( 
.A1(n_2624),
.A2(n_2470),
.B(n_2508),
.Y(n_2686)
);

INVx4_ASAP7_75t_L g2687 ( 
.A(n_2574),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2596),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2575),
.Y(n_2689)
);

AOI22xp33_ASAP7_75t_SL g2690 ( 
.A1(n_2577),
.A2(n_2451),
.B1(n_2511),
.B2(n_2504),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2575),
.Y(n_2691)
);

BUFx8_ASAP7_75t_L g2692 ( 
.A(n_2567),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2567),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2634),
.A2(n_2526),
.B1(n_2496),
.B2(n_2498),
.Y(n_2694)
);

AOI22xp33_ASAP7_75t_L g2695 ( 
.A1(n_2577),
.A2(n_2494),
.B1(n_2454),
.B2(n_2446),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2605),
.Y(n_2696)
);

AO22x1_ASAP7_75t_L g2697 ( 
.A1(n_2631),
.A2(n_2473),
.B1(n_2447),
.B2(n_2458),
.Y(n_2697)
);

BUFx6f_ASAP7_75t_L g2698 ( 
.A(n_2550),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_SL g2699 ( 
.A1(n_2606),
.A2(n_2497),
.B1(n_2487),
.B2(n_2472),
.Y(n_2699)
);

CKINVDCx11_ASAP7_75t_R g2700 ( 
.A(n_2616),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2609),
.A2(n_2477),
.B1(n_2489),
.B2(n_2488),
.Y(n_2701)
);

BUFx12f_ASAP7_75t_L g2702 ( 
.A(n_2631),
.Y(n_2702)
);

AOI22xp33_ASAP7_75t_L g2703 ( 
.A1(n_2606),
.A2(n_2520),
.B1(n_2505),
.B2(n_1136),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2568),
.B(n_2508),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2635),
.A2(n_1139),
.B1(n_1143),
.B2(n_1135),
.Y(n_2705)
);

INVx1_ASAP7_75t_SL g2706 ( 
.A(n_2589),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_SL g2707 ( 
.A1(n_2557),
.A2(n_1146),
.B1(n_1147),
.B2(n_1145),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_L g2708 ( 
.A1(n_2610),
.A2(n_1150),
.B1(n_1151),
.B2(n_1148),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2625),
.B(n_1153),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2585),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2627),
.A2(n_1156),
.B1(n_1158),
.B2(n_1155),
.Y(n_2711)
);

AOI22xp33_ASAP7_75t_SL g2712 ( 
.A1(n_2557),
.A2(n_1161),
.B1(n_1162),
.B2(n_1159),
.Y(n_2712)
);

INVx4_ASAP7_75t_L g2713 ( 
.A(n_2607),
.Y(n_2713)
);

AOI22xp33_ASAP7_75t_L g2714 ( 
.A1(n_2629),
.A2(n_1167),
.B1(n_1168),
.B2(n_1165),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2558),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2542),
.Y(n_2716)
);

CKINVDCx20_ASAP7_75t_R g2717 ( 
.A(n_2616),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2615),
.Y(n_2718)
);

BUFx2_ASAP7_75t_L g2719 ( 
.A(n_2635),
.Y(n_2719)
);

INVx1_ASAP7_75t_SL g2720 ( 
.A(n_2635),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2649),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2641),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2643),
.A2(n_2539),
.B1(n_2607),
.B2(n_2551),
.Y(n_2723)
);

OAI21x1_ASAP7_75t_L g2724 ( 
.A1(n_2685),
.A2(n_2554),
.B(n_2545),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2669),
.B(n_2547),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_SL g2726 ( 
.A(n_2698),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2696),
.Y(n_2727)
);

AOI21xp5_ASAP7_75t_L g2728 ( 
.A1(n_2686),
.A2(n_2542),
.B(n_2551),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_SL g2729 ( 
.A(n_2690),
.B(n_2607),
.Y(n_2729)
);

AOI21x1_ASAP7_75t_L g2730 ( 
.A1(n_2709),
.A2(n_2619),
.B(n_2563),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2641),
.Y(n_2731)
);

AOI21xp5_ASAP7_75t_L g2732 ( 
.A1(n_2695),
.A2(n_2551),
.B(n_2560),
.Y(n_2732)
);

OA21x2_ASAP7_75t_L g2733 ( 
.A1(n_2664),
.A2(n_2559),
.B(n_2599),
.Y(n_2733)
);

OAI22xp5_ASAP7_75t_L g2734 ( 
.A1(n_2670),
.A2(n_2591),
.B1(n_2632),
.B2(n_2588),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2718),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2653),
.Y(n_2736)
);

AOI21xp5_ASAP7_75t_L g2737 ( 
.A1(n_2697),
.A2(n_2560),
.B(n_2536),
.Y(n_2737)
);

AO21x2_ASAP7_75t_L g2738 ( 
.A1(n_2664),
.A2(n_2544),
.B(n_2587),
.Y(n_2738)
);

OA21x2_ASAP7_75t_L g2739 ( 
.A1(n_2716),
.A2(n_2586),
.B(n_2595),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2645),
.Y(n_2740)
);

AOI21xp5_ASAP7_75t_L g2741 ( 
.A1(n_2694),
.A2(n_2621),
.B(n_2571),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2660),
.B(n_2614),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2662),
.B(n_2602),
.Y(n_2743)
);

AOI22xp33_ASAP7_75t_L g2744 ( 
.A1(n_2707),
.A2(n_2629),
.B1(n_2561),
.B2(n_2588),
.Y(n_2744)
);

HB1xp67_ASAP7_75t_L g2745 ( 
.A(n_2710),
.Y(n_2745)
);

AOI21xp5_ASAP7_75t_L g2746 ( 
.A1(n_2701),
.A2(n_2626),
.B(n_2636),
.Y(n_2746)
);

A2O1A1Ixp33_ASAP7_75t_L g2747 ( 
.A1(n_2678),
.A2(n_2613),
.B(n_2608),
.C(n_2603),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2651),
.Y(n_2748)
);

OAI21x1_ASAP7_75t_L g2749 ( 
.A1(n_2716),
.A2(n_2618),
.B(n_2578),
.Y(n_2749)
);

OAI21xp5_ASAP7_75t_L g2750 ( 
.A1(n_2712),
.A2(n_2561),
.B(n_2600),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2644),
.A2(n_2578),
.B(n_2569),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2656),
.B(n_2602),
.Y(n_2752)
);

NAND2x1_ASAP7_75t_L g2753 ( 
.A(n_2652),
.B(n_2590),
.Y(n_2753)
);

INVx2_ASAP7_75t_L g2754 ( 
.A(n_2655),
.Y(n_2754)
);

OAI22xp5_ASAP7_75t_L g2755 ( 
.A1(n_2681),
.A2(n_2591),
.B1(n_2556),
.B2(n_2535),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2688),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2650),
.B(n_2581),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_2719),
.Y(n_2758)
);

A2O1A1Ixp33_ASAP7_75t_L g2759 ( 
.A1(n_2665),
.A2(n_2623),
.B(n_2617),
.C(n_1300),
.Y(n_2759)
);

INVx5_ASAP7_75t_L g2760 ( 
.A(n_2702),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2689),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2691),
.B(n_2581),
.Y(n_2762)
);

OAI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2666),
.A2(n_2590),
.B(n_2569),
.Y(n_2763)
);

AOI21xp5_ASAP7_75t_L g2764 ( 
.A1(n_2699),
.A2(n_2704),
.B(n_2703),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2657),
.B(n_2535),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2661),
.Y(n_2766)
);

AOI221xp5_ASAP7_75t_L g2767 ( 
.A1(n_2714),
.A2(n_1305),
.B1(n_1306),
.B2(n_1302),
.C(n_1299),
.Y(n_2767)
);

AOI21xp5_ASAP7_75t_L g2768 ( 
.A1(n_2652),
.A2(n_2622),
.B(n_2535),
.Y(n_2768)
);

OR2x2_ASAP7_75t_L g2769 ( 
.A(n_2648),
.B(n_2622),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2658),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2675),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2646),
.B(n_2622),
.Y(n_2772)
);

INVx3_ASAP7_75t_L g2773 ( 
.A(n_2677),
.Y(n_2773)
);

BUFx8_ASAP7_75t_L g2774 ( 
.A(n_2698),
.Y(n_2774)
);

AND2x4_ASAP7_75t_L g2775 ( 
.A(n_2720),
.B(n_2),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2715),
.Y(n_2776)
);

OAI21xp5_ASAP7_75t_L g2777 ( 
.A1(n_2684),
.A2(n_1170),
.B(n_1169),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2640),
.B(n_1172),
.Y(n_2778)
);

OAI221xp5_ASAP7_75t_L g2779 ( 
.A1(n_2663),
.A2(n_1176),
.B1(n_1177),
.B2(n_1175),
.C(n_1173),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_2673),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2671),
.A2(n_1180),
.B1(n_1181),
.B2(n_1179),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2683),
.B(n_2541),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2673),
.Y(n_2783)
);

INVx4_ASAP7_75t_L g2784 ( 
.A(n_2654),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2677),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2687),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2687),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2706),
.B(n_1183),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2713),
.A2(n_1186),
.B(n_1185),
.Y(n_2789)
);

OA21x2_ASAP7_75t_L g2790 ( 
.A1(n_2659),
.A2(n_1188),
.B(n_1187),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2713),
.A2(n_1190),
.B(n_1189),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2679),
.B(n_2693),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2693),
.Y(n_2793)
);

OAI222xp33_ASAP7_75t_L g2794 ( 
.A1(n_2764),
.A2(n_2711),
.B1(n_2680),
.B2(n_2708),
.C1(n_2717),
.C2(n_2705),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_L g2795 ( 
.A1(n_2790),
.A2(n_2672),
.B1(n_2667),
.B2(n_2642),
.Y(n_2795)
);

AOI221xp5_ASAP7_75t_L g2796 ( 
.A1(n_2746),
.A2(n_1193),
.B1(n_1194),
.B2(n_1192),
.C(n_1191),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_L g2797 ( 
.A1(n_2790),
.A2(n_2667),
.B1(n_2676),
.B2(n_2642),
.Y(n_2797)
);

AOI22xp33_ASAP7_75t_L g2798 ( 
.A1(n_2741),
.A2(n_2676),
.B1(n_2682),
.B2(n_2693),
.Y(n_2798)
);

AOI22xp33_ASAP7_75t_SL g2799 ( 
.A1(n_2734),
.A2(n_2692),
.B1(n_2682),
.B2(n_2698),
.Y(n_2799)
);

OAI22xp33_ASAP7_75t_L g2800 ( 
.A1(n_2732),
.A2(n_2674),
.B1(n_2654),
.B2(n_2692),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2729),
.A2(n_2700),
.B1(n_2647),
.B2(n_2668),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2723),
.A2(n_2668),
.B1(n_1279),
.B2(n_1280),
.Y(n_2802)
);

AOI222xp33_ASAP7_75t_L g2803 ( 
.A1(n_2777),
.A2(n_1200),
.B1(n_1198),
.B2(n_1205),
.C1(n_1201),
.C2(n_1196),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2745),
.B(n_1197),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2758),
.B(n_3),
.Y(n_2805)
);

OAI22xp33_ASAP7_75t_L g2806 ( 
.A1(n_2737),
.A2(n_1210),
.B1(n_1212),
.B2(n_1208),
.Y(n_2806)
);

AOI22xp33_ASAP7_75t_L g2807 ( 
.A1(n_2750),
.A2(n_1310),
.B1(n_1221),
.B2(n_1223),
.Y(n_2807)
);

INVx4_ASAP7_75t_L g2808 ( 
.A(n_2784),
.Y(n_2808)
);

AOI221xp5_ASAP7_75t_L g2809 ( 
.A1(n_2779),
.A2(n_1227),
.B1(n_1228),
.B2(n_1224),
.C(n_1218),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2785),
.B(n_3),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2742),
.B(n_2776),
.Y(n_2811)
);

BUFx4f_ASAP7_75t_SL g2812 ( 
.A(n_2774),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2722),
.Y(n_2813)
);

BUFx4f_ASAP7_75t_SL g2814 ( 
.A(n_2774),
.Y(n_2814)
);

OAI221xp5_ASAP7_75t_L g2815 ( 
.A1(n_2744),
.A2(n_1237),
.B1(n_1238),
.B2(n_1235),
.C(n_1230),
.Y(n_2815)
);

AOI211xp5_ASAP7_75t_L g2816 ( 
.A1(n_2728),
.A2(n_1240),
.B(n_1243),
.C(n_1239),
.Y(n_2816)
);

HB1xp67_ASAP7_75t_L g2817 ( 
.A(n_2762),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_SL g2818 ( 
.A1(n_2755),
.A2(n_1244),
.B1(n_1248),
.B2(n_1241),
.Y(n_2818)
);

OAI21xp5_ASAP7_75t_L g2819 ( 
.A1(n_2747),
.A2(n_1252),
.B(n_1249),
.Y(n_2819)
);

CKINVDCx5p33_ASAP7_75t_R g2820 ( 
.A(n_2721),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2722),
.Y(n_2821)
);

OAI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2759),
.A2(n_1254),
.B1(n_1256),
.B2(n_1253),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2731),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2770),
.B(n_1257),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2771),
.B(n_1258),
.Y(n_2825)
);

AOI221xp5_ASAP7_75t_SL g2826 ( 
.A1(n_2751),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_2826)
);

AOI22xp33_ASAP7_75t_SL g2827 ( 
.A1(n_2784),
.A2(n_1262),
.B1(n_1265),
.B2(n_1261),
.Y(n_2827)
);

AOI22xp33_ASAP7_75t_L g2828 ( 
.A1(n_2767),
.A2(n_1290),
.B1(n_1291),
.B2(n_1289),
.Y(n_2828)
);

AOI22xp33_ASAP7_75t_L g2829 ( 
.A1(n_2740),
.A2(n_1307),
.B1(n_1293),
.B2(n_1269),
.Y(n_2829)
);

A2O1A1Ixp33_ASAP7_75t_L g2830 ( 
.A1(n_2789),
.A2(n_2791),
.B(n_2775),
.C(n_2788),
.Y(n_2830)
);

AOI22xp33_ASAP7_75t_SL g2831 ( 
.A1(n_2760),
.A2(n_1270),
.B1(n_1273),
.B2(n_1268),
.Y(n_2831)
);

AOI22xp33_ASAP7_75t_L g2832 ( 
.A1(n_2760),
.A2(n_1276),
.B1(n_1278),
.B2(n_1275),
.Y(n_2832)
);

AND2x4_ASAP7_75t_L g2833 ( 
.A(n_2786),
.B(n_4),
.Y(n_2833)
);

OR2x6_ASAP7_75t_L g2834 ( 
.A(n_2753),
.B(n_5),
.Y(n_2834)
);

OAI221xp5_ASAP7_75t_L g2835 ( 
.A1(n_2781),
.A2(n_1287),
.B1(n_1283),
.B2(n_1281),
.C(n_8),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2761),
.Y(n_2836)
);

INVx2_ASAP7_75t_SL g2837 ( 
.A(n_2760),
.Y(n_2837)
);

AOI22xp33_ASAP7_75t_L g2838 ( 
.A1(n_2775),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_2838)
);

NOR2xp33_ASAP7_75t_L g2839 ( 
.A(n_2726),
.B(n_9),
.Y(n_2839)
);

INVx2_ASAP7_75t_L g2840 ( 
.A(n_2813),
.Y(n_2840)
);

AND2x2_ASAP7_75t_L g2841 ( 
.A(n_2817),
.B(n_2769),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2837),
.B(n_2787),
.Y(n_2842)
);

BUFx2_ASAP7_75t_L g2843 ( 
.A(n_2808),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2836),
.B(n_2773),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2821),
.B(n_2773),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2823),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2798),
.B(n_2780),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2811),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2810),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_L g2850 ( 
.A(n_2805),
.B(n_2748),
.Y(n_2850)
);

BUFx3_ASAP7_75t_L g2851 ( 
.A(n_2812),
.Y(n_2851)
);

OR2x2_ASAP7_75t_L g2852 ( 
.A(n_2804),
.B(n_2752),
.Y(n_2852)
);

INVxp33_ASAP7_75t_SL g2853 ( 
.A(n_2820),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_2824),
.B(n_2727),
.Y(n_2854)
);

AND2x2_ASAP7_75t_L g2855 ( 
.A(n_2801),
.B(n_2783),
.Y(n_2855)
);

AOI22xp33_ASAP7_75t_SL g2856 ( 
.A1(n_2819),
.A2(n_2726),
.B1(n_2725),
.B2(n_2778),
.Y(n_2856)
);

BUFx3_ASAP7_75t_L g2857 ( 
.A(n_2814),
.Y(n_2857)
);

BUFx6f_ASAP7_75t_L g2858 ( 
.A(n_2808),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2825),
.B(n_2754),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2810),
.Y(n_2860)
);

OR2x2_ASAP7_75t_L g2861 ( 
.A(n_2800),
.B(n_2735),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2833),
.Y(n_2862)
);

AND2x2_ASAP7_75t_L g2863 ( 
.A(n_2799),
.B(n_2793),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2796),
.B(n_2736),
.Y(n_2864)
);

INVxp67_ASAP7_75t_L g2865 ( 
.A(n_2839),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2833),
.Y(n_2866)
);

OR2x2_ASAP7_75t_L g2867 ( 
.A(n_2834),
.B(n_2743),
.Y(n_2867)
);

AND2x2_ASAP7_75t_L g2868 ( 
.A(n_2834),
.B(n_2766),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2797),
.B(n_2756),
.Y(n_2869)
);

OR2x2_ASAP7_75t_L g2870 ( 
.A(n_2834),
.B(n_2772),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2806),
.Y(n_2871)
);

INVx2_ASAP7_75t_L g2872 ( 
.A(n_2815),
.Y(n_2872)
);

OR2x2_ASAP7_75t_L g2873 ( 
.A(n_2795),
.B(n_2761),
.Y(n_2873)
);

INVx1_ASAP7_75t_L g2874 ( 
.A(n_2816),
.Y(n_2874)
);

AND2x2_ASAP7_75t_L g2875 ( 
.A(n_2802),
.B(n_2763),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2830),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2842),
.B(n_2792),
.Y(n_2877)
);

INVx2_ASAP7_75t_L g2878 ( 
.A(n_2840),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_L g2879 ( 
.A1(n_2876),
.A2(n_2835),
.B1(n_2803),
.B2(n_2807),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2848),
.B(n_2826),
.Y(n_2880)
);

OR2x2_ASAP7_75t_L g2881 ( 
.A(n_2840),
.B(n_2757),
.Y(n_2881)
);

OR2x2_ASAP7_75t_L g2882 ( 
.A(n_2873),
.B(n_2765),
.Y(n_2882)
);

INVx2_ASAP7_75t_SL g2883 ( 
.A(n_2858),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2846),
.Y(n_2884)
);

INVxp67_ASAP7_75t_L g2885 ( 
.A(n_2873),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2846),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2843),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2844),
.Y(n_2888)
);

BUFx2_ASAP7_75t_L g2889 ( 
.A(n_2858),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2844),
.Y(n_2890)
);

AOI21xp5_ASAP7_75t_L g2891 ( 
.A1(n_2864),
.A2(n_2794),
.B(n_2822),
.Y(n_2891)
);

OA21x2_ASAP7_75t_L g2892 ( 
.A1(n_2869),
.A2(n_2768),
.B(n_2749),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2868),
.B(n_2818),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_SL g2894 ( 
.A(n_2858),
.B(n_2782),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2845),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2854),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2868),
.Y(n_2897)
);

INVxp67_ASAP7_75t_SL g2898 ( 
.A(n_2865),
.Y(n_2898)
);

AOI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2872),
.A2(n_2838),
.B(n_2832),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2845),
.Y(n_2900)
);

HB1xp67_ASAP7_75t_L g2901 ( 
.A(n_2841),
.Y(n_2901)
);

NOR2xp33_ASAP7_75t_L g2902 ( 
.A(n_2862),
.B(n_2831),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2859),
.Y(n_2903)
);

AO21x2_ASAP7_75t_L g2904 ( 
.A1(n_2863),
.A2(n_2730),
.B(n_2724),
.Y(n_2904)
);

INVx2_ASAP7_75t_L g2905 ( 
.A(n_2845),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2841),
.Y(n_2906)
);

INVxp67_ASAP7_75t_L g2907 ( 
.A(n_2867),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2842),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2849),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2849),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2860),
.Y(n_2911)
);

INVxp67_ASAP7_75t_L g2912 ( 
.A(n_2860),
.Y(n_2912)
);

AO31x2_ASAP7_75t_L g2913 ( 
.A1(n_2871),
.A2(n_2733),
.A3(n_2739),
.B(n_2738),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2850),
.Y(n_2914)
);

AOI21x1_ASAP7_75t_L g2915 ( 
.A1(n_2863),
.A2(n_2733),
.B(n_2739),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_2858),
.Y(n_2916)
);

INVx1_ASAP7_75t_SL g2917 ( 
.A(n_2887),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2909),
.Y(n_2918)
);

OR2x2_ASAP7_75t_L g2919 ( 
.A(n_2901),
.B(n_2852),
.Y(n_2919)
);

AOI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2891),
.A2(n_2874),
.B(n_2872),
.Y(n_2920)
);

OAI33xp33_ASAP7_75t_L g2921 ( 
.A1(n_2885),
.A2(n_2866),
.A3(n_2861),
.B1(n_2870),
.B2(n_2856),
.B3(n_12),
.Y(n_2921)
);

HB1xp67_ASAP7_75t_L g2922 ( 
.A(n_2898),
.Y(n_2922)
);

OR2x2_ASAP7_75t_L g2923 ( 
.A(n_2906),
.B(n_2847),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2909),
.Y(n_2924)
);

OR2x2_ASAP7_75t_L g2925 ( 
.A(n_2906),
.B(n_2847),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2902),
.B(n_2853),
.Y(n_2926)
);

NOR2x1_ASAP7_75t_L g2927 ( 
.A(n_2916),
.B(n_2851),
.Y(n_2927)
);

OR2x2_ASAP7_75t_L g2928 ( 
.A(n_2912),
.B(n_2875),
.Y(n_2928)
);

BUFx3_ASAP7_75t_L g2929 ( 
.A(n_2889),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2903),
.B(n_2855),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2911),
.Y(n_2931)
);

AND2x2_ASAP7_75t_L g2932 ( 
.A(n_2877),
.B(n_2855),
.Y(n_2932)
);

AOI22xp33_ASAP7_75t_L g2933 ( 
.A1(n_2896),
.A2(n_2875),
.B1(n_2857),
.B2(n_2851),
.Y(n_2933)
);

OAI22xp33_ASAP7_75t_L g2934 ( 
.A1(n_2880),
.A2(n_2907),
.B1(n_2882),
.B2(n_2897),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2914),
.B(n_2857),
.Y(n_2935)
);

INVx3_ASAP7_75t_L g2936 ( 
.A(n_2916),
.Y(n_2936)
);

OAI33xp33_ASAP7_75t_L g2937 ( 
.A1(n_2910),
.A2(n_12),
.A3(n_14),
.B1(n_10),
.B2(n_11),
.B3(n_13),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2877),
.B(n_2738),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_SL g2939 ( 
.A(n_2894),
.B(n_2853),
.Y(n_2939)
);

BUFx2_ASAP7_75t_L g2940 ( 
.A(n_2916),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2911),
.B(n_2829),
.Y(n_2941)
);

AOI221xp5_ASAP7_75t_L g2942 ( 
.A1(n_2899),
.A2(n_2809),
.B1(n_2828),
.B2(n_2827),
.C(n_14),
.Y(n_2942)
);

INVx4_ASAP7_75t_L g2943 ( 
.A(n_2883),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2908),
.B(n_10),
.Y(n_2944)
);

INVx1_ASAP7_75t_SL g2945 ( 
.A(n_2894),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2902),
.B(n_2893),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2895),
.B(n_11),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_SL g2948 ( 
.A(n_2883),
.B(n_15),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2895),
.B(n_15),
.Y(n_2949)
);

AND2x2_ASAP7_75t_L g2950 ( 
.A(n_2900),
.B(n_17),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2884),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2922),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2951),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2932),
.B(n_2900),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2929),
.B(n_2905),
.Y(n_2955)
);

AND2x2_ASAP7_75t_L g2956 ( 
.A(n_2917),
.B(n_2905),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2917),
.B(n_2920),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2946),
.B(n_2945),
.Y(n_2958)
);

AND2x2_ASAP7_75t_L g2959 ( 
.A(n_2927),
.B(n_2888),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_2945),
.B(n_2879),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2943),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2918),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_2943),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2934),
.B(n_2879),
.Y(n_2964)
);

INVx2_ASAP7_75t_L g2965 ( 
.A(n_2940),
.Y(n_2965)
);

AND2x2_ASAP7_75t_L g2966 ( 
.A(n_2936),
.B(n_2888),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2924),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2921),
.B(n_2881),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2936),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2931),
.Y(n_2970)
);

AND2x2_ASAP7_75t_L g2971 ( 
.A(n_2939),
.B(n_2890),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2947),
.B(n_2890),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2949),
.B(n_2950),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2933),
.B(n_2881),
.Y(n_2974)
);

OR2x2_ASAP7_75t_L g2975 ( 
.A(n_2919),
.B(n_2923),
.Y(n_2975)
);

OR2x2_ASAP7_75t_L g2976 ( 
.A(n_2925),
.B(n_2886),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2944),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_2926),
.B(n_2892),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2941),
.B(n_2878),
.Y(n_2979)
);

NAND2x1p5_ASAP7_75t_L g2980 ( 
.A(n_2948),
.B(n_2892),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2935),
.Y(n_2981)
);

NOR3xp33_ASAP7_75t_L g2982 ( 
.A(n_2942),
.B(n_2915),
.C(n_2878),
.Y(n_2982)
);

OR2x2_ASAP7_75t_L g2983 ( 
.A(n_2930),
.B(n_2913),
.Y(n_2983)
);

NOR2xp33_ASAP7_75t_R g2984 ( 
.A(n_2941),
.B(n_2935),
.Y(n_2984)
);

OR2x2_ASAP7_75t_L g2985 ( 
.A(n_2930),
.B(n_2913),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2928),
.Y(n_2986)
);

HB1xp67_ASAP7_75t_L g2987 ( 
.A(n_2938),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_2937),
.B(n_2904),
.Y(n_2988)
);

AND2x2_ASAP7_75t_L g2989 ( 
.A(n_2932),
.B(n_2892),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2922),
.Y(n_2990)
);

NOR3xp33_ASAP7_75t_L g2991 ( 
.A(n_2942),
.B(n_18),
.C(n_19),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2943),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2943),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2943),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2922),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2932),
.B(n_2904),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2932),
.B(n_2913),
.Y(n_2997)
);

OR2x2_ASAP7_75t_L g2998 ( 
.A(n_2922),
.B(n_2913),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2965),
.Y(n_2999)
);

XNOR2x2_ASAP7_75t_L g3000 ( 
.A(n_2988),
.B(n_21),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2965),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2955),
.B(n_2956),
.Y(n_3002)
);

INVx1_ASAP7_75t_SL g3003 ( 
.A(n_2984),
.Y(n_3003)
);

CKINVDCx5p33_ASAP7_75t_R g3004 ( 
.A(n_2984),
.Y(n_3004)
);

OR2x2_ASAP7_75t_L g3005 ( 
.A(n_2975),
.B(n_20),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2952),
.Y(n_3006)
);

NAND4xp75_ASAP7_75t_SL g3007 ( 
.A(n_2968),
.B(n_23),
.C(n_20),
.D(n_22),
.Y(n_3007)
);

BUFx3_ASAP7_75t_L g3008 ( 
.A(n_2961),
.Y(n_3008)
);

INVx1_ASAP7_75t_L g3009 ( 
.A(n_2990),
.Y(n_3009)
);

XOR2x1_ASAP7_75t_L g3010 ( 
.A(n_2961),
.B(n_23),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2995),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2968),
.B(n_24),
.Y(n_3012)
);

OR2x2_ASAP7_75t_L g3013 ( 
.A(n_2958),
.B(n_26),
.Y(n_3013)
);

NAND4xp75_ASAP7_75t_SL g3014 ( 
.A(n_2978),
.B(n_28),
.C(n_26),
.D(n_27),
.Y(n_3014)
);

NAND4xp75_ASAP7_75t_SL g3015 ( 
.A(n_2978),
.B(n_29),
.C(n_27),
.D(n_28),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2962),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2967),
.Y(n_3017)
);

NAND3xp33_ASAP7_75t_SL g3018 ( 
.A(n_2982),
.B(n_30),
.C(n_31),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2970),
.Y(n_3019)
);

NOR3xp33_ASAP7_75t_L g3020 ( 
.A(n_2964),
.B(n_30),
.C(n_31),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2954),
.B(n_33),
.Y(n_3021)
);

OAI22xp5_ASAP7_75t_L g3022 ( 
.A1(n_2960),
.A2(n_35),
.B1(n_36),
.B2(n_34),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2963),
.B(n_33),
.Y(n_3023)
);

NAND4xp75_ASAP7_75t_SL g3024 ( 
.A(n_2971),
.B(n_37),
.C(n_34),
.D(n_36),
.Y(n_3024)
);

INVxp67_ASAP7_75t_SL g3025 ( 
.A(n_2957),
.Y(n_3025)
);

XOR2x2_ASAP7_75t_L g3026 ( 
.A(n_2991),
.B(n_37),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2969),
.Y(n_3027)
);

XNOR2xp5_ASAP7_75t_L g3028 ( 
.A(n_2991),
.B(n_38),
.Y(n_3028)
);

INVx1_ASAP7_75t_SL g3029 ( 
.A(n_2959),
.Y(n_3029)
);

NAND4xp75_ASAP7_75t_L g3030 ( 
.A(n_2963),
.B(n_41),
.C(n_39),
.D(n_40),
.Y(n_3030)
);

OR2x2_ASAP7_75t_L g3031 ( 
.A(n_2981),
.B(n_2977),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2953),
.Y(n_3032)
);

NAND4xp75_ASAP7_75t_SL g3033 ( 
.A(n_2974),
.B(n_41),
.C(n_39),
.D(n_40),
.Y(n_3033)
);

AND2x2_ASAP7_75t_L g3034 ( 
.A(n_2992),
.B(n_42),
.Y(n_3034)
);

INVx3_ASAP7_75t_L g3035 ( 
.A(n_2969),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2992),
.B(n_2993),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2979),
.Y(n_3037)
);

AND4x1_ASAP7_75t_L g3038 ( 
.A(n_2982),
.B(n_45),
.C(n_42),
.D(n_44),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2993),
.B(n_44),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2994),
.Y(n_3040)
);

INVxp67_ASAP7_75t_L g3041 ( 
.A(n_2994),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2981),
.B(n_45),
.Y(n_3042)
);

AND2x2_ASAP7_75t_SL g3043 ( 
.A(n_2973),
.B(n_46),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2966),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2986),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2972),
.B(n_46),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2966),
.B(n_47),
.Y(n_3047)
);

NAND4xp75_ASAP7_75t_L g3048 ( 
.A(n_2996),
.B(n_51),
.C(n_48),
.D(n_50),
.Y(n_3048)
);

OR2x2_ASAP7_75t_L g3049 ( 
.A(n_2976),
.B(n_50),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2998),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2983),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2985),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2980),
.B(n_51),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2980),
.Y(n_3054)
);

NAND4xp75_ASAP7_75t_L g3055 ( 
.A(n_2989),
.B(n_54),
.C(n_52),
.D(n_53),
.Y(n_3055)
);

XNOR2xp5_ASAP7_75t_L g3056 ( 
.A(n_2997),
.B(n_52),
.Y(n_3056)
);

NAND4xp75_ASAP7_75t_SL g3057 ( 
.A(n_2987),
.B(n_56),
.C(n_54),
.D(n_55),
.Y(n_3057)
);

INVx1_ASAP7_75t_L g3058 ( 
.A(n_2987),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2969),
.Y(n_3059)
);

NAND4xp75_ASAP7_75t_L g3060 ( 
.A(n_2988),
.B(n_60),
.C(n_57),
.D(n_58),
.Y(n_3060)
);

XOR2x2_ASAP7_75t_L g3061 ( 
.A(n_2991),
.B(n_58),
.Y(n_3061)
);

AND2x4_ASAP7_75t_L g3062 ( 
.A(n_2965),
.B(n_61),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2965),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2965),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_2965),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_2965),
.B(n_62),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_3010),
.B(n_62),
.Y(n_3067)
);

INVx1_ASAP7_75t_SL g3068 ( 
.A(n_3003),
.Y(n_3068)
);

AOI21xp33_ASAP7_75t_L g3069 ( 
.A1(n_3012),
.A2(n_63),
.B(n_64),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_3002),
.B(n_63),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_3058),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_3058),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_3065),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_3064),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_3043),
.B(n_64),
.Y(n_3075)
);

INVx1_ASAP7_75t_SL g3076 ( 
.A(n_3004),
.Y(n_3076)
);

OR2x2_ASAP7_75t_L g3077 ( 
.A(n_3044),
.B(n_65),
.Y(n_3077)
);

AOI22xp33_ASAP7_75t_SL g3078 ( 
.A1(n_3000),
.A2(n_789),
.B1(n_792),
.B2(n_788),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2999),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_3029),
.B(n_788),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_3064),
.B(n_65),
.Y(n_3081)
);

OR2x2_ASAP7_75t_L g3082 ( 
.A(n_3036),
.B(n_67),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_3008),
.B(n_3038),
.Y(n_3083)
);

OR2x2_ASAP7_75t_L g3084 ( 
.A(n_3005),
.B(n_67),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_3021),
.B(n_793),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_L g3086 ( 
.A(n_3025),
.B(n_68),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_3035),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_3013),
.B(n_69),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_3041),
.B(n_69),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2999),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_3001),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_3040),
.B(n_796),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_3056),
.B(n_70),
.Y(n_3093)
);

OR2x2_ASAP7_75t_L g3094 ( 
.A(n_3018),
.B(n_70),
.Y(n_3094)
);

INVxp67_ASAP7_75t_L g3095 ( 
.A(n_3055),
.Y(n_3095)
);

INVxp33_ASAP7_75t_L g3096 ( 
.A(n_3020),
.Y(n_3096)
);

INVx2_ASAP7_75t_L g3097 ( 
.A(n_3035),
.Y(n_3097)
);

OR2x2_ASAP7_75t_L g3098 ( 
.A(n_3031),
.B(n_71),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_3034),
.B(n_71),
.Y(n_3099)
);

CKINVDCx16_ASAP7_75t_R g3100 ( 
.A(n_3028),
.Y(n_3100)
);

NAND3xp33_ASAP7_75t_L g3101 ( 
.A(n_3054),
.B(n_72),
.C(n_73),
.Y(n_3101)
);

INVx2_ASAP7_75t_L g3102 ( 
.A(n_3062),
.Y(n_3102)
);

OR2x2_ASAP7_75t_L g3103 ( 
.A(n_3045),
.B(n_73),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_3001),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_3062),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_3039),
.B(n_74),
.Y(n_3106)
);

NOR2x1_ASAP7_75t_L g3107 ( 
.A(n_3048),
.B(n_75),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_3053),
.B(n_75),
.Y(n_3108)
);

OR2x2_ASAP7_75t_L g3109 ( 
.A(n_3063),
.B(n_76),
.Y(n_3109)
);

INVx2_ASAP7_75t_SL g3110 ( 
.A(n_3063),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_3042),
.Y(n_3111)
);

OR2x2_ASAP7_75t_L g3112 ( 
.A(n_3047),
.B(n_76),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_3027),
.B(n_77),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_3059),
.Y(n_3114)
);

AND2x2_ASAP7_75t_L g3115 ( 
.A(n_3037),
.B(n_77),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_3049),
.Y(n_3116)
);

NAND3xp33_ASAP7_75t_L g3117 ( 
.A(n_3006),
.B(n_79),
.C(n_80),
.Y(n_3117)
);

OAI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_3060),
.A2(n_79),
.B(n_81),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3026),
.Y(n_3119)
);

OR2x2_ASAP7_75t_L g3120 ( 
.A(n_3009),
.B(n_81),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_3011),
.B(n_82),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_3046),
.B(n_787),
.Y(n_3122)
);

INVxp67_ASAP7_75t_SL g3123 ( 
.A(n_3066),
.Y(n_3123)
);

INVx2_ASAP7_75t_L g3124 ( 
.A(n_3023),
.Y(n_3124)
);

HB1xp67_ASAP7_75t_L g3125 ( 
.A(n_3050),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_3016),
.Y(n_3126)
);

AND2x2_ASAP7_75t_L g3127 ( 
.A(n_3032),
.B(n_3017),
.Y(n_3127)
);

INVx2_ASAP7_75t_L g3128 ( 
.A(n_3030),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_3061),
.B(n_82),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_3022),
.B(n_83),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_3019),
.B(n_84),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_3051),
.B(n_793),
.Y(n_3132)
);

INVxp67_ASAP7_75t_SL g3133 ( 
.A(n_3052),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_3007),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_L g3135 ( 
.A1(n_3014),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.Y(n_3135)
);

BUFx2_ASAP7_75t_L g3136 ( 
.A(n_3015),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3057),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_3033),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_3024),
.B(n_796),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_3002),
.B(n_86),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_3004),
.B(n_87),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_3002),
.B(n_88),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_3058),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_3058),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_3058),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_3002),
.B(n_88),
.Y(n_3146)
);

OAI22xp33_ASAP7_75t_L g3147 ( 
.A1(n_3012),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.Y(n_3147)
);

INVxp33_ASAP7_75t_L g3148 ( 
.A(n_3002),
.Y(n_3148)
);

INVxp67_ASAP7_75t_L g3149 ( 
.A(n_3065),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_3003),
.B(n_93),
.Y(n_3150)
);

OR2x2_ASAP7_75t_L g3151 ( 
.A(n_3003),
.B(n_93),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_3002),
.B(n_94),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_3002),
.B(n_94),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_3058),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_3058),
.Y(n_3155)
);

AOI32xp33_ASAP7_75t_L g3156 ( 
.A1(n_3003),
.A2(n_97),
.A3(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_3156)
);

INVx3_ASAP7_75t_L g3157 ( 
.A(n_3064),
.Y(n_3157)
);

CKINVDCx16_ASAP7_75t_R g3158 ( 
.A(n_3003),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3064),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_3002),
.B(n_785),
.Y(n_3160)
);

NOR2xp33_ASAP7_75t_L g3161 ( 
.A(n_3158),
.B(n_95),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3074),
.Y(n_3162)
);

NAND3xp33_ASAP7_75t_SL g3163 ( 
.A(n_3078),
.B(n_98),
.C(n_99),
.Y(n_3163)
);

OAI21xp33_ASAP7_75t_L g3164 ( 
.A1(n_3148),
.A2(n_99),
.B(n_100),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_3074),
.Y(n_3165)
);

OAI21xp33_ASAP7_75t_SL g3166 ( 
.A1(n_3073),
.A2(n_101),
.B(n_102),
.Y(n_3166)
);

O2A1O1Ixp33_ASAP7_75t_SL g3167 ( 
.A1(n_3067),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_3167)
);

OAI22xp33_ASAP7_75t_L g3168 ( 
.A1(n_3096),
.A2(n_107),
.B1(n_105),
.B2(n_106),
.Y(n_3168)
);

HB1xp67_ASAP7_75t_L g3169 ( 
.A(n_3157),
.Y(n_3169)
);

OAI22xp5_ASAP7_75t_L g3170 ( 
.A1(n_3100),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3073),
.Y(n_3171)
);

OAI31xp33_ASAP7_75t_L g3172 ( 
.A1(n_3147),
.A2(n_111),
.A3(n_109),
.B(n_110),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_3157),
.Y(n_3173)
);

OAI31xp33_ASAP7_75t_SL g3174 ( 
.A1(n_3107),
.A2(n_114),
.A3(n_110),
.B(n_112),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_3071),
.Y(n_3175)
);

OAI22xp5_ASAP7_75t_SL g3176 ( 
.A1(n_3136),
.A2(n_117),
.B1(n_112),
.B2(n_116),
.Y(n_3176)
);

AOI22xp33_ASAP7_75t_L g3177 ( 
.A1(n_3119),
.A2(n_119),
.B1(n_116),
.B2(n_118),
.Y(n_3177)
);

INVx2_ASAP7_75t_L g3178 ( 
.A(n_3159),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_3068),
.B(n_121),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_3083),
.A2(n_3118),
.B(n_3119),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3071),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_3072),
.Y(n_3182)
);

INVx3_ASAP7_75t_L g3183 ( 
.A(n_3087),
.Y(n_3183)
);

OAI221xp5_ASAP7_75t_L g3184 ( 
.A1(n_3095),
.A2(n_124),
.B1(n_121),
.B2(n_122),
.C(n_125),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3072),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_3144),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_3102),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_3135),
.A2(n_128),
.B1(n_125),
.B2(n_126),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_3144),
.Y(n_3189)
);

OAI22xp33_ASAP7_75t_L g3190 ( 
.A1(n_3094),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_3190)
);

AOI22xp5_ASAP7_75t_L g3191 ( 
.A1(n_3128),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_3191)
);

AOI211xp5_ASAP7_75t_L g3192 ( 
.A1(n_3069),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_3192)
);

AOI22xp5_ASAP7_75t_L g3193 ( 
.A1(n_3076),
.A2(n_135),
.B1(n_133),
.B2(n_134),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3090),
.Y(n_3194)
);

OAI21xp5_ASAP7_75t_L g3195 ( 
.A1(n_3149),
.A2(n_134),
.B(n_136),
.Y(n_3195)
);

BUFx2_ASAP7_75t_L g3196 ( 
.A(n_3105),
.Y(n_3196)
);

INVxp67_ASAP7_75t_L g3197 ( 
.A(n_3075),
.Y(n_3197)
);

OAI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_3134),
.A2(n_140),
.B1(n_136),
.B2(n_139),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3090),
.Y(n_3199)
);

OAI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3101),
.A2(n_139),
.B(n_142),
.Y(n_3200)
);

AOI21xp33_ASAP7_75t_SL g3201 ( 
.A1(n_3150),
.A2(n_142),
.B(n_143),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3110),
.Y(n_3202)
);

NOR3xp33_ASAP7_75t_L g3203 ( 
.A(n_3123),
.B(n_144),
.C(n_146),
.Y(n_3203)
);

AOI22xp5_ASAP7_75t_L g3204 ( 
.A1(n_3137),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3125),
.Y(n_3205)
);

OAI221xp5_ASAP7_75t_L g3206 ( 
.A1(n_3156),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_151),
.Y(n_3206)
);

O2A1O1Ixp33_ASAP7_75t_L g3207 ( 
.A1(n_3086),
.A2(n_151),
.B(n_149),
.C(n_150),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3143),
.Y(n_3208)
);

OAI21xp33_ASAP7_75t_L g3209 ( 
.A1(n_3111),
.A2(n_3133),
.B(n_3116),
.Y(n_3209)
);

AND2x4_ASAP7_75t_L g3210 ( 
.A(n_3097),
.B(n_152),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_3145),
.Y(n_3211)
);

NAND3xp33_ASAP7_75t_L g3212 ( 
.A(n_3111),
.B(n_153),
.C(n_154),
.Y(n_3212)
);

XOR2x2_ASAP7_75t_L g3213 ( 
.A(n_3129),
.B(n_154),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_3154),
.Y(n_3214)
);

OAI31xp33_ASAP7_75t_L g3215 ( 
.A1(n_3117),
.A2(n_157),
.A3(n_155),
.B(n_156),
.Y(n_3215)
);

AOI21xp33_ASAP7_75t_SL g3216 ( 
.A1(n_3151),
.A2(n_156),
.B(n_157),
.Y(n_3216)
);

HB1xp67_ASAP7_75t_L g3217 ( 
.A(n_3080),
.Y(n_3217)
);

INVx2_ASAP7_75t_L g3218 ( 
.A(n_3070),
.Y(n_3218)
);

OAI22xp33_ASAP7_75t_SL g3219 ( 
.A1(n_3155),
.A2(n_794),
.B1(n_160),
.B2(n_158),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_3140),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3079),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3142),
.B(n_158),
.Y(n_3222)
);

INVx1_ASAP7_75t_L g3223 ( 
.A(n_3091),
.Y(n_3223)
);

OAI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_3130),
.A2(n_159),
.B(n_161),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3104),
.Y(n_3225)
);

OAI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_3081),
.A2(n_162),
.B(n_163),
.Y(n_3226)
);

AOI22xp5_ASAP7_75t_L g3227 ( 
.A1(n_3138),
.A2(n_3146),
.B1(n_3153),
.B2(n_3152),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3085),
.Y(n_3228)
);

AO21x1_ASAP7_75t_L g3229 ( 
.A1(n_3141),
.A2(n_164),
.B(n_163),
.Y(n_3229)
);

INVx2_ASAP7_75t_L g3230 ( 
.A(n_3160),
.Y(n_3230)
);

AOI21xp33_ASAP7_75t_L g3231 ( 
.A1(n_3124),
.A2(n_162),
.B(n_166),
.Y(n_3231)
);

NAND4xp25_ASAP7_75t_SL g3232 ( 
.A(n_3093),
.B(n_168),
.C(n_166),
.D(n_167),
.Y(n_3232)
);

OAI32xp33_ASAP7_75t_L g3233 ( 
.A1(n_3126),
.A2(n_170),
.A3(n_172),
.B1(n_169),
.B2(n_171),
.Y(n_3233)
);

AOI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3132),
.A2(n_170),
.B1(n_168),
.B2(n_169),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3099),
.Y(n_3235)
);

NOR3xp33_ASAP7_75t_L g3236 ( 
.A(n_3114),
.B(n_171),
.C(n_173),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3092),
.Y(n_3237)
);

OAI21xp33_ASAP7_75t_SL g3238 ( 
.A1(n_3127),
.A2(n_3089),
.B(n_3098),
.Y(n_3238)
);

NAND2x1p5_ASAP7_75t_L g3239 ( 
.A(n_3084),
.B(n_173),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3113),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3109),
.Y(n_3241)
);

INVxp67_ASAP7_75t_SL g3242 ( 
.A(n_3108),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3122),
.B(n_174),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3121),
.A2(n_176),
.B(n_177),
.Y(n_3244)
);

INVxp67_ASAP7_75t_SL g3245 ( 
.A(n_3106),
.Y(n_3245)
);

OAI21xp33_ASAP7_75t_L g3246 ( 
.A1(n_3131),
.A2(n_177),
.B(n_178),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3077),
.Y(n_3247)
);

AOI22xp5_ASAP7_75t_L g3248 ( 
.A1(n_3115),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_3248)
);

NAND2xp5_ASAP7_75t_L g3249 ( 
.A(n_3088),
.B(n_179),
.Y(n_3249)
);

O2A1O1Ixp5_ASAP7_75t_L g3250 ( 
.A1(n_3082),
.A2(n_3103),
.B(n_3120),
.C(n_3139),
.Y(n_3250)
);

OAI211xp5_ASAP7_75t_SL g3251 ( 
.A1(n_3112),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_3251)
);

AOI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_3158),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_3252)
);

OAI221xp5_ASAP7_75t_SL g3253 ( 
.A1(n_3078),
.A2(n_200),
.B1(n_210),
.B2(n_192),
.C(n_183),
.Y(n_3253)
);

INVx3_ASAP7_75t_L g3254 ( 
.A(n_3157),
.Y(n_3254)
);

AOI22xp5_ASAP7_75t_L g3255 ( 
.A1(n_3158),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_3255)
);

NAND2x1_ASAP7_75t_L g3256 ( 
.A(n_3157),
.B(n_786),
.Y(n_3256)
);

AOI22xp33_ASAP7_75t_L g3257 ( 
.A1(n_3096),
.A2(n_188),
.B1(n_186),
.B2(n_187),
.Y(n_3257)
);

AOI22xp5_ASAP7_75t_L g3258 ( 
.A1(n_3158),
.A2(n_192),
.B1(n_189),
.B2(n_191),
.Y(n_3258)
);

AOI22xp5_ASAP7_75t_SL g3259 ( 
.A1(n_3118),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_3259)
);

AOI21xp5_ASAP7_75t_L g3260 ( 
.A1(n_3096),
.A2(n_193),
.B(n_195),
.Y(n_3260)
);

AO21x1_ASAP7_75t_L g3261 ( 
.A1(n_3067),
.A2(n_198),
.B(n_197),
.Y(n_3261)
);

XOR2x2_ASAP7_75t_L g3262 ( 
.A(n_3107),
.B(n_196),
.Y(n_3262)
);

OAI22xp33_ASAP7_75t_SL g3263 ( 
.A1(n_3158),
.A2(n_199),
.B1(n_196),
.B2(n_198),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3074),
.Y(n_3264)
);

AOI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_3158),
.A2(n_202),
.B1(n_199),
.B2(n_201),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3074),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3074),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3074),
.Y(n_3268)
);

OAI211xp5_ASAP7_75t_SL g3269 ( 
.A1(n_3076),
.A2(n_203),
.B(n_201),
.C(n_202),
.Y(n_3269)
);

INVx1_ASAP7_75t_SL g3270 ( 
.A(n_3158),
.Y(n_3270)
);

AOI211xp5_ASAP7_75t_L g3271 ( 
.A1(n_3096),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3074),
.Y(n_3272)
);

INVx3_ASAP7_75t_L g3273 ( 
.A(n_3157),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3100),
.B(n_205),
.Y(n_3274)
);

INVx1_ASAP7_75t_L g3275 ( 
.A(n_3074),
.Y(n_3275)
);

OAI211xp5_ASAP7_75t_L g3276 ( 
.A1(n_3078),
.A2(n_211),
.B(n_206),
.C(n_208),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3074),
.Y(n_3277)
);

XNOR2x2_ASAP7_75t_L g3278 ( 
.A(n_3107),
.B(n_208),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_L g3279 ( 
.A1(n_3096),
.A2(n_215),
.B1(n_211),
.B2(n_214),
.Y(n_3279)
);

OAI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3078),
.A2(n_215),
.B(n_216),
.Y(n_3280)
);

OAI21xp5_ASAP7_75t_SL g3281 ( 
.A1(n_3078),
.A2(n_216),
.B(n_218),
.Y(n_3281)
);

INVx2_ASAP7_75t_L g3282 ( 
.A(n_3157),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3074),
.Y(n_3283)
);

AOI21xp33_ASAP7_75t_L g3284 ( 
.A1(n_3148),
.A2(n_219),
.B(n_220),
.Y(n_3284)
);

OAI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_3096),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_3285)
);

INVx2_ASAP7_75t_SL g3286 ( 
.A(n_3157),
.Y(n_3286)
);

OAI22xp33_ASAP7_75t_SL g3287 ( 
.A1(n_3158),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_3287)
);

BUFx2_ASAP7_75t_SL g3288 ( 
.A(n_3157),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3074),
.Y(n_3289)
);

OAI21xp5_ASAP7_75t_L g3290 ( 
.A1(n_3078),
.A2(n_224),
.B(n_225),
.Y(n_3290)
);

AOI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_3158),
.A2(n_226),
.B1(n_224),
.B2(n_225),
.Y(n_3291)
);

XOR2x2_ASAP7_75t_L g3292 ( 
.A(n_3107),
.B(n_227),
.Y(n_3292)
);

INVx6_ASAP7_75t_L g3293 ( 
.A(n_3158),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3074),
.Y(n_3294)
);

AOI21xp5_ASAP7_75t_L g3295 ( 
.A1(n_3096),
.A2(n_228),
.B(n_230),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_3158),
.B(n_231),
.Y(n_3296)
);

XNOR2xp5_ASAP7_75t_L g3297 ( 
.A(n_3148),
.B(n_231),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3158),
.B(n_232),
.Y(n_3298)
);

AOI21xp33_ASAP7_75t_SL g3299 ( 
.A1(n_3158),
.A2(n_233),
.B(n_234),
.Y(n_3299)
);

NAND3x1_ASAP7_75t_L g3300 ( 
.A(n_3107),
.B(n_235),
.C(n_236),
.Y(n_3300)
);

NOR2x1_ASAP7_75t_SL g3301 ( 
.A(n_3102),
.B(n_236),
.Y(n_3301)
);

A2O1A1Ixp33_ASAP7_75t_L g3302 ( 
.A1(n_3078),
.A2(n_238),
.B(n_235),
.C(n_237),
.Y(n_3302)
);

NAND2xp5_ASAP7_75t_SL g3303 ( 
.A(n_3158),
.B(n_237),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3158),
.B(n_239),
.Y(n_3304)
);

OAI211xp5_ASAP7_75t_SL g3305 ( 
.A1(n_3076),
.A2(n_241),
.B(n_239),
.C(n_240),
.Y(n_3305)
);

AND2x2_ASAP7_75t_L g3306 ( 
.A(n_3158),
.B(n_241),
.Y(n_3306)
);

INVx2_ASAP7_75t_SL g3307 ( 
.A(n_3157),
.Y(n_3307)
);

INVx1_ASAP7_75t_SL g3308 ( 
.A(n_3158),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3074),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3074),
.Y(n_3310)
);

BUFx3_ASAP7_75t_L g3311 ( 
.A(n_3102),
.Y(n_3311)
);

OAI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3096),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3074),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3158),
.B(n_242),
.Y(n_3314)
);

BUFx2_ASAP7_75t_SL g3315 ( 
.A(n_3157),
.Y(n_3315)
);

OAI221xp5_ASAP7_75t_L g3316 ( 
.A1(n_3078),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.C(n_247),
.Y(n_3316)
);

NAND3xp33_ASAP7_75t_L g3317 ( 
.A(n_3078),
.B(n_245),
.C(n_248),
.Y(n_3317)
);

AO21x1_ASAP7_75t_L g3318 ( 
.A1(n_3263),
.A2(n_248),
.B(n_249),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3270),
.B(n_249),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_L g3320 ( 
.A1(n_3308),
.A2(n_250),
.B(n_251),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3169),
.Y(n_3321)
);

AOI221xp5_ASAP7_75t_L g3322 ( 
.A1(n_3180),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.C(n_253),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3306),
.B(n_252),
.Y(n_3323)
);

INVx1_ASAP7_75t_SL g3324 ( 
.A(n_3293),
.Y(n_3324)
);

AOI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_3269),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_3325)
);

OAI221xp5_ASAP7_75t_L g3326 ( 
.A1(n_3174),
.A2(n_257),
.B1(n_254),
.B2(n_256),
.C(n_258),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_3293),
.Y(n_3327)
);

OAI32xp33_ASAP7_75t_L g3328 ( 
.A1(n_3305),
.A2(n_259),
.A3(n_257),
.B1(n_258),
.B2(n_260),
.Y(n_3328)
);

NAND3xp33_ASAP7_75t_L g3329 ( 
.A(n_3205),
.B(n_259),
.C(n_260),
.Y(n_3329)
);

OAI221xp5_ASAP7_75t_L g3330 ( 
.A1(n_3209),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.C(n_265),
.Y(n_3330)
);

AOI211xp5_ASAP7_75t_L g3331 ( 
.A1(n_3163),
.A2(n_3253),
.B(n_3287),
.C(n_3281),
.Y(n_3331)
);

INVx2_ASAP7_75t_SL g3332 ( 
.A(n_3256),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3301),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3196),
.Y(n_3334)
);

NOR2x1p5_ASAP7_75t_L g3335 ( 
.A(n_3296),
.B(n_261),
.Y(n_3335)
);

AOI21xp33_ASAP7_75t_SL g3336 ( 
.A1(n_3303),
.A2(n_262),
.B(n_265),
.Y(n_3336)
);

NAND2xp33_ASAP7_75t_SL g3337 ( 
.A(n_3176),
.B(n_267),
.Y(n_3337)
);

OAI221xp5_ASAP7_75t_L g3338 ( 
.A1(n_3280),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.C(n_270),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_3217),
.Y(n_3339)
);

OAI22xp33_ASAP7_75t_L g3340 ( 
.A1(n_3317),
.A2(n_273),
.B1(n_270),
.B2(n_271),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3311),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3274),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3239),
.Y(n_3343)
);

O2A1O1Ixp33_ASAP7_75t_SL g3344 ( 
.A1(n_3302),
.A2(n_274),
.B(n_271),
.C(n_273),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3161),
.B(n_274),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3218),
.B(n_275),
.Y(n_3346)
);

AOI211xp5_ASAP7_75t_SL g3347 ( 
.A1(n_3202),
.A2(n_278),
.B(n_275),
.C(n_276),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3298),
.Y(n_3348)
);

AOI21xp5_ASAP7_75t_L g3349 ( 
.A1(n_3290),
.A2(n_276),
.B(n_278),
.Y(n_3349)
);

NOR2xp33_ASAP7_75t_L g3350 ( 
.A(n_3304),
.B(n_279),
.Y(n_3350)
);

AOI222xp33_ASAP7_75t_L g3351 ( 
.A1(n_3238),
.A2(n_3262),
.B1(n_3292),
.B2(n_3197),
.C1(n_3166),
.C2(n_3200),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3286),
.B(n_279),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3314),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_3254),
.Y(n_3354)
);

OAI31xp33_ASAP7_75t_SL g3355 ( 
.A1(n_3276),
.A2(n_282),
.A3(n_280),
.B(n_281),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3307),
.B(n_280),
.Y(n_3356)
);

AOI22xp33_ASAP7_75t_L g3357 ( 
.A1(n_3220),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_3357)
);

OAI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_3300),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3254),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3273),
.Y(n_3360)
);

OAI321xp33_ASAP7_75t_L g3361 ( 
.A1(n_3187),
.A2(n_288),
.A3(n_290),
.B1(n_286),
.B2(n_287),
.C(n_289),
.Y(n_3361)
);

INVxp67_ASAP7_75t_L g3362 ( 
.A(n_3288),
.Y(n_3362)
);

OA22x2_ASAP7_75t_L g3363 ( 
.A1(n_3227),
.A2(n_3315),
.B1(n_3173),
.B2(n_3282),
.Y(n_3363)
);

AOI22xp33_ASAP7_75t_L g3364 ( 
.A1(n_3230),
.A2(n_290),
.B1(n_287),
.B2(n_289),
.Y(n_3364)
);

A2O1A1Ixp33_ASAP7_75t_L g3365 ( 
.A1(n_3207),
.A2(n_3259),
.B(n_3215),
.C(n_3299),
.Y(n_3365)
);

HB1xp67_ASAP7_75t_L g3366 ( 
.A(n_3273),
.Y(n_3366)
);

AOI21xp5_ASAP7_75t_L g3367 ( 
.A1(n_3167),
.A2(n_291),
.B(n_292),
.Y(n_3367)
);

OAI222xp33_ASAP7_75t_L g3368 ( 
.A1(n_3316),
.A2(n_3206),
.B1(n_3178),
.B2(n_3228),
.C1(n_3241),
.C2(n_3183),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3183),
.B(n_291),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3201),
.B(n_292),
.Y(n_3370)
);

AOI21xp5_ASAP7_75t_L g3371 ( 
.A1(n_3260),
.A2(n_293),
.B(n_294),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_3216),
.B(n_293),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_3179),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3243),
.Y(n_3374)
);

AO21x1_ASAP7_75t_L g3375 ( 
.A1(n_3175),
.A2(n_294),
.B(n_295),
.Y(n_3375)
);

OAI22xp5_ASAP7_75t_L g3376 ( 
.A1(n_3177),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3181),
.Y(n_3377)
);

OAI22xp5_ASAP7_75t_L g3378 ( 
.A1(n_3252),
.A2(n_3255),
.B1(n_3265),
.B2(n_3258),
.Y(n_3378)
);

AND2x2_ASAP7_75t_L g3379 ( 
.A(n_3235),
.B(n_297),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3182),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3237),
.B(n_299),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_3240),
.B(n_299),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3185),
.Y(n_3383)
);

NAND4xp25_ASAP7_75t_L g3384 ( 
.A(n_3250),
.B(n_302),
.C(n_300),
.D(n_301),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3186),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3291),
.B(n_302),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3210),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3189),
.Y(n_3388)
);

OAI31xp33_ASAP7_75t_L g3389 ( 
.A1(n_3251),
.A2(n_3219),
.A3(n_3285),
.B(n_3168),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3210),
.B(n_304),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_3295),
.B(n_305),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3224),
.A2(n_305),
.B(n_306),
.Y(n_3392)
);

INVx1_ASAP7_75t_SL g3393 ( 
.A(n_3278),
.Y(n_3393)
);

OAI32xp33_ASAP7_75t_L g3394 ( 
.A1(n_3171),
.A2(n_308),
.A3(n_306),
.B1(n_307),
.B2(n_309),
.Y(n_3394)
);

INVx1_ASAP7_75t_SL g3395 ( 
.A(n_3297),
.Y(n_3395)
);

OR2x2_ASAP7_75t_L g3396 ( 
.A(n_3247),
.B(n_307),
.Y(n_3396)
);

INVx3_ASAP7_75t_L g3397 ( 
.A(n_3162),
.Y(n_3397)
);

OAI321xp33_ASAP7_75t_L g3398 ( 
.A1(n_3208),
.A2(n_310),
.A3(n_312),
.B1(n_308),
.B2(n_309),
.C(n_311),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3236),
.B(n_310),
.Y(n_3399)
);

XOR2x2_ASAP7_75t_L g3400 ( 
.A(n_3213),
.B(n_3188),
.Y(n_3400)
);

NOR2xp33_ASAP7_75t_L g3401 ( 
.A(n_3164),
.B(n_311),
.Y(n_3401)
);

AOI322xp5_ASAP7_75t_L g3402 ( 
.A1(n_3203),
.A2(n_318),
.A3(n_317),
.B1(n_315),
.B2(n_312),
.C1(n_313),
.C2(n_316),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3222),
.Y(n_3403)
);

AND2x2_ASAP7_75t_L g3404 ( 
.A(n_3242),
.B(n_313),
.Y(n_3404)
);

OAI22xp5_ASAP7_75t_L g3405 ( 
.A1(n_3257),
.A2(n_319),
.B1(n_315),
.B2(n_316),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_SL g3406 ( 
.A(n_3229),
.B(n_3261),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_3195),
.A2(n_3190),
.B(n_3244),
.Y(n_3407)
);

OAI222xp33_ASAP7_75t_L g3408 ( 
.A1(n_3193),
.A2(n_322),
.B1(n_324),
.B2(n_320),
.C1(n_321),
.C2(n_323),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3245),
.B(n_320),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3194),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3271),
.B(n_3192),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_L g3412 ( 
.A(n_3172),
.B(n_321),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3246),
.B(n_322),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3312),
.B(n_323),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3191),
.B(n_324),
.Y(n_3415)
);

OAI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_3212),
.A2(n_326),
.B(n_328),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3170),
.B(n_328),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3199),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3165),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_3264),
.Y(n_3420)
);

OAI22xp33_ASAP7_75t_SL g3421 ( 
.A1(n_3266),
.A2(n_332),
.B1(n_329),
.B2(n_330),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3267),
.Y(n_3422)
);

AOI21xp33_ASAP7_75t_L g3423 ( 
.A1(n_3268),
.A2(n_329),
.B(n_330),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3272),
.Y(n_3424)
);

INVx2_ASAP7_75t_SL g3425 ( 
.A(n_3275),
.Y(n_3425)
);

OAI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_3204),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3426)
);

HB1xp67_ASAP7_75t_L g3427 ( 
.A(n_3277),
.Y(n_3427)
);

OR2x2_ASAP7_75t_L g3428 ( 
.A(n_3249),
.B(n_335),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3279),
.B(n_337),
.Y(n_3429)
);

AOI21xp33_ASAP7_75t_SL g3430 ( 
.A1(n_3284),
.A2(n_338),
.B(n_339),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_L g3431 ( 
.A1(n_3313),
.A2(n_342),
.B1(n_338),
.B2(n_340),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_3232),
.B(n_340),
.Y(n_3432)
);

AOI211xp5_ASAP7_75t_L g3433 ( 
.A1(n_3233),
.A2(n_3184),
.B(n_3231),
.C(n_3198),
.Y(n_3433)
);

OAI221xp5_ASAP7_75t_L g3434 ( 
.A1(n_3226),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.C(n_345),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3283),
.B(n_344),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3289),
.Y(n_3436)
);

NAND2x1p5_ASAP7_75t_L g3437 ( 
.A(n_3294),
.B(n_345),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3309),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_SL g3439 ( 
.A(n_3234),
.B(n_346),
.Y(n_3439)
);

OAI22xp33_ASAP7_75t_L g3440 ( 
.A1(n_3248),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_3440)
);

AOI322xp5_ASAP7_75t_L g3441 ( 
.A1(n_3211),
.A2(n_3214),
.A3(n_3225),
.B1(n_3223),
.B2(n_3221),
.C1(n_3310),
.C2(n_350),
.Y(n_3441)
);

AOI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3269),
.A2(n_350),
.B1(n_347),
.B2(n_349),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3169),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_3270),
.B(n_351),
.Y(n_3444)
);

AOI211xp5_ASAP7_75t_L g3445 ( 
.A1(n_3393),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_3445)
);

NOR4xp25_ASAP7_75t_SL g3446 ( 
.A(n_3406),
.B(n_355),
.C(n_353),
.D(n_354),
.Y(n_3446)
);

INVx1_ASAP7_75t_L g3447 ( 
.A(n_3366),
.Y(n_3447)
);

OAI322xp33_ASAP7_75t_L g3448 ( 
.A1(n_3363),
.A2(n_360),
.A3(n_359),
.B1(n_357),
.B2(n_355),
.C1(n_356),
.C2(n_358),
.Y(n_3448)
);

AND2x2_ASAP7_75t_L g3449 ( 
.A(n_3324),
.B(n_357),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3337),
.A2(n_358),
.B(n_359),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3332),
.B(n_360),
.Y(n_3451)
);

HB1xp67_ASAP7_75t_L g3452 ( 
.A(n_3333),
.Y(n_3452)
);

O2A1O1Ixp33_ASAP7_75t_L g3453 ( 
.A1(n_3358),
.A2(n_364),
.B(n_362),
.C(n_363),
.Y(n_3453)
);

AOI22xp33_ASAP7_75t_SL g3454 ( 
.A1(n_3334),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3387),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3321),
.Y(n_3456)
);

OAI31xp33_ASAP7_75t_L g3457 ( 
.A1(n_3365),
.A2(n_368),
.A3(n_365),
.B(n_367),
.Y(n_3457)
);

NOR2x1p5_ASAP7_75t_L g3458 ( 
.A(n_3327),
.B(n_3341),
.Y(n_3458)
);

OAI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3362),
.A2(n_365),
.B(n_367),
.Y(n_3459)
);

A2O1A1Ixp33_ASAP7_75t_L g3460 ( 
.A1(n_3325),
.A2(n_371),
.B(n_368),
.C(n_370),
.Y(n_3460)
);

HB1xp67_ASAP7_75t_L g3461 ( 
.A(n_3437),
.Y(n_3461)
);

OR2x2_ASAP7_75t_L g3462 ( 
.A(n_3384),
.B(n_370),
.Y(n_3462)
);

AOI21xp5_ASAP7_75t_L g3463 ( 
.A1(n_3367),
.A2(n_372),
.B(n_373),
.Y(n_3463)
);

NOR2x1_ASAP7_75t_SL g3464 ( 
.A(n_3354),
.B(n_372),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3359),
.B(n_374),
.Y(n_3465)
);

NAND3xp33_ASAP7_75t_SL g3466 ( 
.A(n_3331),
.B(n_376),
.C(n_379),
.Y(n_3466)
);

AOI22xp33_ASAP7_75t_L g3467 ( 
.A1(n_3395),
.A2(n_3342),
.B1(n_3351),
.B2(n_3374),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3443),
.Y(n_3468)
);

NAND4xp75_ASAP7_75t_SL g3469 ( 
.A(n_3389),
.B(n_381),
.C(n_379),
.D(n_380),
.Y(n_3469)
);

INVx1_ASAP7_75t_SL g3470 ( 
.A(n_3404),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3319),
.Y(n_3471)
);

AOI32xp33_ASAP7_75t_L g3472 ( 
.A1(n_3433),
.A2(n_383),
.A3(n_380),
.B1(n_382),
.B2(n_384),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3360),
.B(n_3347),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3355),
.B(n_382),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3444),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3427),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3343),
.B(n_383),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_3375),
.Y(n_3478)
);

AOI22xp5_ASAP7_75t_L g3479 ( 
.A1(n_3378),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_3479)
);

INVx2_ASAP7_75t_SL g3480 ( 
.A(n_3335),
.Y(n_3480)
);

OAI332xp33_ASAP7_75t_L g3481 ( 
.A1(n_3339),
.A2(n_385),
.A3(n_388),
.B1(n_389),
.B2(n_390),
.B3(n_391),
.C1(n_392),
.C2(n_395),
.Y(n_3481)
);

OR2x2_ASAP7_75t_L g3482 ( 
.A(n_3352),
.B(n_389),
.Y(n_3482)
);

OAI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_3320),
.A2(n_391),
.B(n_392),
.Y(n_3483)
);

AND2x4_ASAP7_75t_L g3484 ( 
.A(n_3425),
.B(n_3397),
.Y(n_3484)
);

OAI22xp33_ASAP7_75t_L g3485 ( 
.A1(n_3325),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3323),
.Y(n_3486)
);

OR2x2_ASAP7_75t_L g3487 ( 
.A(n_3356),
.B(n_396),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3397),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3390),
.Y(n_3489)
);

INVx1_ASAP7_75t_L g3490 ( 
.A(n_3369),
.Y(n_3490)
);

OAI22xp33_ASAP7_75t_L g3491 ( 
.A1(n_3442),
.A2(n_401),
.B1(n_399),
.B2(n_400),
.Y(n_3491)
);

INVxp67_ASAP7_75t_L g3492 ( 
.A(n_3432),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3346),
.Y(n_3493)
);

XOR2x2_ASAP7_75t_L g3494 ( 
.A(n_3400),
.B(n_399),
.Y(n_3494)
);

NAND3xp33_ASAP7_75t_SL g3495 ( 
.A(n_3318),
.B(n_400),
.C(n_401),
.Y(n_3495)
);

NOR2xp33_ASAP7_75t_L g3496 ( 
.A(n_3368),
.B(n_3326),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3379),
.B(n_402),
.Y(n_3497)
);

A2O1A1Ixp33_ASAP7_75t_L g3498 ( 
.A1(n_3442),
.A2(n_404),
.B(n_402),
.C(n_403),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3409),
.Y(n_3499)
);

INVx1_ASAP7_75t_SL g3500 ( 
.A(n_3370),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3372),
.B(n_403),
.Y(n_3501)
);

OAI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3338),
.A2(n_407),
.B1(n_404),
.B2(n_405),
.Y(n_3502)
);

OR2x2_ASAP7_75t_L g3503 ( 
.A(n_3411),
.B(n_405),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3396),
.Y(n_3504)
);

OAI221xp5_ASAP7_75t_L g3505 ( 
.A1(n_3322),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.C(n_411),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3428),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3435),
.Y(n_3507)
);

AOI221xp5_ASAP7_75t_L g3508 ( 
.A1(n_3407),
.A2(n_412),
.B1(n_409),
.B2(n_410),
.C(n_413),
.Y(n_3508)
);

INVxp67_ASAP7_75t_L g3509 ( 
.A(n_3350),
.Y(n_3509)
);

OAI322xp33_ASAP7_75t_L g3510 ( 
.A1(n_3419),
.A2(n_413),
.A3(n_414),
.B1(n_415),
.B2(n_416),
.C1(n_418),
.C2(n_419),
.Y(n_3510)
);

INVx2_ASAP7_75t_SL g3511 ( 
.A(n_3420),
.Y(n_3511)
);

OAI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3349),
.A2(n_3371),
.B(n_3392),
.Y(n_3512)
);

NAND2xp33_ASAP7_75t_L g3513 ( 
.A(n_3391),
.B(n_414),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3348),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3353),
.B(n_3373),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3345),
.Y(n_3516)
);

HB1xp67_ASAP7_75t_L g3517 ( 
.A(n_3422),
.Y(n_3517)
);

OAI33xp33_ASAP7_75t_L g3518 ( 
.A1(n_3424),
.A2(n_420),
.A3(n_422),
.B1(n_416),
.B2(n_419),
.B3(n_421),
.Y(n_3518)
);

OAI32xp33_ASAP7_75t_L g3519 ( 
.A1(n_3412),
.A2(n_424),
.A3(n_420),
.B1(n_423),
.B2(n_425),
.Y(n_3519)
);

INVx1_ASAP7_75t_SL g3520 ( 
.A(n_3414),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3403),
.B(n_3416),
.Y(n_3521)
);

OAI21xp5_ASAP7_75t_L g3522 ( 
.A1(n_3441),
.A2(n_425),
.B(n_427),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3381),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3382),
.Y(n_3524)
);

OAI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_3439),
.A2(n_427),
.B(n_428),
.Y(n_3525)
);

AO21x1_ASAP7_75t_L g3526 ( 
.A1(n_3421),
.A2(n_428),
.B(n_429),
.Y(n_3526)
);

CKINVDCx16_ASAP7_75t_R g3527 ( 
.A(n_3401),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3436),
.Y(n_3528)
);

OAI21xp5_ASAP7_75t_SL g3529 ( 
.A1(n_3408),
.A2(n_431),
.B(n_433),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_L g3530 ( 
.A(n_3336),
.B(n_433),
.Y(n_3530)
);

OAI22xp5_ASAP7_75t_L g3531 ( 
.A1(n_3330),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_3531)
);

AND2x4_ASAP7_75t_L g3532 ( 
.A(n_3438),
.B(n_434),
.Y(n_3532)
);

INVx2_ASAP7_75t_SL g3533 ( 
.A(n_3377),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_SL g3534 ( 
.A1(n_3430),
.A2(n_436),
.B(n_437),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3380),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3383),
.B(n_437),
.Y(n_3536)
);

O2A1O1Ixp33_ASAP7_75t_L g3537 ( 
.A1(n_3344),
.A2(n_441),
.B(n_438),
.C(n_439),
.Y(n_3537)
);

NOR3xp33_ASAP7_75t_L g3538 ( 
.A(n_3434),
.B(n_3340),
.C(n_3426),
.Y(n_3538)
);

AOI22xp33_ASAP7_75t_SL g3539 ( 
.A1(n_3328),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3385),
.Y(n_3540)
);

AOI211xp5_ASAP7_75t_L g3541 ( 
.A1(n_3361),
.A2(n_446),
.B(n_442),
.C(n_443),
.Y(n_3541)
);

OR2x2_ASAP7_75t_L g3542 ( 
.A(n_3417),
.B(n_3399),
.Y(n_3542)
);

NOR2xp33_ASAP7_75t_L g3543 ( 
.A(n_3413),
.B(n_447),
.Y(n_3543)
);

AOI321xp33_ASAP7_75t_L g3544 ( 
.A1(n_3388),
.A2(n_449),
.A3(n_452),
.B1(n_447),
.B2(n_448),
.C(n_450),
.Y(n_3544)
);

NAND2x1_ASAP7_75t_L g3545 ( 
.A(n_3410),
.B(n_3418),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3402),
.B(n_449),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3329),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3386),
.Y(n_3548)
);

AOI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3376),
.A2(n_453),
.B1(n_450),
.B2(n_452),
.Y(n_3549)
);

INVxp67_ASAP7_75t_L g3550 ( 
.A(n_3415),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3394),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3429),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3405),
.Y(n_3553)
);

OAI22xp33_ASAP7_75t_L g3554 ( 
.A1(n_3398),
.A2(n_455),
.B1(n_453),
.B2(n_454),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3440),
.B(n_454),
.Y(n_3555)
);

OAI21xp33_ASAP7_75t_L g3556 ( 
.A1(n_3357),
.A2(n_3364),
.B(n_3431),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3423),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3366),
.Y(n_3558)
);

NAND3xp33_ASAP7_75t_L g3559 ( 
.A(n_3337),
.B(n_457),
.C(n_458),
.Y(n_3559)
);

OAI31xp33_ASAP7_75t_L g3560 ( 
.A1(n_3337),
.A2(n_463),
.A3(n_459),
.B(n_461),
.Y(n_3560)
);

OR2x2_ASAP7_75t_L g3561 ( 
.A(n_3393),
.B(n_459),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3324),
.B(n_461),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_3332),
.Y(n_3563)
);

OR2x2_ASAP7_75t_L g3564 ( 
.A(n_3393),
.B(n_463),
.Y(n_3564)
);

INVx1_ASAP7_75t_SL g3565 ( 
.A(n_3324),
.Y(n_3565)
);

INVx1_ASAP7_75t_SL g3566 ( 
.A(n_3324),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3324),
.B(n_464),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_3327),
.A2(n_466),
.B1(n_464),
.B2(n_465),
.Y(n_3568)
);

AOI21xp5_ASAP7_75t_L g3569 ( 
.A1(n_3406),
.A2(n_467),
.B(n_468),
.Y(n_3569)
);

OAI221xp5_ASAP7_75t_L g3570 ( 
.A1(n_3393),
.A2(n_470),
.B1(n_467),
.B2(n_469),
.C(n_471),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3324),
.B(n_469),
.Y(n_3571)
);

OR2x2_ASAP7_75t_L g3572 ( 
.A(n_3393),
.B(n_471),
.Y(n_3572)
);

NOR2xp33_ASAP7_75t_L g3573 ( 
.A(n_3324),
.B(n_472),
.Y(n_3573)
);

NAND3xp33_ASAP7_75t_L g3574 ( 
.A(n_3337),
.B(n_472),
.C(n_473),
.Y(n_3574)
);

INVxp67_ASAP7_75t_L g3575 ( 
.A(n_3366),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3332),
.Y(n_3576)
);

NOR2xp67_ASAP7_75t_SL g3577 ( 
.A(n_3327),
.B(n_473),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3366),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3324),
.B(n_474),
.Y(n_3579)
);

INVx1_ASAP7_75t_L g3580 ( 
.A(n_3366),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3324),
.B(n_474),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3366),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3366),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3324),
.B(n_475),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3366),
.Y(n_3585)
);

AOI32xp33_ASAP7_75t_L g3586 ( 
.A1(n_3393),
.A2(n_478),
.A3(n_476),
.B1(n_477),
.B2(n_479),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3406),
.A2(n_478),
.B(n_479),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3324),
.B(n_480),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_L g3589 ( 
.A(n_3324),
.B(n_480),
.Y(n_3589)
);

INVx1_ASAP7_75t_SL g3590 ( 
.A(n_3324),
.Y(n_3590)
);

OAI211xp5_ASAP7_75t_L g3591 ( 
.A1(n_3406),
.A2(n_483),
.B(n_481),
.C(n_482),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3324),
.B(n_481),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3324),
.B(n_483),
.Y(n_3593)
);

INVx1_ASAP7_75t_L g3594 ( 
.A(n_3366),
.Y(n_3594)
);

OAI21xp33_ASAP7_75t_L g3595 ( 
.A1(n_3324),
.A2(n_484),
.B(n_486),
.Y(n_3595)
);

INVx2_ASAP7_75t_L g3596 ( 
.A(n_3332),
.Y(n_3596)
);

INVxp67_ASAP7_75t_L g3597 ( 
.A(n_3366),
.Y(n_3597)
);

INVx2_ASAP7_75t_L g3598 ( 
.A(n_3332),
.Y(n_3598)
);

AOI22xp5_ASAP7_75t_L g3599 ( 
.A1(n_3324),
.A2(n_487),
.B1(n_484),
.B2(n_486),
.Y(n_3599)
);

NAND2x1_ASAP7_75t_SL g3600 ( 
.A(n_3333),
.B(n_487),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3324),
.B(n_488),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3366),
.Y(n_3602)
);

INVx2_ASAP7_75t_SL g3603 ( 
.A(n_3600),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3563),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3565),
.B(n_489),
.Y(n_3605)
);

OAI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3450),
.A2(n_3597),
.B(n_3575),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3566),
.B(n_491),
.Y(n_3607)
);

NOR2x1_ASAP7_75t_L g3608 ( 
.A(n_3559),
.B(n_492),
.Y(n_3608)
);

OAI322xp33_ASAP7_75t_L g3609 ( 
.A1(n_3496),
.A2(n_493),
.A3(n_494),
.B1(n_495),
.B2(n_496),
.C1(n_497),
.C2(n_498),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3452),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_3513),
.A2(n_493),
.B(n_496),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3484),
.B(n_497),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_SL g3613 ( 
.A(n_3484),
.B(n_498),
.Y(n_3613)
);

O2A1O1Ixp33_ASAP7_75t_SL g3614 ( 
.A1(n_3478),
.A2(n_501),
.B(n_499),
.C(n_500),
.Y(n_3614)
);

HB1xp67_ASAP7_75t_L g3615 ( 
.A(n_3461),
.Y(n_3615)
);

AOI221xp5_ASAP7_75t_L g3616 ( 
.A1(n_3448),
.A2(n_3522),
.B1(n_3495),
.B2(n_3466),
.C(n_3554),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3464),
.Y(n_3617)
);

AOI211x1_ASAP7_75t_L g3618 ( 
.A1(n_3526),
.A2(n_502),
.B(n_500),
.C(n_501),
.Y(n_3618)
);

NAND2xp5_ASAP7_75t_L g3619 ( 
.A(n_3590),
.B(n_503),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3576),
.B(n_503),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3561),
.Y(n_3621)
);

NOR2xp33_ASAP7_75t_L g3622 ( 
.A(n_3596),
.B(n_504),
.Y(n_3622)
);

NOR3xp33_ASAP7_75t_L g3623 ( 
.A(n_3527),
.B(n_504),
.C(n_505),
.Y(n_3623)
);

OAI21xp5_ASAP7_75t_SL g3624 ( 
.A1(n_3529),
.A2(n_505),
.B(n_507),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_3537),
.B(n_3560),
.Y(n_3625)
);

INVx1_ASAP7_75t_L g3626 ( 
.A(n_3564),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3598),
.B(n_508),
.Y(n_3627)
);

CKINVDCx20_ASAP7_75t_R g3628 ( 
.A(n_3494),
.Y(n_3628)
);

NOR2xp33_ASAP7_75t_L g3629 ( 
.A(n_3470),
.B(n_508),
.Y(n_3629)
);

AOI211xp5_ASAP7_75t_L g3630 ( 
.A1(n_3570),
.A2(n_512),
.B(n_509),
.C(n_510),
.Y(n_3630)
);

NOR3xp33_ASAP7_75t_L g3631 ( 
.A(n_3492),
.B(n_509),
.C(n_512),
.Y(n_3631)
);

AOI211xp5_ASAP7_75t_L g3632 ( 
.A1(n_3556),
.A2(n_515),
.B(n_513),
.C(n_514),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3447),
.B(n_514),
.Y(n_3633)
);

OAI211xp5_ASAP7_75t_SL g3634 ( 
.A1(n_3467),
.A2(n_521),
.B(n_516),
.C(n_519),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3558),
.B(n_516),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_SL g3636 ( 
.A(n_3586),
.B(n_519),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3449),
.B(n_522),
.Y(n_3637)
);

AOI22xp5_ASAP7_75t_L g3638 ( 
.A1(n_3551),
.A2(n_526),
.B1(n_523),
.B2(n_525),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_3578),
.B(n_525),
.Y(n_3639)
);

NAND4xp25_ASAP7_75t_SL g3640 ( 
.A(n_3472),
.B(n_529),
.C(n_527),
.D(n_528),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3572),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3567),
.Y(n_3642)
);

NAND4xp25_ASAP7_75t_L g3643 ( 
.A(n_3538),
.B(n_530),
.C(n_527),
.D(n_529),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3580),
.B(n_530),
.Y(n_3644)
);

AOI211xp5_ASAP7_75t_L g3645 ( 
.A1(n_3582),
.A2(n_534),
.B(n_532),
.C(n_533),
.Y(n_3645)
);

OR2x2_ASAP7_75t_L g3646 ( 
.A(n_3473),
.B(n_532),
.Y(n_3646)
);

NOR3xp33_ASAP7_75t_SL g3647 ( 
.A(n_3583),
.B(n_534),
.C(n_535),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_SL g3648 ( 
.A(n_3539),
.B(n_535),
.Y(n_3648)
);

NOR2xp67_ASAP7_75t_L g3649 ( 
.A(n_3574),
.B(n_538),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_L g3650 ( 
.A(n_3585),
.B(n_538),
.Y(n_3650)
);

HB1xp67_ASAP7_75t_L g3651 ( 
.A(n_3469),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3594),
.B(n_539),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_L g3653 ( 
.A(n_3602),
.B(n_3480),
.Y(n_3653)
);

NOR2xp33_ASAP7_75t_L g3654 ( 
.A(n_3499),
.B(n_541),
.Y(n_3654)
);

INVxp67_ASAP7_75t_SL g3655 ( 
.A(n_3577),
.Y(n_3655)
);

NOR3xp33_ASAP7_75t_L g3656 ( 
.A(n_3455),
.B(n_541),
.C(n_542),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3571),
.B(n_543),
.Y(n_3657)
);

INVxp67_ASAP7_75t_L g3658 ( 
.A(n_3573),
.Y(n_3658)
);

NAND2xp33_ASAP7_75t_L g3659 ( 
.A(n_3476),
.B(n_543),
.Y(n_3659)
);

NAND2xp5_ASAP7_75t_L g3660 ( 
.A(n_3497),
.B(n_544),
.Y(n_3660)
);

AOI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_3463),
.A2(n_545),
.B(n_546),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3454),
.B(n_545),
.Y(n_3662)
);

NOR3xp33_ASAP7_75t_L g3663 ( 
.A(n_3557),
.B(n_546),
.C(n_547),
.Y(n_3663)
);

NOR3x1_ASAP7_75t_L g3664 ( 
.A(n_3534),
.B(n_547),
.C(n_548),
.Y(n_3664)
);

NOR2xp67_ASAP7_75t_L g3665 ( 
.A(n_3488),
.B(n_548),
.Y(n_3665)
);

AOI31xp33_ASAP7_75t_L g3666 ( 
.A1(n_3541),
.A2(n_551),
.A3(n_549),
.B(n_550),
.Y(n_3666)
);

OAI21xp5_ASAP7_75t_L g3667 ( 
.A1(n_3569),
.A2(n_549),
.B(n_550),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3445),
.B(n_551),
.Y(n_3668)
);

AOI211xp5_ASAP7_75t_L g3669 ( 
.A1(n_3587),
.A2(n_555),
.B(n_552),
.C(n_553),
.Y(n_3669)
);

NOR3x1_ASAP7_75t_L g3670 ( 
.A(n_3591),
.B(n_3483),
.C(n_3512),
.Y(n_3670)
);

XOR2x2_ASAP7_75t_L g3671 ( 
.A(n_3474),
.B(n_552),
.Y(n_3671)
);

NAND2x1p5_ASAP7_75t_L g3672 ( 
.A(n_3545),
.B(n_3458),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_3595),
.B(n_553),
.Y(n_3673)
);

OAI22xp5_ASAP7_75t_L g3674 ( 
.A1(n_3462),
.A2(n_3479),
.B1(n_3549),
.B2(n_3546),
.Y(n_3674)
);

NAND3xp33_ASAP7_75t_L g3675 ( 
.A(n_3457),
.B(n_555),
.C(n_556),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3519),
.B(n_556),
.Y(n_3676)
);

O2A1O1Ixp33_ASAP7_75t_SL g3677 ( 
.A1(n_3460),
.A2(n_560),
.B(n_558),
.C(n_559),
.Y(n_3677)
);

OAI21xp33_ASAP7_75t_L g3678 ( 
.A1(n_3553),
.A2(n_558),
.B(n_560),
.Y(n_3678)
);

NOR2x1_ASAP7_75t_SL g3679 ( 
.A(n_3511),
.B(n_562),
.Y(n_3679)
);

NOR2xp33_ASAP7_75t_SL g3680 ( 
.A(n_3504),
.B(n_562),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3451),
.Y(n_3681)
);

OAI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3456),
.A2(n_564),
.B(n_565),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3562),
.B(n_564),
.Y(n_3683)
);

NOR3xp33_ASAP7_75t_SL g3684 ( 
.A(n_3547),
.B(n_565),
.C(n_568),
.Y(n_3684)
);

OAI211xp5_ASAP7_75t_SL g3685 ( 
.A1(n_3550),
.A2(n_571),
.B(n_568),
.C(n_570),
.Y(n_3685)
);

OAI21xp5_ASAP7_75t_L g3686 ( 
.A1(n_3468),
.A2(n_570),
.B(n_571),
.Y(n_3686)
);

OAI211xp5_ASAP7_75t_L g3687 ( 
.A1(n_3446),
.A2(n_575),
.B(n_572),
.C(n_574),
.Y(n_3687)
);

AOI221xp5_ASAP7_75t_L g3688 ( 
.A1(n_3485),
.A2(n_3491),
.B1(n_3535),
.B2(n_3517),
.C(n_3520),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3453),
.A2(n_572),
.B(n_576),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3544),
.B(n_577),
.Y(n_3690)
);

NOR3x1_ASAP7_75t_L g3691 ( 
.A(n_3505),
.B(n_578),
.C(n_579),
.Y(n_3691)
);

NOR2x1_ASAP7_75t_L g3692 ( 
.A(n_3510),
.B(n_578),
.Y(n_3692)
);

HB1xp67_ASAP7_75t_L g3693 ( 
.A(n_3532),
.Y(n_3693)
);

OAI21xp5_ASAP7_75t_L g3694 ( 
.A1(n_3498),
.A2(n_580),
.B(n_581),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_3579),
.B(n_581),
.Y(n_3695)
);

A2O1A1Ixp33_ASAP7_75t_L g3696 ( 
.A1(n_3603),
.A2(n_3653),
.B(n_3665),
.C(n_3617),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3655),
.A2(n_3584),
.B(n_3581),
.Y(n_3697)
);

OAI211xp5_ASAP7_75t_SL g3698 ( 
.A1(n_3688),
.A2(n_3509),
.B(n_3500),
.C(n_3471),
.Y(n_3698)
);

OA22x2_ASAP7_75t_L g3699 ( 
.A1(n_3624),
.A2(n_3533),
.B1(n_3493),
.B2(n_3475),
.Y(n_3699)
);

AOI32xp33_ASAP7_75t_L g3700 ( 
.A1(n_3634),
.A2(n_3521),
.A3(n_3515),
.B1(n_3552),
.B2(n_3548),
.Y(n_3700)
);

NOR3x1_ASAP7_75t_L g3701 ( 
.A(n_3687),
.B(n_3525),
.C(n_3588),
.Y(n_3701)
);

NOR2x1_ASAP7_75t_L g3702 ( 
.A(n_3628),
.B(n_3643),
.Y(n_3702)
);

NAND3xp33_ASAP7_75t_L g3703 ( 
.A(n_3618),
.B(n_3540),
.C(n_3528),
.Y(n_3703)
);

OAI22xp33_ASAP7_75t_L g3704 ( 
.A1(n_3672),
.A2(n_3589),
.B1(n_3593),
.B2(n_3592),
.Y(n_3704)
);

NOR3xp33_ASAP7_75t_L g3705 ( 
.A(n_3606),
.B(n_3489),
.C(n_3490),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3693),
.B(n_3477),
.Y(n_3706)
);

OAI21xp33_ASAP7_75t_L g3707 ( 
.A1(n_3604),
.A2(n_3516),
.B(n_3486),
.Y(n_3707)
);

OAI221xp5_ASAP7_75t_L g3708 ( 
.A1(n_3672),
.A2(n_3616),
.B1(n_3678),
.B2(n_3610),
.C(n_3615),
.Y(n_3708)
);

OAI221xp5_ASAP7_75t_L g3709 ( 
.A1(n_3667),
.A2(n_3514),
.B1(n_3508),
.B2(n_3601),
.C(n_3465),
.Y(n_3709)
);

NAND4xp25_ASAP7_75t_L g3710 ( 
.A(n_3670),
.B(n_3542),
.C(n_3506),
.D(n_3524),
.Y(n_3710)
);

AOI22xp5_ASAP7_75t_L g3711 ( 
.A1(n_3690),
.A2(n_3531),
.B1(n_3502),
.B2(n_3543),
.Y(n_3711)
);

AOI22xp33_ASAP7_75t_SL g3712 ( 
.A1(n_3679),
.A2(n_3523),
.B1(n_3507),
.B2(n_3555),
.Y(n_3712)
);

NOR2xp33_ASAP7_75t_R g3713 ( 
.A(n_3640),
.B(n_3659),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_3637),
.B(n_3532),
.Y(n_3714)
);

AOI221xp5_ASAP7_75t_L g3715 ( 
.A1(n_3666),
.A2(n_3518),
.B1(n_3481),
.B2(n_3459),
.C(n_3501),
.Y(n_3715)
);

OAI211xp5_ASAP7_75t_L g3716 ( 
.A1(n_3651),
.A2(n_3599),
.B(n_3568),
.C(n_3503),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3642),
.B(n_3536),
.Y(n_3717)
);

AOI211xp5_ASAP7_75t_SL g3718 ( 
.A1(n_3674),
.A2(n_3530),
.B(n_3487),
.C(n_3482),
.Y(n_3718)
);

NOR3x1_ASAP7_75t_L g3719 ( 
.A(n_3675),
.B(n_3536),
.C(n_582),
.Y(n_3719)
);

AOI211xp5_ASAP7_75t_L g3720 ( 
.A1(n_3614),
.A2(n_3609),
.B(n_3677),
.C(n_3685),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_SL g3721 ( 
.A(n_3680),
.B(n_582),
.Y(n_3721)
);

OAI21xp5_ASAP7_75t_L g3722 ( 
.A1(n_3692),
.A2(n_583),
.B(n_584),
.Y(n_3722)
);

OAI21xp33_ASAP7_75t_L g3723 ( 
.A1(n_3625),
.A2(n_583),
.B(n_585),
.Y(n_3723)
);

OAI21xp5_ASAP7_75t_SL g3724 ( 
.A1(n_3638),
.A2(n_585),
.B(n_586),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3605),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3664),
.B(n_586),
.Y(n_3726)
);

NOR3x1_ASAP7_75t_L g3727 ( 
.A(n_3694),
.B(n_587),
.C(n_588),
.Y(n_3727)
);

AOI311xp33_ASAP7_75t_L g3728 ( 
.A1(n_3621),
.A2(n_588),
.A3(n_589),
.B(n_590),
.C(n_591),
.Y(n_3728)
);

NAND3xp33_ASAP7_75t_SL g3729 ( 
.A(n_3630),
.B(n_590),
.C(n_591),
.Y(n_3729)
);

AOI21xp33_ASAP7_75t_L g3730 ( 
.A1(n_3646),
.A2(n_594),
.B(n_595),
.Y(n_3730)
);

NOR3xp33_ASAP7_75t_L g3731 ( 
.A(n_3658),
.B(n_596),
.C(n_597),
.Y(n_3731)
);

OAI322xp33_ASAP7_75t_L g3732 ( 
.A1(n_3636),
.A2(n_598),
.A3(n_599),
.B1(n_601),
.B2(n_602),
.C1(n_603),
.C2(n_604),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_L g3733 ( 
.A(n_3612),
.B(n_598),
.Y(n_3733)
);

AOI21xp33_ASAP7_75t_SL g3734 ( 
.A1(n_3613),
.A2(n_599),
.B(n_602),
.Y(n_3734)
);

AND2x2_ASAP7_75t_L g3735 ( 
.A(n_3626),
.B(n_603),
.Y(n_3735)
);

INVxp67_ASAP7_75t_L g3736 ( 
.A(n_3629),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3676),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_3737)
);

OAI21xp33_ASAP7_75t_L g3738 ( 
.A1(n_3671),
.A2(n_605),
.B(n_607),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3683),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3607),
.Y(n_3740)
);

OAI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3689),
.A2(n_607),
.B(n_608),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3641),
.B(n_609),
.Y(n_3742)
);

NAND3xp33_ASAP7_75t_L g3743 ( 
.A(n_3632),
.B(n_610),
.C(n_611),
.Y(n_3743)
);

NAND3xp33_ASAP7_75t_L g3744 ( 
.A(n_3684),
.B(n_610),
.C(n_611),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3660),
.Y(n_3745)
);

O2A1O1Ixp5_ASAP7_75t_L g3746 ( 
.A1(n_3648),
.A2(n_614),
.B(n_612),
.C(n_613),
.Y(n_3746)
);

AOI221xp5_ASAP7_75t_L g3747 ( 
.A1(n_3681),
.A2(n_613),
.B1(n_617),
.B2(n_618),
.C(n_619),
.Y(n_3747)
);

OAI211xp5_ASAP7_75t_L g3748 ( 
.A1(n_3608),
.A2(n_619),
.B(n_617),
.C(n_618),
.Y(n_3748)
);

AOI222xp33_ASAP7_75t_L g3749 ( 
.A1(n_3649),
.A2(n_620),
.B1(n_621),
.B2(n_622),
.C1(n_623),
.C2(n_624),
.Y(n_3749)
);

NAND3xp33_ASAP7_75t_L g3750 ( 
.A(n_3669),
.B(n_620),
.C(n_622),
.Y(n_3750)
);

INVxp67_ASAP7_75t_SL g3751 ( 
.A(n_3619),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3657),
.Y(n_3752)
);

AOI221xp5_ASAP7_75t_L g3753 ( 
.A1(n_3663),
.A2(n_624),
.B1(n_625),
.B2(n_626),
.C(n_627),
.Y(n_3753)
);

NAND3xp33_ASAP7_75t_L g3754 ( 
.A(n_3647),
.B(n_626),
.C(n_628),
.Y(n_3754)
);

AOI21xp33_ASAP7_75t_L g3755 ( 
.A1(n_3633),
.A2(n_629),
.B(n_630),
.Y(n_3755)
);

O2A1O1Ixp33_ASAP7_75t_L g3756 ( 
.A1(n_3661),
.A2(n_629),
.B(n_632),
.C(n_633),
.Y(n_3756)
);

OAI221xp5_ASAP7_75t_L g3757 ( 
.A1(n_3620),
.A2(n_634),
.B1(n_635),
.B2(n_636),
.C(n_637),
.Y(n_3757)
);

OAI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3737),
.A2(n_3662),
.B1(n_3668),
.B2(n_3627),
.Y(n_3758)
);

OAI221xp5_ASAP7_75t_L g3759 ( 
.A1(n_3696),
.A2(n_3650),
.B1(n_3639),
.B2(n_3652),
.C(n_3635),
.Y(n_3759)
);

HB1xp67_ASAP7_75t_L g3760 ( 
.A(n_3726),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3706),
.Y(n_3761)
);

OAI221xp5_ASAP7_75t_L g3762 ( 
.A1(n_3708),
.A2(n_3644),
.B1(n_3622),
.B2(n_3686),
.C(n_3682),
.Y(n_3762)
);

AOI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3698),
.A2(n_3673),
.B1(n_3623),
.B2(n_3656),
.Y(n_3763)
);

OAI22xp5_ASAP7_75t_L g3764 ( 
.A1(n_3711),
.A2(n_3645),
.B1(n_3695),
.B2(n_3654),
.Y(n_3764)
);

OAI211xp5_ASAP7_75t_L g3765 ( 
.A1(n_3722),
.A2(n_3700),
.B(n_3716),
.C(n_3707),
.Y(n_3765)
);

INVx1_ASAP7_75t_L g3766 ( 
.A(n_3714),
.Y(n_3766)
);

AOI22xp5_ASAP7_75t_L g3767 ( 
.A1(n_3702),
.A2(n_3631),
.B1(n_3611),
.B2(n_3691),
.Y(n_3767)
);

HB1xp67_ASAP7_75t_L g3768 ( 
.A(n_3713),
.Y(n_3768)
);

INVx2_ASAP7_75t_L g3769 ( 
.A(n_3735),
.Y(n_3769)
);

OAI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_3754),
.A2(n_634),
.B1(n_637),
.B2(n_638),
.Y(n_3770)
);

INVx2_ASAP7_75t_SL g3771 ( 
.A(n_3742),
.Y(n_3771)
);

AOI22xp5_ASAP7_75t_L g3772 ( 
.A1(n_3705),
.A2(n_639),
.B1(n_640),
.B2(n_641),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3717),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3699),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3703),
.Y(n_3775)
);

HB1xp67_ASAP7_75t_L g3776 ( 
.A(n_3727),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3744),
.Y(n_3777)
);

AOI22xp5_ASAP7_75t_L g3778 ( 
.A1(n_3715),
.A2(n_3738),
.B1(n_3729),
.B2(n_3710),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3739),
.Y(n_3779)
);

A2O1A1Ixp33_ASAP7_75t_L g3780 ( 
.A1(n_3756),
.A2(n_639),
.B(n_640),
.C(n_641),
.Y(n_3780)
);

BUFx2_ASAP7_75t_L g3781 ( 
.A(n_3741),
.Y(n_3781)
);

INVx1_ASAP7_75t_SL g3782 ( 
.A(n_3721),
.Y(n_3782)
);

AOI221xp5_ASAP7_75t_L g3783 ( 
.A1(n_3704),
.A2(n_642),
.B1(n_643),
.B2(n_644),
.C(n_645),
.Y(n_3783)
);

OAI22xp5_ASAP7_75t_L g3784 ( 
.A1(n_3743),
.A2(n_642),
.B1(n_644),
.B2(n_645),
.Y(n_3784)
);

BUFx8_ASAP7_75t_L g3785 ( 
.A(n_3725),
.Y(n_3785)
);

INVx1_ASAP7_75t_L g3786 ( 
.A(n_3733),
.Y(n_3786)
);

OAI22xp5_ASAP7_75t_L g3787 ( 
.A1(n_3712),
.A2(n_3750),
.B1(n_3720),
.B2(n_3736),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3748),
.Y(n_3788)
);

INVxp33_ASAP7_75t_SL g3789 ( 
.A(n_3701),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3732),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3723),
.Y(n_3791)
);

AO22x2_ASAP7_75t_L g3792 ( 
.A1(n_3724),
.A2(n_649),
.B1(n_650),
.B2(n_651),
.Y(n_3792)
);

OAI221xp5_ASAP7_75t_SL g3793 ( 
.A1(n_3720),
.A2(n_649),
.B1(n_650),
.B2(n_651),
.C(n_652),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3709),
.A2(n_652),
.B1(n_653),
.B2(n_654),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3746),
.Y(n_3795)
);

A2O1A1Ixp33_ASAP7_75t_L g3796 ( 
.A1(n_3775),
.A2(n_3734),
.B(n_3697),
.C(n_3718),
.Y(n_3796)
);

AOI222xp33_ASAP7_75t_L g3797 ( 
.A1(n_3789),
.A2(n_3774),
.B1(n_3765),
.B2(n_3787),
.C1(n_3788),
.C2(n_3795),
.Y(n_3797)
);

NAND3xp33_ASAP7_75t_SL g3798 ( 
.A(n_3767),
.B(n_3749),
.C(n_3753),
.Y(n_3798)
);

AOI22xp5_ASAP7_75t_L g3799 ( 
.A1(n_3773),
.A2(n_3751),
.B1(n_3740),
.B2(n_3745),
.Y(n_3799)
);

AOI221xp5_ASAP7_75t_L g3800 ( 
.A1(n_3762),
.A2(n_3752),
.B1(n_3730),
.B2(n_3755),
.C(n_3757),
.Y(n_3800)
);

A2O1A1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_3783),
.A2(n_3731),
.B(n_3747),
.C(n_3728),
.Y(n_3801)
);

OAI222xp33_ASAP7_75t_L g3802 ( 
.A1(n_3763),
.A2(n_3719),
.B1(n_655),
.B2(n_656),
.C1(n_657),
.C2(n_658),
.Y(n_3802)
);

OAI211xp5_ASAP7_75t_L g3803 ( 
.A1(n_3778),
.A2(n_3768),
.B(n_3776),
.C(n_3760),
.Y(n_3803)
);

AOI221xp5_ASAP7_75t_L g3804 ( 
.A1(n_3764),
.A2(n_654),
.B1(n_655),
.B2(n_656),
.C(n_658),
.Y(n_3804)
);

INVx1_ASAP7_75t_L g3805 ( 
.A(n_3792),
.Y(n_3805)
);

AOI221xp5_ASAP7_75t_L g3806 ( 
.A1(n_3759),
.A2(n_659),
.B1(n_660),
.B2(n_661),
.C(n_662),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3794),
.A2(n_660),
.B(n_661),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3771),
.B(n_662),
.Y(n_3808)
);

INVx1_ASAP7_75t_L g3809 ( 
.A(n_3792),
.Y(n_3809)
);

OAI22xp5_ASAP7_75t_L g3810 ( 
.A1(n_3793),
.A2(n_663),
.B1(n_664),
.B2(n_665),
.Y(n_3810)
);

INVx1_ASAP7_75t_L g3811 ( 
.A(n_3769),
.Y(n_3811)
);

NOR2x1_ASAP7_75t_L g3812 ( 
.A(n_3779),
.B(n_663),
.Y(n_3812)
);

CKINVDCx5p33_ASAP7_75t_R g3813 ( 
.A(n_3785),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_R g3814 ( 
.A(n_3777),
.B(n_3785),
.Y(n_3814)
);

BUFx2_ASAP7_75t_L g3815 ( 
.A(n_3812),
.Y(n_3815)
);

OAI221xp5_ASAP7_75t_L g3816 ( 
.A1(n_3796),
.A2(n_3780),
.B1(n_3782),
.B2(n_3790),
.C(n_3791),
.Y(n_3816)
);

AOI21xp5_ASAP7_75t_L g3817 ( 
.A1(n_3803),
.A2(n_3770),
.B(n_3758),
.Y(n_3817)
);

AO22x2_ASAP7_75t_L g3818 ( 
.A1(n_3805),
.A2(n_3766),
.B1(n_3761),
.B2(n_3786),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3813),
.B(n_3772),
.Y(n_3819)
);

AOI222xp33_ASAP7_75t_L g3820 ( 
.A1(n_3798),
.A2(n_3781),
.B1(n_3784),
.B2(n_667),
.C1(n_668),
.C2(n_670),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3809),
.Y(n_3821)
);

OAI211xp5_ASAP7_75t_SL g3822 ( 
.A1(n_3797),
.A2(n_3800),
.B(n_3799),
.C(n_3811),
.Y(n_3822)
);

NAND4xp75_ASAP7_75t_L g3823 ( 
.A(n_3808),
.B(n_664),
.C(n_666),
.D(n_667),
.Y(n_3823)
);

AOI221xp5_ASAP7_75t_L g3824 ( 
.A1(n_3802),
.A2(n_666),
.B1(n_668),
.B2(n_670),
.C(n_671),
.Y(n_3824)
);

AOI322xp5_ASAP7_75t_L g3825 ( 
.A1(n_3801),
.A2(n_671),
.A3(n_672),
.B1(n_673),
.B2(n_674),
.C1(n_676),
.C2(n_678),
.Y(n_3825)
);

AOI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_3807),
.A2(n_672),
.B(n_674),
.Y(n_3826)
);

AOI222xp33_ASAP7_75t_L g3827 ( 
.A1(n_3810),
.A2(n_676),
.B1(n_678),
.B2(n_679),
.C1(n_680),
.C2(n_681),
.Y(n_3827)
);

XNOR2xp5_ASAP7_75t_L g3828 ( 
.A(n_3823),
.B(n_3816),
.Y(n_3828)
);

OAI32xp33_ASAP7_75t_L g3829 ( 
.A1(n_3821),
.A2(n_3814),
.A3(n_3806),
.B1(n_3804),
.B2(n_684),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3815),
.Y(n_3830)
);

OAI211xp5_ASAP7_75t_L g3831 ( 
.A1(n_3824),
.A2(n_681),
.B(n_682),
.C(n_683),
.Y(n_3831)
);

AOI22xp33_ASAP7_75t_SL g3832 ( 
.A1(n_3818),
.A2(n_682),
.B1(n_683),
.B2(n_684),
.Y(n_3832)
);

NOR3xp33_ASAP7_75t_L g3833 ( 
.A(n_3822),
.B(n_3819),
.C(n_3817),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3818),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_SL g3835 ( 
.A(n_3827),
.B(n_685),
.Y(n_3835)
);

NAND3xp33_ASAP7_75t_SL g3836 ( 
.A(n_3820),
.B(n_3826),
.C(n_3825),
.Y(n_3836)
);

AND2x2_ASAP7_75t_L g3837 ( 
.A(n_3818),
.B(n_686),
.Y(n_3837)
);

AND2x2_ASAP7_75t_L g3838 ( 
.A(n_3837),
.B(n_687),
.Y(n_3838)
);

OAI321xp33_ASAP7_75t_L g3839 ( 
.A1(n_3834),
.A2(n_687),
.A3(n_689),
.B1(n_690),
.B2(n_691),
.C(n_692),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3830),
.Y(n_3840)
);

INVxp67_ASAP7_75t_SL g3841 ( 
.A(n_3832),
.Y(n_3841)
);

AND2x4_ASAP7_75t_L g3842 ( 
.A(n_3833),
.B(n_690),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3840),
.A2(n_3828),
.B1(n_3831),
.B2(n_3835),
.Y(n_3843)
);

INVx1_ASAP7_75t_L g3844 ( 
.A(n_3838),
.Y(n_3844)
);

AOI21xp5_ASAP7_75t_L g3845 ( 
.A1(n_3841),
.A2(n_3836),
.B(n_3829),
.Y(n_3845)
);

NAND3xp33_ASAP7_75t_SL g3846 ( 
.A(n_3842),
.B(n_691),
.C(n_692),
.Y(n_3846)
);

XNOR2x2_ASAP7_75t_SL g3847 ( 
.A(n_3844),
.B(n_3839),
.Y(n_3847)
);

INVx1_ASAP7_75t_L g3848 ( 
.A(n_3847),
.Y(n_3848)
);

AOI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3848),
.A2(n_3843),
.B1(n_3846),
.B2(n_3845),
.Y(n_3849)
);

OAI22xp5_ASAP7_75t_SL g3850 ( 
.A1(n_3849),
.A2(n_693),
.B1(n_694),
.B2(n_695),
.Y(n_3850)
);

AOI22xp33_ASAP7_75t_L g3851 ( 
.A1(n_3850),
.A2(n_693),
.B1(n_694),
.B2(n_696),
.Y(n_3851)
);

OAI22xp5_ASAP7_75t_SL g3852 ( 
.A1(n_3851),
.A2(n_696),
.B1(n_697),
.B2(n_698),
.Y(n_3852)
);

OAI21xp5_ASAP7_75t_L g3853 ( 
.A1(n_3852),
.A2(n_700),
.B(n_701),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3853),
.Y(n_3854)
);

INVx1_ASAP7_75t_SL g3855 ( 
.A(n_3854),
.Y(n_3855)
);

AO21x2_ASAP7_75t_L g3856 ( 
.A1(n_3855),
.A2(n_700),
.B(n_701),
.Y(n_3856)
);

AOI221xp5_ASAP7_75t_L g3857 ( 
.A1(n_3856),
.A2(n_702),
.B1(n_703),
.B2(n_704),
.C(n_705),
.Y(n_3857)
);

AOI211xp5_ASAP7_75t_L g3858 ( 
.A1(n_3857),
.A2(n_703),
.B(n_704),
.C(n_705),
.Y(n_3858)
);


endmodule