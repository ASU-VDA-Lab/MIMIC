module fake_jpeg_28140_n_309 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_27),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_51),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_54),
.B1(n_33),
.B2(n_25),
.Y(n_70)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_56),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_23),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_16),
.B1(n_32),
.B2(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_62),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_64),
.Y(n_71)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_84),
.B1(n_86),
.B2(n_68),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_79),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_30),
.B1(n_31),
.B2(n_25),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_19),
.B1(n_31),
.B2(n_25),
.Y(n_101)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_33),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_84),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_83),
.B(n_86),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_34),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.C(n_57),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_42),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_43),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_57),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_102),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_41),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_78),
.B1(n_80),
.B2(n_66),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_19),
.A3(n_31),
.B1(n_44),
.B2(n_41),
.Y(n_103)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_109),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_106),
.B1(n_81),
.B2(n_39),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_71),
.A2(n_39),
.B1(n_66),
.B2(n_59),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_82),
.B(n_75),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_18),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_17),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_90),
.B1(n_39),
.B2(n_85),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_39),
.B1(n_85),
.B2(n_91),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_79),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_121),
.B(n_131),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_81),
.B(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_139),
.B1(n_73),
.B2(n_24),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_107),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_75),
.B(n_2),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_133),
.B(n_135),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_140),
.Y(n_156)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_138),
.B1(n_112),
.B2(n_143),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_118),
.B(n_109),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_76),
.B1(n_49),
.B2(n_60),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_80),
.B1(n_38),
.B2(n_76),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_113),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_143),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_58),
.B1(n_55),
.B2(n_34),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_142),
.A2(n_145),
.B1(n_112),
.B2(n_108),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_115),
.A2(n_34),
.B1(n_27),
.B2(n_22),
.Y(n_145)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_153),
.B1(n_165),
.B2(n_175),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_151),
.B1(n_170),
.B2(n_138),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_124),
.B(n_133),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_150),
.A2(n_164),
.B(n_120),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_95),
.B1(n_111),
.B2(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_152),
.B(n_159),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_100),
.B1(n_99),
.B2(n_118),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_108),
.C(n_107),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_132),
.C(n_127),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_128),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_93),
.B1(n_34),
.B2(n_27),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_126),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_73),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_174),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_73),
.Y(n_173)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_137),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_121),
.B(n_132),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_157),
.B(n_152),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_123),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_197),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_195),
.B1(n_18),
.B2(n_9),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_17),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_185),
.C(n_189),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_127),
.C(n_145),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_169),
.B1(n_148),
.B2(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_202),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_151),
.B(n_140),
.C(n_122),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_147),
.C(n_22),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.C(n_198),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_147),
.C(n_24),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_156),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_193),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_176),
.B1(n_149),
.B2(n_158),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_24),
.C(n_17),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_199),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_165),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_168),
.B1(n_157),
.B2(n_175),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_218),
.B1(n_5),
.B2(n_6),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_221),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_194),
.B1(n_187),
.B2(n_203),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_1),
.B(n_2),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_178),
.B1(n_195),
.B2(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_1),
.Y(n_220)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_220),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_10),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_183),
.B(n_10),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_11),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_9),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_226),
.B(n_228),
.C(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_227),
.B(n_188),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_184),
.B(n_9),
.Y(n_228)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_233),
.B1(n_239),
.B2(n_245),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_232),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_180),
.B1(n_207),
.B2(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_237),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_191),
.C(n_188),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_213),
.C(n_215),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_202),
.B1(n_198),
.B2(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_4),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_214),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_243),
.Y(n_263)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_206),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_246),
.A2(n_223),
.B1(n_211),
.B2(n_222),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_6),
.C(n_8),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_221),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_248),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_213),
.C(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_255),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_241),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_228),
.C(n_210),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_216),
.B(n_218),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_261),
.B(n_5),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_246),
.A2(n_225),
.B1(n_219),
.B2(n_8),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_259),
.Y(n_267)
);

OA21x2_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_235),
.B(n_244),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_244),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_266),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_245),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_229),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_257),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_240),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_262),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_249),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_273),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_259),
.B(n_258),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_8),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_268),
.A2(n_253),
.B1(n_256),
.B2(n_254),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

BUFx12f_ASAP7_75t_SL g279 ( 
.A(n_267),
.Y(n_279)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_279),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_267),
.B(n_275),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_287),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_12),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_13),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_292),
.Y(n_296)
);

AOI221xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_266),
.B1(n_270),
.B2(n_265),
.C(n_15),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_290),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_14),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_14),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_289),
.B1(n_15),
.B2(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_286),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_301),
.C(n_296),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_283),
.B(n_278),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_299),
.A2(n_15),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_277),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_302),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_303),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_304),
.Y(n_309)
);


endmodule