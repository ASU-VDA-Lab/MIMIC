module fake_jpeg_1733_n_695 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_695);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_695;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_554;
wire n_280;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_9),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_63),
.Y(n_147)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_11),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_R g218 ( 
.A(n_65),
.B(n_115),
.Y(n_218)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_67),
.Y(n_217)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_73),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_11),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_80),
.Y(n_135)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_75),
.Y(n_175)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

BUFx4f_ASAP7_75t_SL g215 ( 
.A(n_78),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_54),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_81),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

BUFx16f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_87),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_88),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_90),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

CKINVDCx9p33_ASAP7_75t_R g196 ( 
.A(n_91),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_92),
.B(n_117),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_23),
.B(n_11),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_94),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_23),
.B(n_10),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

BUFx16f_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_98),
.B(n_109),
.Y(n_151)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_108),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_41),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_38),
.Y(n_110)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_110),
.Y(n_188)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_35),
.Y(n_111)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_41),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_112),
.B(n_120),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_36),
.B(n_10),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_12),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_118),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_12),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_119),
.B(n_122),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_53),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_54),
.B(n_7),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_56),
.B(n_7),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_125),
.B(n_130),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_56),
.B(n_13),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_40),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_29),
.Y(n_127)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_127),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_29),
.Y(n_128)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_42),
.Y(n_129)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_53),
.Y(n_130)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_36),
.Y(n_131)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_131),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_27),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_132),
.Y(n_174)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_57),
.Y(n_133)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_58),
.C(n_49),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_142),
.B(n_0),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_67),
.A2(n_49),
.B1(n_36),
.B2(n_42),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_143),
.A2(n_154),
.B1(n_157),
.B2(n_197),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_124),
.A2(n_42),
.B1(n_25),
.B2(n_45),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_145),
.A2(n_192),
.B1(n_33),
.B2(n_24),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_146),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_152),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_153),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_53),
.B1(n_42),
.B2(n_40),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_155),
.B(n_13),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_77),
.A2(n_47),
.B1(n_37),
.B2(n_55),
.Y(n_157)
);

INVx6_ASAP7_75t_SL g161 ( 
.A(n_96),
.Y(n_161)
);

INVx13_ASAP7_75t_L g305 ( 
.A(n_161),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_123),
.A2(n_58),
.B(n_33),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_163),
.B(n_164),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_69),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_121),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_168),
.B(n_169),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_133),
.B(n_46),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_190),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_78),
.B(n_47),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_110),
.A2(n_37),
.B1(n_55),
.B2(n_51),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_78),
.B(n_51),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_195),
.B(n_222),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_62),
.A2(n_46),
.B1(n_39),
.B2(n_45),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_64),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_198),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_128),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_219),
.Y(n_229)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_101),
.Y(n_205)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_111),
.Y(n_206)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_63),
.B(n_49),
.Y(n_219)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_73),
.B(n_39),
.C(n_25),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_114),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_87),
.B(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_103),
.Y(n_223)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_88),
.Y(n_225)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_196),
.A2(n_132),
.B1(n_105),
.B2(n_24),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_227),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_228),
.A2(n_271),
.B1(n_191),
.B2(n_202),
.Y(n_309)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_231),
.Y(n_362)
);

BUFx8_ASAP7_75t_L g234 ( 
.A(n_149),
.Y(n_234)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_234),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_151),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g353 ( 
.A(n_237),
.B(n_257),
.C(n_264),
.Y(n_353)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_239),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_136),
.Y(n_240)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_240),
.Y(n_335)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_246),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_219),
.A2(n_33),
.B1(n_24),
.B2(n_116),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_242),
.A2(n_245),
.B1(n_265),
.B2(n_275),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_186),
.A2(n_129),
.B1(n_71),
.B2(n_118),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_243),
.A2(n_277),
.B1(n_279),
.B2(n_288),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_136),
.Y(n_244)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_244),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_170),
.A2(n_68),
.B1(n_90),
.B2(n_131),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_213),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_137),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_248),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_137),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_249),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_61),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_250),
.B(n_254),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_183),
.Y(n_251)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_251),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_253),
.B(n_256),
.C(n_162),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_0),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_160),
.Y(n_255)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx2_ASAP7_75t_R g256 ( 
.A(n_138),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_0),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_259),
.B(n_297),
.Y(n_317)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_260),
.B(n_263),
.Y(n_320)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_175),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_174),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_193),
.A2(n_84),
.B1(n_79),
.B2(n_100),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_135),
.B(n_113),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_266),
.B(n_286),
.Y(n_327)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_138),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_267),
.B(n_269),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

BUFx24_ASAP7_75t_L g364 ( 
.A(n_268),
.Y(n_364)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_204),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_145),
.A2(n_82),
.B1(n_89),
.B2(n_81),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_199),
.Y(n_272)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_272),
.Y(n_312)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_208),
.Y(n_273)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_183),
.A2(n_59),
.B1(n_95),
.B2(n_91),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_147),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_276),
.B(n_281),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_220),
.A2(n_59),
.B1(n_97),
.B2(n_95),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_141),
.A2(n_59),
.B1(n_91),
.B2(n_43),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_147),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_282),
.Y(n_330)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_200),
.A2(n_106),
.B1(n_34),
.B2(n_43),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_284),
.A2(n_295),
.B1(n_177),
.B2(n_187),
.Y(n_313)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_150),
.Y(n_285)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_285),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_215),
.B(n_14),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_143),
.A2(n_34),
.B1(n_43),
.B2(n_2),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_176),
.Y(n_289)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_181),
.B(n_166),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_290),
.B(n_291),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_215),
.B(n_14),
.Y(n_291)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_207),
.Y(n_292)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_139),
.A2(n_34),
.B1(n_43),
.B2(n_2),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_293),
.A2(n_226),
.B1(n_167),
.B2(n_194),
.Y(n_322)
);

INVx11_ASAP7_75t_L g294 ( 
.A(n_134),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_294),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_140),
.A2(n_34),
.B1(n_43),
.B2(n_15),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_189),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_298),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_144),
.B(n_212),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_173),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_148),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_300),
.Y(n_351)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_184),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_301),
.B(n_303),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_212),
.B(n_0),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_0),
.Y(n_365)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_158),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_217),
.B(n_6),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_304),
.B(n_177),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_173),
.B(n_224),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_306),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_234),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_307),
.B(n_311),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_309),
.A2(n_322),
.B1(n_331),
.B2(n_339),
.Y(n_377)
);

AO22x1_ASAP7_75t_SL g310 ( 
.A1(n_252),
.A2(n_209),
.B1(n_208),
.B2(n_158),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_310),
.B(n_313),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_234),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_159),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_238),
.B(n_254),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_243),
.A2(n_209),
.B1(n_188),
.B2(n_202),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_329),
.A2(n_295),
.B1(n_303),
.B2(n_255),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_228),
.A2(n_188),
.B1(n_191),
.B2(n_167),
.Y(n_331)
);

NAND3xp33_ASAP7_75t_L g408 ( 
.A(n_333),
.B(n_340),
.C(n_305),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_270),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_337),
.B(n_349),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_232),
.A2(n_226),
.B1(n_194),
.B2(n_171),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_301),
.A2(n_178),
.B1(n_171),
.B2(n_187),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_342),
.A2(n_344),
.B1(n_350),
.B2(n_352),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_301),
.A2(n_178),
.B1(n_185),
.B2(n_208),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_259),
.B(n_184),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_302),
.A2(n_172),
.B1(n_165),
.B2(n_179),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_250),
.A2(n_172),
.B1(n_165),
.B2(n_134),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_306),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_356),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_229),
.A2(n_179),
.B1(n_148),
.B2(n_216),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_355),
.A2(n_360),
.B1(n_363),
.B2(n_230),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_306),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_297),
.A2(n_216),
.B1(n_162),
.B2(n_149),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_284),
.A2(n_134),
.B1(n_34),
.B2(n_153),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_365),
.B(n_2),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_235),
.B(n_1),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_1),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_233),
.B(n_289),
.C(n_285),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_368),
.B(n_274),
.Y(n_401)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_319),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_370),
.B(n_374),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_326),
.A2(n_288),
.B1(n_239),
.B2(n_283),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_371),
.A2(n_394),
.B1(n_405),
.B2(n_407),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_372),
.B(n_384),
.Y(n_434)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_337),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_336),
.B(n_235),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_376),
.B(n_406),
.Y(n_429)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_354),
.A2(n_256),
.B(n_251),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_379),
.A2(n_398),
.B(n_399),
.Y(n_421)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_338),
.Y(n_380)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_380),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g457 ( 
.A1(n_381),
.A2(n_398),
.B1(n_375),
.B2(n_378),
.Y(n_457)
);

INVx5_ASAP7_75t_SL g382 ( 
.A(n_307),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_382),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_319),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_383),
.B(n_392),
.Y(n_436)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_385),
.Y(n_442)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_338),
.Y(n_386)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_386),
.Y(n_450)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

INVx8_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

BUFx4f_ASAP7_75t_SL g390 ( 
.A(n_364),
.Y(n_390)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_390),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_317),
.B(n_272),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_391),
.B(n_396),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g392 ( 
.A(n_328),
.B(n_305),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_393),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_320),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_395),
.B(n_408),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_317),
.B(n_236),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_339),
.A2(n_230),
.B(n_299),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_356),
.A2(n_327),
.B(n_340),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_314),
.A2(n_329),
.B1(n_310),
.B2(n_323),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_400),
.A2(n_410),
.B1(n_331),
.B2(n_342),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_321),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_357),
.B(n_236),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_411),
.B(n_415),
.Y(n_444)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_314),
.A2(n_249),
.B1(n_240),
.B2(n_248),
.Y(n_410)
);

O2A1O1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_313),
.A2(n_261),
.B(n_258),
.C(n_247),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_336),
.B(n_296),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_412),
.B(n_414),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_365),
.B(n_287),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_416),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_320),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_323),
.A2(n_274),
.B(n_261),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_247),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_346),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_417),
.B(n_358),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_420),
.A2(n_456),
.B1(n_377),
.B2(n_394),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_328),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_428),
.C(n_430),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_388),
.A2(n_310),
.B1(n_327),
.B2(n_322),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_425),
.A2(n_433),
.B1(n_377),
.B2(n_407),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_400),
.A2(n_310),
.B1(n_344),
.B2(n_357),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_427),
.A2(n_432),
.B1(n_435),
.B2(n_440),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_341),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_341),
.C(n_368),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_388),
.A2(n_341),
.B1(n_350),
.B2(n_352),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_388),
.A2(n_353),
.B1(n_316),
.B2(n_308),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_363),
.B1(n_351),
.B2(n_316),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_SL g439 ( 
.A1(n_381),
.A2(n_373),
.B1(n_397),
.B2(n_385),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_389),
.A2(n_351),
.B1(n_293),
.B2(n_308),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_334),
.C(n_311),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_443),
.C(n_452),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_396),
.B(n_334),
.C(n_321),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_258),
.Y(n_489)
);

OAI32xp33_ASAP7_75t_L g448 ( 
.A1(n_391),
.A2(n_359),
.A3(n_347),
.B1(n_361),
.B2(n_358),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_448),
.B(n_394),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_359),
.Y(n_452)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_453),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_389),
.A2(n_282),
.B1(n_244),
.B2(n_330),
.Y(n_456)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_397),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_395),
.Y(n_464)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_461),
.A2(n_487),
.B1(n_433),
.B2(n_456),
.Y(n_527)
);

INVx13_ASAP7_75t_L g463 ( 
.A(n_437),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_464),
.B(n_483),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_425),
.A2(n_370),
.B1(n_383),
.B2(n_414),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_467),
.A2(n_450),
.B1(n_440),
.B2(n_449),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_421),
.A2(n_415),
.B(n_379),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_468),
.A2(n_472),
.B(n_478),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_441),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_469),
.B(n_479),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_453),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_470),
.B(n_476),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_421),
.A2(n_392),
.B(n_411),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_418),
.Y(n_473)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_473),
.Y(n_514)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_418),
.Y(n_474)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_423),
.Y(n_475)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_475),
.Y(n_520)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_423),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_SL g477 ( 
.A(n_446),
.B(n_380),
.C(n_386),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_477),
.B(n_480),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_444),
.A2(n_382),
.B(n_403),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_424),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_442),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_481),
.Y(n_505)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_448),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_485),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_458),
.B(n_412),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_420),
.A2(n_376),
.B1(n_413),
.B2(n_416),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_484),
.A2(n_482),
.B1(n_471),
.B2(n_483),
.Y(n_517)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_426),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_436),
.A2(n_403),
.B(n_417),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_452),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_427),
.A2(n_372),
.B1(n_384),
.B2(n_406),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_447),
.B(n_347),
.C(n_361),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_488),
.B(n_455),
.C(n_424),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_489),
.B(n_422),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_454),
.B(n_393),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_490),
.B(n_493),
.Y(n_513)
);

AOI21xp33_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_382),
.B(n_390),
.Y(n_491)
);

OAI21xp33_ASAP7_75t_L g523 ( 
.A1(n_491),
.A2(n_451),
.B(n_419),
.Y(n_523)
);

NAND2x1p5_ASAP7_75t_R g492 ( 
.A(n_444),
.B(n_390),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_492),
.A2(n_496),
.B(n_432),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_454),
.B(n_369),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_495),
.Y(n_511)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_450),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_498),
.B(n_499),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_428),
.Y(n_499)
);

OAI21xp33_ASAP7_75t_L g555 ( 
.A1(n_503),
.A2(n_523),
.B(n_364),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_504),
.A2(n_527),
.B1(n_461),
.B2(n_462),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_430),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_509),
.B(n_526),
.C(n_529),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_510),
.B(n_481),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_486),
.B(n_431),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_534),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_443),
.Y(n_515)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_515),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_465),
.Y(n_535)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_518),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_449),
.Y(n_519)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_519),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_429),
.Y(n_521)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_521),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_490),
.B(n_445),
.Y(n_522)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_522),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_488),
.B(n_442),
.Y(n_524)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_524),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_485),
.Y(n_525)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_525),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_484),
.A2(n_438),
.B1(n_435),
.B2(n_434),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_528),
.A2(n_533),
.B1(n_324),
.B2(n_330),
.Y(n_558)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_434),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_468),
.B(n_332),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_530),
.B(n_531),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_472),
.B(n_465),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_478),
.B(n_455),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_532),
.B(n_324),
.C(n_362),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_496),
.A2(n_451),
.B1(n_437),
.B2(n_405),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_494),
.B(n_362),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_535),
.B(n_557),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_493),
.Y(n_537)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_537),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_506),
.A2(n_459),
.B1(n_470),
.B2(n_471),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_539),
.A2(n_543),
.B1(n_556),
.B2(n_558),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_540),
.Y(n_585)
);

FAx1_ASAP7_75t_SL g542 ( 
.A(n_497),
.B(n_492),
.CI(n_491),
.CON(n_542),
.SN(n_542)
);

MAJIxp5_ASAP7_75t_SL g573 ( 
.A(n_542),
.B(n_531),
.C(n_508),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_506),
.A2(n_460),
.B1(n_462),
.B2(n_495),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_502),
.B(n_511),
.Y(n_545)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_545),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_509),
.B(n_460),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_546),
.B(n_553),
.Y(n_579)
);

XNOR2x1_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_533),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_502),
.A2(n_476),
.B1(n_475),
.B2(n_474),
.Y(n_549)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_549),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_505),
.Y(n_551)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_551),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_499),
.B(n_473),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_511),
.B(n_390),
.Y(n_554)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_554),
.Y(n_591)
);

CKINVDCx14_ASAP7_75t_R g590 ( 
.A(n_555),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_508),
.A2(n_463),
.B1(n_335),
.B2(n_366),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_507),
.A2(n_463),
.B(n_325),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_500),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_560),
.B(n_565),
.Y(n_596)
);

INVx13_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_563),
.B(n_498),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_497),
.A2(n_335),
.B1(n_366),
.B2(n_325),
.Y(n_564)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_564),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_526),
.B(n_312),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_528),
.A2(n_312),
.B1(n_231),
.B2(n_387),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_566),
.A2(n_501),
.B1(n_520),
.B2(n_516),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_517),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_569),
.B(n_577),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_532),
.C(n_529),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_575),
.C(n_595),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_573),
.B(n_584),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_583),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_559),
.B(n_530),
.C(n_507),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_536),
.B(n_513),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_567),
.B(n_541),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_594),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_SL g583 ( 
.A(n_548),
.B(n_519),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_568),
.Y(n_586)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_586),
.Y(n_600)
);

XNOR2xp5_ASAP7_75t_SL g587 ( 
.A(n_548),
.B(n_546),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_587),
.B(n_562),
.Y(n_618)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_588),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_550),
.A2(n_518),
.B1(n_500),
.B2(n_527),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_592),
.A2(n_576),
.B1(n_571),
.B2(n_552),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_537),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_553),
.B(n_520),
.C(n_516),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_596),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_598),
.B(n_599),
.Y(n_628)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_588),
.Y(n_599)
);

INVx13_ASAP7_75t_L g602 ( 
.A(n_589),
.Y(n_602)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_602),
.Y(n_625)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_572),
.B(n_563),
.C(n_538),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_603),
.B(n_612),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_585),
.A2(n_550),
.B1(n_535),
.B2(n_539),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_604),
.A2(n_607),
.B1(n_609),
.B2(n_364),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_591),
.A2(n_547),
.B(n_542),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_606),
.A2(n_364),
.B(n_300),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_582),
.A2(n_552),
.B1(n_545),
.B2(n_558),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_592),
.A2(n_576),
.B1(n_581),
.B2(n_570),
.Y(n_609)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_589),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_611),
.B(n_614),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_579),
.B(n_551),
.Y(n_612)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_578),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_615),
.A2(n_556),
.B1(n_513),
.B2(n_578),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_579),
.B(n_543),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_616),
.B(n_292),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_575),
.B(n_538),
.C(n_547),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_617),
.B(n_619),
.Y(n_621)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_618),
.B(n_387),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_587),
.B(n_557),
.C(n_554),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_573),
.B(n_566),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_620),
.B(n_584),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_597),
.B(n_595),
.C(n_574),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_622),
.B(n_626),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_623),
.B(n_636),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_606),
.A2(n_542),
.B(n_562),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_624),
.A2(n_635),
.B(n_614),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_610),
.B(n_593),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_627),
.A2(n_639),
.B1(n_607),
.B2(n_602),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_608),
.B(n_590),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_629),
.B(n_630),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_618),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_603),
.B(n_583),
.C(n_514),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_631),
.B(n_638),
.Y(n_644)
);

FAx1_ASAP7_75t_SL g633 ( 
.A(n_613),
.B(n_561),
.CI(n_514),
.CON(n_633),
.SN(n_633)
);

OAI22xp5_ASAP7_75t_SL g651 ( 
.A1(n_633),
.A2(n_624),
.B1(n_605),
.B2(n_627),
.Y(n_651)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_611),
.B(n_335),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g643 ( 
.A(n_637),
.B(n_619),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_600),
.B(n_273),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_617),
.B(n_268),
.C(n_294),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_641),
.B(n_601),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_622),
.B(n_630),
.C(n_631),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_642),
.B(n_645),
.Y(n_670)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_643),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_640),
.B(n_605),
.C(n_615),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_646),
.B(n_656),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_628),
.B(n_600),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g659 ( 
.A(n_647),
.B(n_649),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_621),
.A2(n_613),
.B(n_620),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_648),
.A2(n_641),
.B(n_637),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_625),
.B(n_609),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_651),
.A2(n_636),
.B1(n_633),
.B2(n_632),
.Y(n_661)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_652),
.B(n_280),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g656 ( 
.A(n_639),
.B(n_604),
.C(n_601),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_657),
.B(n_635),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_623),
.B(n_632),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_SL g671 ( 
.A(n_658),
.B(n_17),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_SL g678 ( 
.A1(n_661),
.A2(n_663),
.B1(n_664),
.B2(n_659),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_646),
.A2(n_657),
.B1(n_650),
.B2(n_654),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_662),
.B(n_665),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_642),
.A2(n_633),
.B(n_268),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_666),
.A2(n_667),
.B(n_668),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_644),
.A2(n_268),
.B(n_278),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_656),
.A2(n_280),
.B(n_278),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g679 ( 
.A(n_669),
.B(n_6),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_671),
.B(n_655),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_660),
.A2(n_651),
.B(n_653),
.Y(n_673)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_673),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_674),
.B(n_680),
.Y(n_684)
);

AOI322xp5_ASAP7_75t_L g676 ( 
.A1(n_670),
.A2(n_643),
.A3(n_653),
.B1(n_280),
.B2(n_278),
.C1(n_153),
.C2(n_152),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_SL g683 ( 
.A1(n_676),
.A2(n_16),
.B1(n_18),
.B2(n_2),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_SL g677 ( 
.A1(n_664),
.A2(n_15),
.B1(n_17),
.B2(n_5),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_677),
.A2(n_672),
.B(n_673),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_678),
.A2(n_679),
.B1(n_15),
.B2(n_16),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_665),
.B(n_6),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_675),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_681),
.B(n_682),
.Y(n_689)
);

MAJIxp5_ASAP7_75t_L g687 ( 
.A(n_683),
.B(n_685),
.C(n_677),
.Y(n_687)
);

XNOR2xp5_ASAP7_75t_L g690 ( 
.A(n_687),
.B(n_686),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_SL g688 ( 
.A1(n_681),
.A2(n_16),
.B(n_18),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_688),
.A2(n_684),
.B(n_3),
.Y(n_691)
);

XOR2xp5_ASAP7_75t_L g692 ( 
.A(n_690),
.B(n_691),
.Y(n_692)
);

MAJIxp5_ASAP7_75t_L g693 ( 
.A(n_692),
.B(n_689),
.C(n_3),
.Y(n_693)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_693),
.B(n_3),
.Y(n_694)
);

XOR2xp5_ASAP7_75t_L g695 ( 
.A(n_694),
.B(n_3),
.Y(n_695)
);


endmodule