module fake_ibex_1008_n_1892 (n_151, n_85, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_165, n_452, n_86, n_70, n_255, n_175, n_586, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_545, n_583, n_194, n_249, n_334, n_312, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_421, n_475, n_166, n_163, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_7, n_109, n_127, n_121, n_527, n_465, n_48, n_325, n_57, n_301, n_496, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_13, n_122, n_523, n_116, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_150, n_286, n_321, n_133, n_569, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_459, n_30, n_518, n_367, n_221, n_437, n_355, n_474, n_407, n_102, n_490, n_568, n_52, n_448, n_99, n_466, n_269, n_156, n_570, n_126, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_536, n_352, n_290, n_558, n_174, n_467, n_427, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_267, n_245, n_571, n_229, n_209, n_472, n_347, n_473, n_445, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_137, n_338, n_173, n_477, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_365, n_4, n_6, n_539, n_100, n_179, n_354, n_206, n_392, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_495, n_410, n_308, n_463, n_411, n_135, n_520, n_512, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_409, n_582, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_532, n_95, n_405, n_415, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_311, n_406, n_97, n_197, n_528, n_181, n_131, n_123, n_260, n_462, n_302, n_450, n_443, n_572, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_492, n_232, n_380, n_281, n_559, n_425, n_1892);

input n_151;
input n_85;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_165;
input n_452;
input n_86;
input n_70;
input n_255;
input n_175;
input n_586;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_194;
input n_249;
input n_334;
input n_312;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_421;
input n_475;
input n_166;
input n_163;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_13;
input n_122;
input n_523;
input n_116;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_437;
input n_355;
input n_474;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_536;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_267;
input n_245;
input n_571;
input n_229;
input n_209;
input n_472;
input n_347;
input n_473;
input n_445;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_137;
input n_338;
input n_173;
input n_477;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_365;
input n_4;
input n_6;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_495;
input n_410;
input n_308;
input n_463;
input n_411;
input n_135;
input n_520;
input n_512;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_409;
input n_582;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_532;
input n_95;
input n_405;
input n_415;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_260;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_492;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_1892;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_1308;
wire n_1138;
wire n_708;
wire n_1096;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_876;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_641;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_694;
wire n_787;
wire n_614;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_1155;
wire n_1292;
wire n_1576;
wire n_1664;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_1778;
wire n_646;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_605;
wire n_630;
wire n_1869;
wire n_1853;
wire n_745;
wire n_1753;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_709;
wire n_1296;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_606;
wire n_737;
wire n_1571;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_981;
wire n_1591;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_1036;
wire n_974;
wire n_1831;
wire n_608;
wire n_864;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_846;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_1334;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_1200;
wire n_1120;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_705;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1704;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_817;
wire n_951;
wire n_1580;
wire n_1574;
wire n_780;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_1785;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_628;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_887;
wire n_1162;
wire n_634;
wire n_961;
wire n_991;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_1323;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_595;
wire n_1001;
wire n_1396;
wire n_1224;
wire n_1538;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_1726;
wire n_830;
wire n_1241;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1337;
wire n_1647;
wire n_839;
wire n_768;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_1057;
wire n_1473;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_934;
wire n_775;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_815;
wire n_919;
wire n_681;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_1621;
wire n_1342;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_885;
wire n_1530;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1361;
wire n_1187;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_755;
wire n_1029;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1734;
wire n_1876;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_1262;
wire n_1692;
wire n_1012;
wire n_1805;
wire n_960;
wire n_689;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_1092;
wire n_1808;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1158;
wire n_763;
wire n_1882;
wire n_940;
wire n_1762;
wire n_1404;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_1333;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_1335;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_970;
wire n_921;
wire n_1534;
wire n_908;
wire n_1346;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_649;
wire n_1854;
wire n_866;

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_275),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_510),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_573),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_121),
.Y(n_590)
);

CKINVDCx14_ASAP7_75t_R g591 ( 
.A(n_529),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_422),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_60),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_54),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_455),
.Y(n_595)
);

INVx1_ASAP7_75t_SL g596 ( 
.A(n_295),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_47),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_185),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_440),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_103),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_539),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_102),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_46),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_143),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_571),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_332),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_346),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_217),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_338),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_434),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_266),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_72),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_80),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_184),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_403),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_557),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_547),
.Y(n_617)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_553),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_299),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_221),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_363),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_217),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_59),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_399),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_555),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_44),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_552),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_492),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_521),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_350),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_559),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_302),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_392),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_383),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_67),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_373),
.Y(n_637)
);

INVxp67_ASAP7_75t_R g638 ( 
.A(n_249),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_372),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_202),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_201),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_128),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_546),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_504),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_581),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_305),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_450),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_400),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_466),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_234),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_181),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_404),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_394),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_577),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_85),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_104),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_77),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_538),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_254),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_340),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_247),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_569),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_570),
.Y(n_663)
);

BUFx10_ASAP7_75t_L g664 ( 
.A(n_155),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_11),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_121),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_584),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_585),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_541),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_278),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_189),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_549),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_568),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_454),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_343),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_401),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_498),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_574),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_465),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_376),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_509),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_190),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_131),
.Y(n_684)
);

BUFx2_ASAP7_75t_L g685 ( 
.A(n_122),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_464),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_508),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_81),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_496),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_299),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_563),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_113),
.Y(n_692)
);

BUFx10_ASAP7_75t_L g693 ( 
.A(n_530),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_54),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_86),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_275),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_146),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_536),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_567),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_567),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_566),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_105),
.Y(n_702)
);

BUFx5_ASAP7_75t_L g703 ( 
.A(n_341),
.Y(n_703)
);

BUFx8_ASAP7_75t_SL g704 ( 
.A(n_365),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_488),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_572),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_124),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_244),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_519),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_409),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_544),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_499),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_172),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_450),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_579),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_562),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_354),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_59),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_20),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_290),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_556),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_92),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_239),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_540),
.Y(n_724)
);

INVx1_ASAP7_75t_SL g725 ( 
.A(n_56),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_514),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_522),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_277),
.Y(n_728)
);

BUFx10_ASAP7_75t_L g729 ( 
.A(n_505),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_389),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_30),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_468),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_235),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_534),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_582),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_576),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_28),
.Y(n_737)
);

BUFx5_ASAP7_75t_L g738 ( 
.A(n_561),
.Y(n_738)
);

BUFx10_ASAP7_75t_L g739 ( 
.A(n_580),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_457),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_382),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_139),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_506),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_480),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_159),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_331),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_192),
.Y(n_747)
);

CKINVDCx16_ASAP7_75t_R g748 ( 
.A(n_114),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_93),
.Y(n_749)
);

CKINVDCx14_ASAP7_75t_R g750 ( 
.A(n_507),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_283),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_143),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_351),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_537),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_560),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_202),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_491),
.Y(n_757)
);

BUFx10_ASAP7_75t_L g758 ( 
.A(n_272),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_565),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_497),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_308),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_550),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_479),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_548),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_31),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_303),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_467),
.Y(n_767)
);

BUFx10_ASAP7_75t_L g768 ( 
.A(n_205),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_502),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_426),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_462),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_272),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_493),
.Y(n_773)
);

BUFx10_ASAP7_75t_L g774 ( 
.A(n_517),
.Y(n_774)
);

BUFx10_ASAP7_75t_L g775 ( 
.A(n_554),
.Y(n_775)
);

BUFx10_ASAP7_75t_L g776 ( 
.A(n_55),
.Y(n_776)
);

INVx1_ASAP7_75t_SL g777 ( 
.A(n_544),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_423),
.Y(n_778)
);

CKINVDCx11_ASAP7_75t_R g779 ( 
.A(n_558),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_164),
.Y(n_780)
);

CKINVDCx14_ASAP7_75t_R g781 ( 
.A(n_583),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_524),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_575),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_494),
.Y(n_784)
);

CKINVDCx14_ASAP7_75t_R g785 ( 
.A(n_186),
.Y(n_785)
);

BUFx5_ASAP7_75t_L g786 ( 
.A(n_495),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_551),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_106),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_339),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_578),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_503),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_545),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_542),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_540),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_564),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_785),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_655),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_590),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_659),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_592),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_594),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_713),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_704),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_591),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_772),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_616),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_600),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_676),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_685),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_608),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_692),
.Y(n_811)
);

CKINVDCx20_ASAP7_75t_R g812 ( 
.A(n_620),
.Y(n_812)
);

CKINVDCx16_ASAP7_75t_R g813 ( 
.A(n_748),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_749),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_622),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_635),
.Y(n_817)
);

INVxp67_ASAP7_75t_SL g818 ( 
.A(n_661),
.Y(n_818)
);

INVxp33_ASAP7_75t_SL g819 ( 
.A(n_638),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_781),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_597),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_750),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_598),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_738),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_779),
.Y(n_825)
);

CKINVDCx20_ASAP7_75t_R g826 ( 
.A(n_671),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_675),
.B(n_0),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_691),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_587),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_633),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_627),
.B(n_1),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_717),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_695),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_712),
.B(n_2),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_641),
.Y(n_836)
);

INVxp33_ASAP7_75t_L g837 ( 
.A(n_588),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_602),
.Y(n_838)
);

INVxp67_ASAP7_75t_SL g839 ( 
.A(n_717),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_738),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_665),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_603),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_731),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_726),
.B(n_2),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_740),
.B(n_2),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_604),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_606),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_738),
.Y(n_848)
);

CKINVDCx16_ASAP7_75t_R g849 ( 
.A(n_599),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_609),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_736),
.B(n_3),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_610),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_751),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_612),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_613),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_615),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_853),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_846),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_797),
.B(n_799),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_814),
.B(n_751),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_818),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_815),
.B(n_766),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_852),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_813),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_846),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_840),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_848),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_798),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_833),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_829),
.B(n_664),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_839),
.Y(n_871)
);

CKINVDCx6p67_ASAP7_75t_R g872 ( 
.A(n_796),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_802),
.Y(n_873)
);

OA21x2_ASAP7_75t_L g874 ( 
.A1(n_821),
.A2(n_607),
.B(n_593),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_805),
.B(n_619),
.Y(n_875)
);

OA21x2_ASAP7_75t_L g876 ( 
.A1(n_823),
.A2(n_611),
.B(n_607),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_837),
.B(n_664),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_830),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_808),
.B(n_809),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_831),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_811),
.B(n_669),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_846),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_819),
.B(n_804),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_841),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_838),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_842),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_847),
.B(n_758),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_845),
.B(n_679),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_850),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_832),
.Y(n_891)
);

OA21x2_ASAP7_75t_L g892 ( 
.A1(n_835),
.A2(n_614),
.B(n_611),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_844),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_854),
.B(n_768),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_827),
.Y(n_895)
);

BUFx8_ASAP7_75t_L g896 ( 
.A(n_825),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_851),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_855),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_856),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_820),
.Y(n_900)
);

AND2x4_ASAP7_75t_L g901 ( 
.A(n_822),
.B(n_679),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_803),
.B(n_714),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_800),
.B(n_621),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_801),
.B(n_623),
.Y(n_904)
);

INVx3_ASAP7_75t_L g905 ( 
.A(n_807),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_810),
.B(n_714),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_812),
.B(n_626),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_816),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_817),
.Y(n_909)
);

AND2x4_ASAP7_75t_L g910 ( 
.A(n_826),
.B(n_764),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_834),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_843),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_846),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_797),
.B(n_764),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_849),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_806),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_846),
.Y(n_917)
);

INVxp67_ASAP7_75t_L g918 ( 
.A(n_852),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_828),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_849),
.B(n_703),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_806),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_828),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_828),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_814),
.B(n_780),
.Y(n_924)
);

AND2x6_ASAP7_75t_L g925 ( 
.A(n_814),
.B(n_780),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_806),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_828),
.B(n_631),
.Y(n_927)
);

XOR2xp5_ASAP7_75t_L g928 ( 
.A(n_798),
.B(n_770),
.Y(n_928)
);

CKINVDCx16_ASAP7_75t_R g929 ( 
.A(n_849),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_806),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_849),
.B(n_703),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_797),
.B(n_776),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_806),
.Y(n_933)
);

OA21x2_ASAP7_75t_L g934 ( 
.A1(n_824),
.A2(n_737),
.B(n_710),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_828),
.B(n_634),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_846),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_849),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_806),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_806),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_929),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_874),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_874),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_891),
.B(n_636),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_876),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_860),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_937),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_934),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_863),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_883),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_860),
.Y(n_950)
);

INVxp33_ASAP7_75t_L g951 ( 
.A(n_870),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_859),
.B(n_596),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_877),
.B(n_589),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_893),
.B(n_637),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_885),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_886),
.Y(n_956)
);

INVx1_ASAP7_75t_SL g957 ( 
.A(n_899),
.Y(n_957)
);

INVx5_ASAP7_75t_L g958 ( 
.A(n_860),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_927),
.B(n_639),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_895),
.Y(n_960)
);

BUFx10_ASAP7_75t_L g961 ( 
.A(n_864),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_861),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_921),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_892),
.Y(n_964)
);

INVxp67_ASAP7_75t_SL g965 ( 
.A(n_918),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_892),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_897),
.A2(n_697),
.B1(n_702),
.B2(n_696),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_935),
.B(n_640),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_933),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_862),
.Y(n_970)
);

OR2x2_ASAP7_75t_L g971 ( 
.A(n_903),
.B(n_725),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_938),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_932),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_857),
.B(n_642),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_904),
.B(n_907),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_869),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_880),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_871),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_884),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_926),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_939),
.Y(n_981)
);

OA22x2_ASAP7_75t_L g982 ( 
.A1(n_928),
.A2(n_648),
.B1(n_650),
.B2(n_646),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_924),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_919),
.B(n_651),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_868),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_914),
.B(n_881),
.Y(n_986)
);

AND2x6_ASAP7_75t_L g987 ( 
.A(n_888),
.B(n_753),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_925),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_922),
.B(n_652),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_923),
.B(n_653),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_887),
.Y(n_991)
);

BUFx4f_ASAP7_75t_L g992 ( 
.A(n_898),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_906),
.B(n_733),
.Y(n_993)
);

AND2x6_ASAP7_75t_L g994 ( 
.A(n_894),
.B(n_753),
.Y(n_994)
);

BUFx8_ASAP7_75t_SL g995 ( 
.A(n_905),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_872),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_896),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_901),
.B(n_660),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_910),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_916),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_910),
.B(n_666),
.Y(n_1001)
);

XNOR2xp5_ASAP7_75t_L g1002 ( 
.A(n_928),
.B(n_618),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_930),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_878),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_898),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_866),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_875),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_908),
.B(n_890),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_889),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_900),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_858),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_902),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_867),
.A2(n_756),
.B(n_752),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_920),
.B(n_931),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_858),
.Y(n_1016)
);

CKINVDCx16_ASAP7_75t_R g1017 ( 
.A(n_911),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_L g1018 ( 
.A(n_865),
.B(n_738),
.Y(n_1018)
);

INVx4_ASAP7_75t_SL g1019 ( 
.A(n_909),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_882),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_912),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_913),
.Y(n_1022)
);

OR2x6_ASAP7_75t_L g1023 ( 
.A(n_913),
.B(n_668),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_917),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_936),
.Y(n_1025)
);

INVx4_ASAP7_75t_SL g1026 ( 
.A(n_936),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_877),
.B(n_672),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_873),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_915),
.Y(n_1029)
);

INVx6_ASAP7_75t_L g1030 ( 
.A(n_915),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_874),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_877),
.B(n_789),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_859),
.A2(n_681),
.B1(n_683),
.B2(n_677),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_891),
.B(n_684),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_915),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_863),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1007),
.B(n_943),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_975),
.B(n_688),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_958),
.B(n_694),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_954),
.B(n_690),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_973),
.B(n_595),
.Y(n_1041)
);

AND2x4_ASAP7_75t_SL g1042 ( 
.A(n_961),
.B(n_724),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_958),
.B(n_707),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_957),
.B(n_724),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_946),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_945),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_962),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1034),
.B(n_708),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_945),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_976),
.B(n_978),
.Y(n_1050)
);

NOR2xp67_ASAP7_75t_L g1051 ( 
.A(n_991),
.B(n_4),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1033),
.B(n_718),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_953),
.A2(n_720),
.B1(n_722),
.B2(n_719),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_948),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_948),
.B(n_729),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_1030),
.B(n_668),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_950),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_1036),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_970),
.Y(n_1059)
);

OAI22x1_ASAP7_75t_R g1060 ( 
.A1(n_997),
.A2(n_769),
.B1(n_706),
.B2(n_730),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1019),
.B(n_617),
.Y(n_1061)
);

NOR3xp33_ASAP7_75t_L g1062 ( 
.A(n_1017),
.B(n_777),
.C(n_734),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_1036),
.B(n_1004),
.Y(n_1063)
);

BUFx8_ASAP7_75t_L g1064 ( 
.A(n_1004),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_1027),
.B(n_745),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_1032),
.B(n_746),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_971),
.B(n_747),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_964),
.Y(n_1068)
);

INVxp67_ASAP7_75t_L g1069 ( 
.A(n_993),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_953),
.B(n_761),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_959),
.B(n_968),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_966),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1001),
.B(n_765),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_941),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_SL g1075 ( 
.A(n_988),
.B(n_778),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_986),
.B(n_998),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_982),
.A2(n_794),
.B1(n_795),
.B2(n_793),
.Y(n_1077)
);

AOI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_967),
.A2(n_629),
.B1(n_632),
.B2(n_628),
.C(n_625),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1028),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_995),
.Y(n_1080)
);

INVx4_ASAP7_75t_SL g1081 ( 
.A(n_987),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_944),
.Y(n_1082)
);

INVx8_ASAP7_75t_L g1083 ( 
.A(n_1008),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_1023),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_1031),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_977),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_947),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_1002),
.B(n_630),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_992),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_960),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_1008),
.B(n_673),
.Y(n_1091)
);

INVx8_ASAP7_75t_L g1092 ( 
.A(n_994),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_SL g1093 ( 
.A(n_961),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_979),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_994),
.A2(n_604),
.B1(n_656),
.B2(n_624),
.Y(n_1095)
);

BUFx2_ASAP7_75t_SL g1096 ( 
.A(n_1029),
.Y(n_1096)
);

INVx5_ASAP7_75t_L g1097 ( 
.A(n_1023),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_SL g1098 ( 
.A1(n_1002),
.A2(n_985),
.B1(n_940),
.B2(n_996),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_999),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_974),
.B(n_644),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_984),
.B(n_645),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1000),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1009),
.A2(n_604),
.B1(n_656),
.B2(n_624),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_989),
.B(n_654),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_990),
.B(n_658),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1035),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1012),
.B(n_674),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1019),
.B(n_643),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_1015),
.B(n_686),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_949),
.B(n_739),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1005),
.B(n_687),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_980),
.B(n_673),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1021),
.B(n_744),
.Y(n_1113)
);

OR2x2_ASAP7_75t_L g1114 ( 
.A(n_981),
.B(n_698),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_963),
.B(n_700),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_981),
.B(n_701),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_1010),
.B(n_715),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_1003),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_969),
.B(n_716),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_972),
.B(n_721),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1006),
.A2(n_649),
.B1(n_662),
.B2(n_647),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1013),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_955),
.B(n_735),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_SL g1124 ( 
.A(n_1025),
.B(n_775),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1026),
.B(n_775),
.Y(n_1125)
);

BUFx3_ASAP7_75t_L g1126 ( 
.A(n_1020),
.Y(n_1126)
);

INVx8_ASAP7_75t_L g1127 ( 
.A(n_1020),
.Y(n_1127)
);

NAND2xp33_ASAP7_75t_L g1128 ( 
.A(n_1011),
.B(n_738),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1018),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_1011),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1011),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1016),
.B(n_743),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_1022),
.B(n_754),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1024),
.B(n_755),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_942),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_956),
.B(n_775),
.Y(n_1136)
);

NOR2xp67_ASAP7_75t_L g1137 ( 
.A(n_991),
.B(n_4),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1007),
.A2(n_723),
.B1(n_728),
.B2(n_657),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_952),
.B(n_757),
.Y(n_1139)
);

OAI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_956),
.A2(n_790),
.B1(n_791),
.B2(n_787),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_1031),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_965),
.A2(n_760),
.B1(n_762),
.B2(n_759),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1030),
.Y(n_1143)
);

AO22x2_ASAP7_75t_L g1144 ( 
.A1(n_956),
.A2(n_667),
.B1(n_670),
.B2(n_663),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_951),
.B(n_763),
.Y(n_1145)
);

NAND2xp33_ASAP7_75t_L g1146 ( 
.A(n_983),
.B(n_786),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_965),
.A2(n_771),
.B1(n_773),
.B2(n_767),
.Y(n_1147)
);

INVx8_ASAP7_75t_L g1148 ( 
.A(n_1008),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1014),
.A2(n_680),
.B(n_682),
.C(n_678),
.Y(n_1149)
);

AND2x6_ASAP7_75t_L g1150 ( 
.A(n_983),
.B(n_741),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_1030),
.Y(n_1151)
);

BUFx10_ASAP7_75t_L g1152 ( 
.A(n_1030),
.Y(n_1152)
);

OAI21xp33_ASAP7_75t_L g1153 ( 
.A1(n_1038),
.A2(n_705),
.B(n_699),
.Y(n_1153)
);

OAI21xp33_ASAP7_75t_L g1154 ( 
.A1(n_1067),
.A2(n_711),
.B(n_709),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1071),
.A2(n_732),
.B(n_727),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1073),
.A2(n_783),
.B(n_782),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1054),
.B(n_792),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1050),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1075),
.B(n_693),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1082),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1045),
.B(n_774),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_1088),
.B(n_784),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1047),
.B(n_786),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1085),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_1064),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1064),
.B(n_788),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1149),
.A2(n_6),
.B(n_4),
.C(n_5),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1056),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_1124),
.B(n_601),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1080),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1087),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1097),
.B(n_605),
.Y(n_1172)
);

OR2x2_ASAP7_75t_SL g1173 ( 
.A(n_1060),
.B(n_689),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1081),
.B(n_7),
.Y(n_1174)
);

NOR2xp67_ASAP7_75t_L g1175 ( 
.A(n_1089),
.B(n_8),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1127),
.Y(n_1176)
);

INVx3_ASAP7_75t_L g1177 ( 
.A(n_1127),
.Y(n_1177)
);

AOI22x1_ASAP7_75t_L g1178 ( 
.A1(n_1129),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1040),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1135),
.A2(n_12),
.B(n_13),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_1076),
.B(n_13),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_R g1182 ( 
.A(n_1096),
.B(n_14),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1081),
.B(n_15),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1068),
.A2(n_16),
.B(n_17),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_SL g1185 ( 
.A(n_1152),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_1085),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1048),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1140),
.B(n_19),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1079),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1072),
.A2(n_18),
.B(n_19),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1070),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_1191)
);

BUFx4f_ASAP7_75t_L g1192 ( 
.A(n_1092),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1112),
.Y(n_1193)
);

OR2x6_ASAP7_75t_L g1194 ( 
.A(n_1083),
.B(n_24),
.Y(n_1194)
);

INVx11_ASAP7_75t_L g1195 ( 
.A(n_1093),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1139),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1196)
);

INVx5_ASAP7_75t_L g1197 ( 
.A(n_1150),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1055),
.B(n_29),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1099),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1101),
.A2(n_32),
.B(n_33),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1053),
.B(n_32),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1148),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1062),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1086),
.A2(n_35),
.B(n_37),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1104),
.A2(n_38),
.B(n_39),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1141),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1102),
.B(n_1118),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1105),
.A2(n_38),
.B(n_39),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1094),
.Y(n_1209)
);

INVx6_ASAP7_75t_L g1210 ( 
.A(n_1151),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1041),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1144),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1113),
.B(n_45),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1052),
.A2(n_48),
.B(n_49),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1100),
.A2(n_49),
.B(n_50),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1044),
.B(n_51),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1136),
.B(n_52),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1091),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1078),
.B(n_53),
.Y(n_1219)
);

OR2x2_ASAP7_75t_L g1220 ( 
.A(n_1114),
.B(n_56),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_SL g1221 ( 
.A(n_1150),
.B(n_57),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1110),
.B(n_58),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1102),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1090),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_L g1225 ( 
.A(n_1095),
.B(n_61),
.C(n_62),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1109),
.A2(n_62),
.B(n_63),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1051),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1227)
);

INVx11_ASAP7_75t_L g1228 ( 
.A(n_1150),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1137),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1131),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1115),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1065),
.B(n_66),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1042),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1066),
.B(n_67),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1142),
.B(n_68),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1119),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_SL g1237 ( 
.A(n_1130),
.B(n_69),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1132),
.Y(n_1238)
);

INVx11_ASAP7_75t_L g1239 ( 
.A(n_1098),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1147),
.B(n_70),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1084),
.A2(n_74),
.B1(n_71),
.B2(n_73),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1126),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1134),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1046),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1046),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1121),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1145),
.B(n_76),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1138),
.A2(n_77),
.B(n_78),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1123),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1120),
.B(n_78),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1111),
.B(n_79),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1084),
.B(n_80),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1125),
.Y(n_1253)
);

INVx3_ASAP7_75t_L g1254 ( 
.A(n_1049),
.Y(n_1254)
);

INVx5_ASAP7_75t_L g1255 ( 
.A(n_1143),
.Y(n_1255)
);

AO21x1_ASAP7_75t_L g1256 ( 
.A1(n_1146),
.A2(n_452),
.B(n_451),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1106),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1057),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1039),
.A2(n_82),
.B(n_83),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1043),
.A2(n_83),
.B(n_84),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1107),
.B(n_83),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1061),
.B(n_1108),
.Y(n_1262)
);

AND2x6_ASAP7_75t_L g1263 ( 
.A(n_1059),
.B(n_87),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1061),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1108),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1128),
.A2(n_88),
.B(n_89),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1117),
.B(n_88),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1103),
.A2(n_90),
.B(n_91),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1116),
.Y(n_1269)
);

AND2x6_ASAP7_75t_SL g1270 ( 
.A(n_1133),
.B(n_93),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_SL g1271 ( 
.A(n_1058),
.B(n_95),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1038),
.B(n_94),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1127),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1064),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1069),
.B(n_96),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1071),
.A2(n_97),
.B(n_98),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1038),
.B(n_97),
.Y(n_1277)
);

BUFx8_ASAP7_75t_L g1278 ( 
.A(n_1093),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1038),
.B(n_99),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1069),
.B(n_100),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1038),
.B(n_101),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1064),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1050),
.Y(n_1283)
);

BUFx4f_ASAP7_75t_L g1284 ( 
.A(n_1092),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1038),
.B(n_106),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1069),
.B(n_107),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1071),
.A2(n_108),
.B(n_109),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1071),
.A2(n_108),
.B(n_109),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1058),
.B(n_111),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1069),
.B(n_110),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1071),
.A2(n_112),
.B(n_113),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1127),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1050),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1081),
.B(n_118),
.Y(n_1294)
);

BUFx4f_ASAP7_75t_L g1295 ( 
.A(n_1092),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1071),
.A2(n_119),
.B(n_120),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1074),
.Y(n_1297)
);

AND2x2_ASAP7_75t_SL g1298 ( 
.A(n_1075),
.B(n_123),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1127),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1038),
.B(n_125),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1038),
.B(n_126),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1081),
.B(n_127),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1080),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1097),
.B(n_128),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1071),
.A2(n_128),
.B(n_129),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1071),
.A2(n_129),
.B(n_130),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1122),
.A2(n_132),
.B(n_133),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1071),
.A2(n_132),
.B(n_133),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1144),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1071),
.A2(n_135),
.B(n_136),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1152),
.Y(n_1311)
);

OAI321xp33_ASAP7_75t_L g1312 ( 
.A1(n_1077),
.A2(n_140),
.A3(n_142),
.B1(n_137),
.B2(n_138),
.C(n_141),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_141),
.B1(n_138),
.B2(n_140),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_SL g1314 ( 
.A(n_1075),
.B(n_142),
.Y(n_1314)
);

INVxp67_ASAP7_75t_SL g1315 ( 
.A(n_1045),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1071),
.A2(n_143),
.B(n_144),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1038),
.B(n_144),
.Y(n_1317)
);

AND2x6_ASAP7_75t_L g1318 ( 
.A(n_1046),
.B(n_144),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1069),
.B(n_145),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_SL g1320 ( 
.A(n_1058),
.B(n_146),
.Y(n_1320)
);

BUFx4f_ASAP7_75t_L g1321 ( 
.A(n_1092),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1038),
.B(n_147),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1063),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1323)
);

AND2x2_ASAP7_75t_SL g1324 ( 
.A(n_1075),
.B(n_149),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1069),
.B(n_149),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1071),
.A2(n_150),
.B(n_151),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1058),
.B(n_153),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1071),
.A2(n_152),
.B(n_153),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1058),
.B(n_155),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1071),
.A2(n_154),
.B(n_155),
.Y(n_1330)
);

NOR3xp33_ASAP7_75t_L g1331 ( 
.A(n_1037),
.B(n_157),
.C(n_156),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1144),
.A2(n_159),
.B1(n_157),
.B2(n_158),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1050),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1071),
.A2(n_160),
.B(n_161),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1045),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1127),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1071),
.A2(n_161),
.B(n_162),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1071),
.A2(n_163),
.B(n_164),
.Y(n_1338)
);

OAI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1071),
.A2(n_165),
.B(n_166),
.Y(n_1339)
);

OAI321xp33_ASAP7_75t_L g1340 ( 
.A1(n_1077),
.A2(n_167),
.A3(n_169),
.B1(n_165),
.B2(n_166),
.C(n_168),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1071),
.A2(n_165),
.B(n_166),
.Y(n_1341)
);

NAND2x1_ASAP7_75t_L g1342 ( 
.A(n_1150),
.B(n_167),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1071),
.A2(n_167),
.B(n_168),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_SL g1344 ( 
.A(n_1075),
.B(n_170),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1071),
.A2(n_171),
.B(n_172),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1144),
.A2(n_174),
.B1(n_171),
.B2(n_173),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1071),
.A2(n_173),
.B(n_174),
.Y(n_1347)
);

NOR3xp33_ASAP7_75t_L g1348 ( 
.A(n_1037),
.B(n_177),
.C(n_176),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1038),
.B(n_175),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1063),
.B(n_178),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1038),
.B(n_178),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1071),
.A2(n_179),
.B(n_180),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1071),
.A2(n_182),
.B(n_183),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1058),
.B(n_188),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1038),
.B(n_187),
.Y(n_1355)
);

NAND2x1p5_ASAP7_75t_L g1356 ( 
.A(n_1097),
.B(n_191),
.Y(n_1356)
);

BUFx2_ASAP7_75t_L g1357 ( 
.A(n_1045),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1050),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_SL g1359 ( 
.A(n_1058),
.B(n_193),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1127),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1038),
.B(n_192),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1069),
.B(n_194),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1071),
.A2(n_194),
.B(n_195),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1127),
.Y(n_1364)
);

NAND2x1p5_ASAP7_75t_L g1365 ( 
.A(n_1097),
.B(n_195),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1071),
.A2(n_196),
.B(n_197),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1071),
.A2(n_198),
.B(n_199),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1050),
.Y(n_1368)
);

NOR2xp33_ASAP7_75t_L g1369 ( 
.A(n_1069),
.B(n_200),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1071),
.A2(n_200),
.B(n_201),
.Y(n_1370)
);

INVx5_ASAP7_75t_L g1371 ( 
.A(n_1299),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1158),
.B(n_1283),
.Y(n_1372)
);

BUFx8_ASAP7_75t_SL g1373 ( 
.A(n_1170),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1169),
.B(n_1314),
.Y(n_1374)
);

INVxp67_ASAP7_75t_L g1375 ( 
.A(n_1357),
.Y(n_1375)
);

OAI21xp33_ASAP7_75t_L g1376 ( 
.A1(n_1314),
.A2(n_203),
.B(n_204),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1253),
.B(n_204),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1164),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_SL g1379 ( 
.A(n_1274),
.B(n_206),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1253),
.B(n_207),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1364),
.Y(n_1381)
);

AO22x1_ASAP7_75t_L g1382 ( 
.A1(n_1278),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_1382)
);

O2A1O1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1153),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_L g1384 ( 
.A(n_1153),
.B(n_212),
.C(n_213),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1272),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1168),
.B(n_215),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1186),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1344),
.B(n_453),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1315),
.B(n_216),
.Y(n_1389)
);

AND2x2_ASAP7_75t_SL g1390 ( 
.A(n_1298),
.B(n_1324),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1168),
.B(n_218),
.Y(n_1391)
);

NOR3xp33_ASAP7_75t_SL g1392 ( 
.A(n_1166),
.B(n_219),
.C(n_220),
.Y(n_1392)
);

INVx3_ASAP7_75t_L g1393 ( 
.A(n_1282),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_SL g1394 ( 
.A(n_1344),
.B(n_455),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1237),
.B(n_456),
.Y(n_1395)
);

O2A1O1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1277),
.A2(n_224),
.B(n_222),
.C(n_223),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1279),
.A2(n_226),
.B(n_224),
.C(n_225),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1335),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1303),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1333),
.A2(n_227),
.B1(n_225),
.B2(n_226),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1160),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1237),
.B(n_456),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1218),
.B(n_228),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1155),
.A2(n_229),
.B(n_230),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1358),
.A2(n_229),
.B(n_230),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1189),
.Y(n_1406)
);

BUFx2_ASAP7_75t_R g1407 ( 
.A(n_1165),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1368),
.A2(n_231),
.B(n_232),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1194),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1194),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1224),
.Y(n_1411)
);

NAND2x1p5_ASAP7_75t_L g1412 ( 
.A(n_1192),
.B(n_1284),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1171),
.Y(n_1413)
);

NAND3xp33_ASAP7_75t_SL g1414 ( 
.A(n_1212),
.B(n_233),
.C(n_234),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1221),
.B(n_457),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1201),
.A2(n_238),
.B1(n_236),
.B2(n_237),
.Y(n_1416)
);

NOR2xp67_ASAP7_75t_L g1417 ( 
.A(n_1176),
.B(n_237),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_SL g1418 ( 
.A(n_1309),
.B(n_240),
.C(n_241),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1281),
.A2(n_241),
.B(n_242),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1193),
.B(n_458),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1309),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1285),
.A2(n_243),
.B(n_245),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1195),
.Y(n_1423)
);

AND2x6_ASAP7_75t_L g1424 ( 
.A(n_1174),
.B(n_248),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_R g1425 ( 
.A(n_1192),
.B(n_249),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1156),
.B(n_250),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1173),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_1427)
);

OAI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1313),
.A2(n_255),
.B1(n_252),
.B2(n_253),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1213),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1350),
.B(n_255),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1177),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1154),
.B(n_256),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1313),
.A2(n_1346),
.B1(n_1332),
.B2(n_1181),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1209),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1332),
.A2(n_259),
.B1(n_257),
.B2(n_258),
.Y(n_1435)
);

CKINVDCx8_ASAP7_75t_R g1436 ( 
.A(n_1270),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_SL g1437 ( 
.A(n_1175),
.B(n_459),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1273),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1346),
.A2(n_262),
.B1(n_260),
.B2(n_261),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1154),
.B(n_261),
.Y(n_1440)
);

AOI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1300),
.A2(n_262),
.B(n_263),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1301),
.A2(n_263),
.B(n_264),
.Y(n_1442)
);

CKINVDCx14_ASAP7_75t_R g1443 ( 
.A(n_1284),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1231),
.B(n_265),
.Y(n_1444)
);

NAND2xp33_ASAP7_75t_L g1445 ( 
.A(n_1263),
.B(n_265),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1317),
.A2(n_267),
.B(n_268),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1322),
.A2(n_267),
.B(n_269),
.Y(n_1447)
);

AOI222xp33_ASAP7_75t_L g1448 ( 
.A1(n_1182),
.A2(n_271),
.B1(n_273),
.B2(n_269),
.C1(n_270),
.C2(n_272),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1199),
.Y(n_1449)
);

INVx6_ASAP7_75t_L g1450 ( 
.A(n_1242),
.Y(n_1450)
);

NAND2x1p5_ASAP7_75t_L g1451 ( 
.A(n_1295),
.B(n_274),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1236),
.B(n_276),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1307),
.A2(n_277),
.B(n_278),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1273),
.Y(n_1454)
);

OAI21xp33_ASAP7_75t_L g1455 ( 
.A1(n_1247),
.A2(n_278),
.B(n_279),
.Y(n_1455)
);

NOR2x1_ASAP7_75t_L g1456 ( 
.A(n_1292),
.B(n_280),
.Y(n_1456)
);

OAI22x1_ASAP7_75t_L g1457 ( 
.A1(n_1227),
.A2(n_1229),
.B1(n_1356),
.B2(n_1304),
.Y(n_1457)
);

INVx3_ASAP7_75t_SL g1458 ( 
.A(n_1292),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1257),
.B(n_460),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1349),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1263),
.Y(n_1461)
);

INVx3_ASAP7_75t_SL g1462 ( 
.A(n_1336),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1162),
.B(n_282),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_SL g1464 ( 
.A(n_1257),
.B(n_461),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1351),
.A2(n_284),
.B(n_285),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1360),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1287),
.A2(n_288),
.B(n_286),
.C(n_287),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1275),
.B(n_289),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1360),
.B(n_289),
.Y(n_1469)
);

A2O1A1Ixp33_ASAP7_75t_L g1470 ( 
.A1(n_1288),
.A2(n_292),
.B(n_290),
.C(n_291),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1297),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1219),
.B(n_292),
.Y(n_1472)
);

A2O1A1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1291),
.A2(n_295),
.B(n_293),
.C(n_294),
.Y(n_1473)
);

AND2x6_ASAP7_75t_L g1474 ( 
.A(n_1174),
.B(n_293),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1197),
.B(n_1258),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1321),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1355),
.A2(n_298),
.B1(n_296),
.B2(n_297),
.Y(n_1477)
);

INVx5_ASAP7_75t_L g1478 ( 
.A(n_1263),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1243),
.B(n_1238),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1361),
.A2(n_300),
.B(n_301),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1232),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1249),
.B(n_306),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1269),
.B(n_306),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1239),
.Y(n_1484)
);

INVx5_ASAP7_75t_L g1485 ( 
.A(n_1318),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1280),
.B(n_307),
.Y(n_1486)
);

INVx3_ASAP7_75t_L g1487 ( 
.A(n_1185),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1365),
.B(n_1233),
.Y(n_1488)
);

BUFx12f_ASAP7_75t_L g1489 ( 
.A(n_1202),
.Y(n_1489)
);

NOR3xp33_ASAP7_75t_SL g1490 ( 
.A(n_1312),
.B(n_309),
.C(n_310),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1286),
.B(n_310),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1210),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1290),
.A2(n_313),
.B1(n_311),
.B2(n_312),
.Y(n_1493)
);

NAND2x1_ASAP7_75t_L g1494 ( 
.A(n_1318),
.B(n_312),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1210),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1220),
.B(n_314),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1319),
.B(n_315),
.Y(n_1497)
);

NAND2x1p5_ASAP7_75t_L g1498 ( 
.A(n_1197),
.B(n_1183),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1163),
.A2(n_316),
.B(n_317),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1325),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_1500)
);

NOR3xp33_ASAP7_75t_L g1501 ( 
.A(n_1167),
.B(n_317),
.C(n_318),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1318),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1331),
.B(n_320),
.C(n_321),
.Y(n_1503)
);

OAI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1246),
.A2(n_322),
.B1(n_320),
.B2(n_321),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1252),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1362),
.B(n_323),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1262),
.B(n_324),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1369),
.B(n_325),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1246),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1229),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1269),
.B(n_330),
.Y(n_1511)
);

INVx4_ASAP7_75t_L g1512 ( 
.A(n_1228),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1222),
.B(n_333),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1203),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_1514)
);

OAI22x1_ASAP7_75t_L g1515 ( 
.A1(n_1178),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_SL g1516 ( 
.A(n_1340),
.B(n_337),
.C(n_338),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1270),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1294),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1250),
.A2(n_342),
.B(n_343),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1261),
.A2(n_345),
.B(n_342),
.C(n_344),
.Y(n_1520)
);

INVx5_ASAP7_75t_L g1521 ( 
.A(n_1206),
.Y(n_1521)
);

INVx3_ASAP7_75t_L g1522 ( 
.A(n_1207),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1265),
.B(n_347),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1157),
.B(n_347),
.Y(n_1524)
);

INVx4_ASAP7_75t_L g1525 ( 
.A(n_1302),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1198),
.B(n_348),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1161),
.B(n_349),
.Y(n_1527)
);

NOR3x1_ASAP7_75t_L g1528 ( 
.A(n_1159),
.B(n_351),
.C(n_349),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1339),
.B(n_462),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_SL g1530 ( 
.A(n_1347),
.B(n_463),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1311),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1352),
.B(n_463),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1216),
.B(n_350),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1293),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1217),
.B(n_352),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1367),
.A2(n_355),
.B1(n_353),
.B2(n_354),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1370),
.A2(n_356),
.B1(n_353),
.B2(n_355),
.Y(n_1537)
);

O2A1O1Ixp33_ASAP7_75t_L g1538 ( 
.A1(n_1234),
.A2(n_358),
.B(n_356),
.C(n_357),
.Y(n_1538)
);

AND2x4_ASAP7_75t_L g1539 ( 
.A(n_1264),
.B(n_359),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1211),
.A2(n_361),
.B1(n_359),
.B2(n_360),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1348),
.A2(n_365),
.B1(n_362),
.B2(n_364),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1235),
.B(n_364),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1240),
.B(n_366),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1255),
.Y(n_1544)
);

O2A1O1Ixp5_ASAP7_75t_L g1545 ( 
.A1(n_1172),
.A2(n_369),
.B(n_367),
.C(n_368),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1241),
.Y(n_1546)
);

OR2x6_ASAP7_75t_L g1547 ( 
.A(n_1342),
.B(n_370),
.Y(n_1547)
);

NAND3xp33_ASAP7_75t_SL g1548 ( 
.A(n_1191),
.B(n_371),
.C(n_373),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1204),
.A2(n_374),
.B(n_375),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1223),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1200),
.A2(n_377),
.B(n_378),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1223),
.B(n_1244),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1205),
.A2(n_377),
.B(n_378),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1271),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1208),
.A2(n_379),
.B(n_380),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1390),
.A2(n_1323),
.B1(n_1214),
.B2(n_1225),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1433),
.A2(n_1188),
.B1(n_1267),
.B2(n_1251),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1373),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1372),
.B(n_1289),
.Y(n_1559)
);

NOR2xp67_ASAP7_75t_L g1560 ( 
.A(n_1371),
.B(n_1381),
.Y(n_1560)
);

A2O1A1Ixp33_ASAP7_75t_L g1561 ( 
.A1(n_1445),
.A2(n_1196),
.B(n_1179),
.C(n_1187),
.Y(n_1561)
);

NOR2xp67_ASAP7_75t_L g1562 ( 
.A(n_1371),
.B(n_1215),
.Y(n_1562)
);

NOR2xp67_ASAP7_75t_R g1563 ( 
.A(n_1410),
.B(n_1244),
.Y(n_1563)
);

BUFx8_ASAP7_75t_L g1564 ( 
.A(n_1399),
.Y(n_1564)
);

AOI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1374),
.A2(n_1256),
.B(n_1180),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1453),
.A2(n_1190),
.B(n_1184),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1479),
.B(n_1276),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1478),
.B(n_1248),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1479),
.B(n_1296),
.Y(n_1569)
);

AO31x2_ASAP7_75t_L g1570 ( 
.A1(n_1457),
.A2(n_1266),
.A3(n_1306),
.B(n_1305),
.Y(n_1570)
);

AND3x2_ASAP7_75t_L g1571 ( 
.A(n_1409),
.B(n_1268),
.C(n_381),
.Y(n_1571)
);

AO31x2_ASAP7_75t_L g1572 ( 
.A1(n_1515),
.A2(n_1308),
.A3(n_1316),
.B(n_1310),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1475),
.A2(n_1254),
.B(n_1245),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_R g1574 ( 
.A(n_1410),
.B(n_1484),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1412),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1529),
.A2(n_1328),
.B(n_1326),
.Y(n_1576)
);

AO22x2_ASAP7_75t_L g1577 ( 
.A1(n_1510),
.A2(n_1320),
.B1(n_1329),
.B2(n_1327),
.Y(n_1577)
);

INVx4_ASAP7_75t_L g1578 ( 
.A(n_1458),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_SL g1579 ( 
.A(n_1478),
.B(n_1330),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_SL g1580 ( 
.A1(n_1494),
.A2(n_1402),
.B(n_1395),
.C(n_1394),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1485),
.B(n_1461),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1530),
.A2(n_1337),
.B(n_1334),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1376),
.A2(n_1353),
.B(n_1345),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1406),
.Y(n_1584)
);

AO22x2_ASAP7_75t_L g1585 ( 
.A1(n_1421),
.A2(n_1359),
.B1(n_1354),
.B2(n_1338),
.Y(n_1585)
);

OAI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1448),
.A2(n_1343),
.B(n_1341),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1532),
.A2(n_1366),
.B(n_1363),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1398),
.Y(n_1588)
);

NAND2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1485),
.B(n_1245),
.Y(n_1589)
);

O2A1O1Ixp33_ASAP7_75t_SL g1590 ( 
.A1(n_1388),
.A2(n_1470),
.B(n_1473),
.C(n_1467),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1502),
.A2(n_1415),
.B(n_1534),
.Y(n_1591)
);

BUFx6f_ASAP7_75t_L g1592 ( 
.A(n_1462),
.Y(n_1592)
);

BUFx10_ASAP7_75t_L g1593 ( 
.A(n_1423),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1489),
.Y(n_1594)
);

AOI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1554),
.A2(n_1226),
.B1(n_1260),
.B2(n_1259),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1512),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1501),
.A2(n_1230),
.B1(n_382),
.B2(n_381),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1512),
.Y(n_1598)
);

BUFx2_ASAP7_75t_R g1599 ( 
.A(n_1436),
.Y(n_1599)
);

AOI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1505),
.A2(n_383),
.B(n_384),
.Y(n_1600)
);

AOI221x1_ASAP7_75t_L g1601 ( 
.A1(n_1384),
.A2(n_1455),
.B1(n_1435),
.B2(n_1439),
.C(n_1428),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1488),
.B(n_385),
.Y(n_1602)
);

OR2x6_ASAP7_75t_L g1603 ( 
.A(n_1451),
.B(n_386),
.Y(n_1603)
);

AO32x2_ASAP7_75t_L g1604 ( 
.A1(n_1427),
.A2(n_389),
.A3(n_387),
.B1(n_388),
.B2(n_390),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1518),
.A2(n_393),
.B1(n_391),
.B2(n_392),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1424),
.A2(n_394),
.B1(n_391),
.B2(n_393),
.Y(n_1606)
);

OAI21x1_ASAP7_75t_L g1607 ( 
.A1(n_1498),
.A2(n_396),
.B(n_395),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1434),
.Y(n_1608)
);

AOI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1546),
.A2(n_397),
.B(n_398),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1424),
.A2(n_1474),
.B1(n_1514),
.B2(n_1426),
.Y(n_1610)
);

OAI22x1_ASAP7_75t_L g1611 ( 
.A1(n_1517),
.A2(n_403),
.B1(n_401),
.B2(n_402),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1496),
.B(n_401),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1525),
.A2(n_406),
.B1(n_404),
.B2(n_405),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1401),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1414),
.A2(n_409),
.B1(n_407),
.B2(n_408),
.Y(n_1615)
);

OA21x2_ASAP7_75t_L g1616 ( 
.A1(n_1545),
.A2(n_407),
.B(n_408),
.Y(n_1616)
);

AO31x2_ASAP7_75t_L g1617 ( 
.A1(n_1536),
.A2(n_412),
.A3(n_410),
.B(n_411),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1418),
.A2(n_414),
.B1(n_411),
.B2(n_413),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1413),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1424),
.A2(n_415),
.B1(n_411),
.B2(n_414),
.Y(n_1620)
);

BUFx6f_ASAP7_75t_L g1621 ( 
.A(n_1521),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1463),
.B(n_416),
.Y(n_1622)
);

AO31x2_ASAP7_75t_L g1623 ( 
.A1(n_1537),
.A2(n_419),
.A3(n_417),
.B(n_418),
.Y(n_1623)
);

AO32x2_ASAP7_75t_L g1624 ( 
.A1(n_1504),
.A2(n_420),
.A3(n_418),
.B1(n_419),
.B2(n_421),
.Y(n_1624)
);

BUFx6f_ASAP7_75t_L g1625 ( 
.A(n_1521),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1503),
.A2(n_420),
.B(n_421),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1531),
.Y(n_1627)
);

INVx1_ASAP7_75t_SL g1628 ( 
.A(n_1407),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1472),
.B(n_424),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1526),
.A2(n_1535),
.B(n_1533),
.Y(n_1630)
);

AND2x6_ASAP7_75t_L g1631 ( 
.A(n_1539),
.B(n_425),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1521),
.Y(n_1632)
);

O2A1O1Ixp33_ASAP7_75t_SL g1633 ( 
.A1(n_1437),
.A2(n_428),
.B(n_426),
.C(n_427),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1549),
.A2(n_429),
.B(n_430),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1471),
.A2(n_431),
.B(n_432),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1438),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1469),
.B(n_433),
.Y(n_1637)
);

INVx4_ASAP7_75t_L g1638 ( 
.A(n_1393),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1476),
.Y(n_1639)
);

INVxp67_ASAP7_75t_L g1640 ( 
.A(n_1411),
.Y(n_1640)
);

CKINVDCx20_ASAP7_75t_R g1641 ( 
.A(n_1443),
.Y(n_1641)
);

AOI221xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1509),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.C(n_438),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1548),
.A2(n_437),
.B1(n_435),
.B2(n_436),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1404),
.A2(n_441),
.B(n_439),
.C(n_440),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1547),
.B(n_439),
.Y(n_1645)
);

AO31x2_ASAP7_75t_L g1646 ( 
.A1(n_1432),
.A2(n_441),
.A3(n_439),
.B(n_440),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1499),
.A2(n_441),
.B(n_442),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1538),
.A2(n_1520),
.B(n_1385),
.C(n_1396),
.Y(n_1648)
);

AOI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1441),
.A2(n_444),
.B1(n_442),
.B2(n_443),
.C(n_445),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1389),
.B(n_443),
.Y(n_1650)
);

NAND3xp33_ASAP7_75t_L g1651 ( 
.A(n_1392),
.B(n_444),
.C(n_445),
.Y(n_1651)
);

AO31x2_ASAP7_75t_L g1652 ( 
.A1(n_1440),
.A2(n_448),
.A3(n_446),
.B(n_447),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_SL g1653 ( 
.A(n_1425),
.B(n_447),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1378),
.A2(n_448),
.B(n_449),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1378),
.A2(n_448),
.B(n_449),
.Y(n_1655)
);

NOR2xp67_ASAP7_75t_L g1656 ( 
.A(n_1544),
.B(n_449),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_SL g1657 ( 
.A1(n_1419),
.A2(n_469),
.B(n_470),
.Y(n_1657)
);

INVx5_ASAP7_75t_L g1658 ( 
.A(n_1474),
.Y(n_1658)
);

NAND2x1_ASAP7_75t_L g1659 ( 
.A(n_1474),
.B(n_1547),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1450),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1449),
.B(n_586),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1468),
.B(n_471),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1375),
.Y(n_1663)
);

CKINVDCx14_ASAP7_75t_R g1664 ( 
.A(n_1641),
.Y(n_1664)
);

BUFx2_ASAP7_75t_SL g1665 ( 
.A(n_1560),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1592),
.Y(n_1666)
);

INVx11_ASAP7_75t_L g1667 ( 
.A(n_1564),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1645),
.A2(n_1541),
.B1(n_1507),
.B2(n_1481),
.Y(n_1668)
);

NAND2x1p5_ASAP7_75t_L g1669 ( 
.A(n_1578),
.B(n_1379),
.Y(n_1669)
);

BUFx10_ASAP7_75t_L g1670 ( 
.A(n_1594),
.Y(n_1670)
);

OAI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1429),
.B1(n_1416),
.B2(n_1417),
.Y(n_1671)
);

INVx4_ASAP7_75t_L g1672 ( 
.A(n_1594),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1610),
.A2(n_1516),
.B1(n_1490),
.B2(n_1456),
.Y(n_1673)
);

CKINVDCx20_ASAP7_75t_R g1674 ( 
.A(n_1558),
.Y(n_1674)
);

BUFx10_ASAP7_75t_L g1675 ( 
.A(n_1602),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1556),
.A2(n_1508),
.B1(n_1486),
.B2(n_1540),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1614),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1621),
.Y(n_1678)
);

BUFx10_ASAP7_75t_L g1679 ( 
.A(n_1602),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1621),
.Y(n_1680)
);

INVx5_ASAP7_75t_L g1681 ( 
.A(n_1603),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1631),
.A2(n_1523),
.B1(n_1391),
.B2(n_1386),
.Y(n_1682)
);

INVx2_ASAP7_75t_SL g1683 ( 
.A(n_1593),
.Y(n_1683)
);

OAI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1658),
.A2(n_1400),
.B1(n_1500),
.B2(n_1493),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1619),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_SL g1686 ( 
.A1(n_1631),
.A2(n_1380),
.B1(n_1377),
.B2(n_1422),
.Y(n_1686)
);

AOI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1631),
.A2(n_1480),
.B1(n_1465),
.B2(n_1483),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1653),
.A2(n_1511),
.B1(n_1460),
.B2(n_1477),
.Y(n_1688)
);

INVx6_ASAP7_75t_L g1689 ( 
.A(n_1638),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1627),
.Y(n_1690)
);

AOI22x1_ASAP7_75t_SL g1691 ( 
.A1(n_1628),
.A2(n_1487),
.B1(n_1382),
.B2(n_1528),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1608),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1557),
.A2(n_1420),
.B1(n_1527),
.B2(n_1497),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1625),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1577),
.A2(n_1506),
.B1(n_1491),
.B2(n_1403),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1632),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1636),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1606),
.A2(n_1464),
.B1(n_1459),
.B2(n_1430),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1575),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1596),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1571),
.A2(n_1542),
.B1(n_1543),
.B2(n_1519),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1598),
.Y(n_1702)
);

OAI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1620),
.A2(n_1656),
.B1(n_1615),
.B2(n_1618),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1597),
.A2(n_1442),
.B1(n_1447),
.B2(n_1446),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1588),
.Y(n_1705)
);

CKINVDCx11_ASAP7_75t_R g1706 ( 
.A(n_1599),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1639),
.Y(n_1707)
);

INVx3_ASAP7_75t_L g1708 ( 
.A(n_1589),
.Y(n_1708)
);

CKINVDCx20_ASAP7_75t_R g1709 ( 
.A(n_1663),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1586),
.A2(n_1452),
.B1(n_1482),
.B2(n_1444),
.Y(n_1710)
);

BUFx2_ASAP7_75t_L g1711 ( 
.A(n_1574),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1584),
.Y(n_1712)
);

BUFx12f_ASAP7_75t_L g1713 ( 
.A(n_1637),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1652),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1559),
.B(n_1522),
.Y(n_1715)
);

INVx2_ASAP7_75t_SL g1716 ( 
.A(n_1660),
.Y(n_1716)
);

BUFx2_ASAP7_75t_SL g1717 ( 
.A(n_1562),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1652),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1601),
.A2(n_1513),
.B1(n_1405),
.B2(n_1408),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1635),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1644),
.A2(n_1383),
.B1(n_1524),
.B2(n_1397),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_SL g1722 ( 
.A1(n_1657),
.A2(n_1550),
.B1(n_1552),
.B2(n_1495),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1640),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1646),
.Y(n_1724)
);

OAI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1643),
.A2(n_1651),
.B1(n_1648),
.B2(n_1561),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1612),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1662),
.Y(n_1727)
);

BUFx12f_ASAP7_75t_L g1728 ( 
.A(n_1650),
.Y(n_1728)
);

INVx6_ASAP7_75t_L g1729 ( 
.A(n_1622),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1617),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_SL g1731 ( 
.A1(n_1585),
.A2(n_1552),
.B1(n_1492),
.B2(n_1387),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1607),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1649),
.A2(n_1551),
.B1(n_1555),
.B2(n_1553),
.Y(n_1733)
);

INVx6_ASAP7_75t_L g1734 ( 
.A(n_1563),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_1616),
.Y(n_1735)
);

BUFx8_ASAP7_75t_L g1736 ( 
.A(n_1604),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1611),
.A2(n_1454),
.B1(n_1466),
.B2(n_1431),
.Y(n_1737)
);

CKINVDCx6p67_ASAP7_75t_R g1738 ( 
.A(n_1581),
.Y(n_1738)
);

CKINVDCx11_ASAP7_75t_R g1739 ( 
.A(n_1605),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1712),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1689),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1730),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1739),
.A2(n_1568),
.B1(n_1626),
.B2(n_1647),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1725),
.A2(n_1630),
.B(n_1634),
.Y(n_1744)
);

NOR2x1_ASAP7_75t_SL g1745 ( 
.A(n_1665),
.B(n_1579),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1677),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1668),
.A2(n_1736),
.B1(n_1687),
.B2(n_1684),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1697),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1727),
.B(n_1705),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1720),
.A2(n_1591),
.B(n_1565),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1734),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1685),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1734),
.Y(n_1753)
);

INVx3_ASAP7_75t_L g1754 ( 
.A(n_1738),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1681),
.B(n_1567),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1703),
.A2(n_1642),
.B1(n_1595),
.B2(n_1613),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1724),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1681),
.B(n_1569),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1714),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1718),
.Y(n_1760)
);

CKINVDCx20_ASAP7_75t_R g1761 ( 
.A(n_1674),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1692),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1700),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1702),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1678),
.B(n_1623),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1696),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1729),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1729),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1735),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1680),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1695),
.A2(n_1566),
.B(n_1573),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1694),
.Y(n_1772)
);

AND2x2_ASAP7_75t_L g1773 ( 
.A(n_1715),
.B(n_1661),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1675),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1679),
.Y(n_1775)
);

AND2x4_ASAP7_75t_L g1776 ( 
.A(n_1711),
.B(n_1570),
.Y(n_1776)
);

BUFx2_ASAP7_75t_L g1777 ( 
.A(n_1709),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1716),
.B(n_1624),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1732),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1690),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1732),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1717),
.Y(n_1782)
);

OR2x6_ASAP7_75t_L g1783 ( 
.A(n_1748),
.B(n_1669),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1761),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1749),
.B(n_1728),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1747),
.A2(n_1673),
.B1(n_1671),
.B2(n_1737),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1741),
.B(n_1672),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1744),
.A2(n_1686),
.B(n_1726),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1767),
.B(n_1666),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1768),
.B(n_1731),
.Y(n_1790)
);

OAI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1743),
.A2(n_1682),
.B1(n_1723),
.B2(n_1676),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1756),
.A2(n_1701),
.B1(n_1710),
.B2(n_1691),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1754),
.A2(n_1664),
.B(n_1683),
.C(n_1708),
.Y(n_1793)
);

AND2x4_ASAP7_75t_SL g1794 ( 
.A(n_1763),
.B(n_1670),
.Y(n_1794)
);

NOR2x1_ASAP7_75t_SL g1795 ( 
.A(n_1782),
.B(n_1713),
.Y(n_1795)
);

AND2x4_ASAP7_75t_L g1796 ( 
.A(n_1776),
.B(n_1707),
.Y(n_1796)
);

AO21x2_ASAP7_75t_L g1797 ( 
.A1(n_1781),
.A2(n_1719),
.B(n_1609),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1755),
.A2(n_1693),
.B1(n_1721),
.B2(n_1698),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1745),
.A2(n_1580),
.B(n_1590),
.Y(n_1799)
);

A2O1A1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1751),
.A2(n_1688),
.B(n_1722),
.C(n_1600),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1746),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1772),
.B(n_1699),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1780),
.B(n_1706),
.Y(n_1803)
);

INVx4_ASAP7_75t_L g1804 ( 
.A(n_1753),
.Y(n_1804)
);

NOR2xp67_ASAP7_75t_L g1805 ( 
.A(n_1774),
.B(n_1775),
.Y(n_1805)
);

CKINVDCx11_ASAP7_75t_R g1806 ( 
.A(n_1777),
.Y(n_1806)
);

BUFx2_ASAP7_75t_L g1807 ( 
.A(n_1770),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1807),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1796),
.B(n_1769),
.Y(n_1809)
);

AO22x1_ASAP7_75t_L g1810 ( 
.A1(n_1796),
.A2(n_1758),
.B1(n_1765),
.B2(n_1778),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1805),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1801),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1789),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1787),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_SL g1815 ( 
.A1(n_1795),
.A2(n_1745),
.B1(n_1765),
.B2(n_1764),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1802),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1790),
.B(n_1785),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1804),
.B(n_1762),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1798),
.B(n_1740),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1783),
.Y(n_1820)
);

INVx5_ASAP7_75t_L g1821 ( 
.A(n_1783),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_L g1822 ( 
.A1(n_1788),
.A2(n_1792),
.B1(n_1791),
.B2(n_1786),
.Y(n_1822)
);

AND2x4_ASAP7_75t_L g1823 ( 
.A(n_1794),
.B(n_1779),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1806),
.B(n_1773),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1784),
.Y(n_1825)
);

NOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1793),
.B(n_1803),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1797),
.B(n_1752),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1811),
.B(n_1771),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1821),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1809),
.B(n_1742),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1825),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1812),
.Y(n_1832)
);

AOI31xp33_ASAP7_75t_L g1833 ( 
.A1(n_1826),
.A2(n_1799),
.A3(n_1667),
.B(n_1800),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1821),
.A2(n_1814),
.B1(n_1822),
.B2(n_1815),
.Y(n_1834)
);

AO31x2_ASAP7_75t_L g1835 ( 
.A1(n_1820),
.A2(n_1759),
.A3(n_1760),
.B(n_1757),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1808),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1827),
.Y(n_1837)
);

OAI211xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1819),
.A2(n_1704),
.B(n_1629),
.C(n_1733),
.Y(n_1838)
);

AOI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1810),
.A2(n_1766),
.B(n_1633),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1821),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1816),
.B(n_1750),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1818),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1817),
.A2(n_1655),
.B1(n_1654),
.B2(n_1583),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1840),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1833),
.B(n_1813),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1836),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1835),
.Y(n_1847)
);

NOR2xp67_ASAP7_75t_L g1848 ( 
.A(n_1834),
.B(n_1824),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1829),
.B(n_1823),
.Y(n_1849)
);

BUFx3_ASAP7_75t_L g1850 ( 
.A(n_1831),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1835),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1828),
.B(n_1572),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1850),
.B(n_1837),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1850),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1846),
.Y(n_1855)
);

AOI22xp5_ASAP7_75t_L g1856 ( 
.A1(n_1848),
.A2(n_1830),
.B1(n_1842),
.B2(n_1838),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1844),
.B(n_1832),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1849),
.Y(n_1858)
);

OAI211xp5_ASAP7_75t_L g1859 ( 
.A1(n_1845),
.A2(n_1839),
.B(n_1843),
.C(n_1841),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1847),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1851),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1854),
.B(n_1852),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1853),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1855),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1858),
.Y(n_1865)
);

INVx2_ASAP7_75t_SL g1866 ( 
.A(n_1857),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1861),
.Y(n_1867)
);

OAI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1859),
.A2(n_1856),
.B(n_1860),
.Y(n_1868)
);

AOI221x1_ASAP7_75t_L g1869 ( 
.A1(n_1868),
.A2(n_1863),
.B1(n_1864),
.B2(n_1862),
.C(n_1865),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1866),
.A2(n_1582),
.B1(n_1587),
.B2(n_1576),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1867),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1869),
.A2(n_472),
.B(n_473),
.Y(n_1872)
);

OAI322xp33_ASAP7_75t_L g1873 ( 
.A1(n_1871),
.A2(n_480),
.A3(n_478),
.B1(n_476),
.B2(n_474),
.C1(n_475),
.C2(n_477),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1870),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1872),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.C(n_484),
.Y(n_1875)
);

AOI222xp33_ASAP7_75t_L g1876 ( 
.A1(n_1873),
.A2(n_487),
.B1(n_490),
.B2(n_485),
.C1(n_486),
.C2(n_489),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1874),
.B(n_490),
.Y(n_1877)
);

NAND3xp33_ASAP7_75t_L g1878 ( 
.A(n_1877),
.B(n_1876),
.C(n_1875),
.Y(n_1878)
);

OAI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1878),
.A2(n_500),
.B(n_501),
.Y(n_1879)
);

AOI211x1_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_513),
.B(n_511),
.C(n_512),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1880),
.Y(n_1881)
);

OAI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_517),
.B1(n_515),
.B2(n_516),
.C(n_518),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1882),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1883),
.Y(n_1884)
);

INVx3_ASAP7_75t_L g1885 ( 
.A(n_1884),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_L g1886 ( 
.A(n_1885),
.B(n_520),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_L g1887 ( 
.A1(n_1886),
.A2(n_523),
.B(n_525),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_L g1888 ( 
.A(n_1887),
.B(n_526),
.C(n_527),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1888),
.Y(n_1889)
);

XOR2xp5_ASAP7_75t_L g1890 ( 
.A(n_1889),
.B(n_528),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_R g1891 ( 
.A1(n_1890),
.A2(n_531),
.B1(n_528),
.B2(n_530),
.C(n_532),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1891),
.A2(n_536),
.B(n_533),
.C(n_535),
.Y(n_1892)
);


endmodule