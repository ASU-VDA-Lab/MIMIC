module real_aes_6991_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g244 ( .A1(n_0), .A2(n_245), .B(n_246), .C(n_249), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_1), .B(n_233), .Y(n_250) );
INVx1_ASAP7_75t_L g446 ( .A(n_2), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_3), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_4), .A2(n_122), .B(n_125), .C(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_5), .A2(n_117), .B(n_573), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_6), .A2(n_117), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_7), .B(n_233), .Y(n_579) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_8), .A2(n_152), .B(n_189), .Y(n_188) );
AND2x6_ASAP7_75t_L g122 ( .A(n_9), .B(n_123), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_10), .A2(n_122), .B(n_125), .C(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g517 ( .A(n_11), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_12), .B(n_40), .Y(n_447) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_13), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_13), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_14), .B(n_209), .Y(n_551) );
INVx1_ASAP7_75t_L g143 ( .A(n_15), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_16), .B(n_161), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_17), .A2(n_162), .B(n_535), .C(n_537), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_18), .B(n_233), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_19), .B(n_137), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_20), .A2(n_125), .B(n_128), .C(n_136), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_21), .A2(n_197), .B(n_248), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_22), .B(n_209), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g435 ( .A1(n_23), .A2(n_56), .B1(n_436), .B2(n_437), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_23), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_24), .B(n_209), .Y(n_490) );
CKINVDCx16_ASAP7_75t_R g564 ( .A(n_25), .Y(n_564) );
INVx1_ASAP7_75t_L g489 ( .A(n_26), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_27), .A2(n_125), .B(n_136), .C(n_192), .Y(n_191) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_29), .Y(n_547) );
INVx1_ASAP7_75t_L g505 ( .A(n_30), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_31), .A2(n_117), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g120 ( .A(n_32), .Y(n_120) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_33), .A2(n_165), .B(n_174), .C(n_176), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_34), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_35), .A2(n_248), .B(n_576), .C(n_578), .Y(n_575) );
INVxp67_ASAP7_75t_L g506 ( .A(n_36), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_37), .B(n_194), .Y(n_193) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_38), .A2(n_125), .B(n_136), .C(n_488), .Y(n_487) );
CKINVDCx14_ASAP7_75t_R g574 ( .A(n_39), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_L g514 ( .A1(n_41), .A2(n_249), .B(n_515), .C(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_42), .B(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_43), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_44), .B(n_161), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_45), .B(n_117), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_46), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_47), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_48), .A2(n_165), .B(n_174), .C(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_49), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g247 ( .A(n_50), .Y(n_247) );
OAI22xp5_ASAP7_75t_SL g433 ( .A1(n_51), .A2(n_434), .B1(n_435), .B2(n_438), .Y(n_433) );
CKINVDCx16_ASAP7_75t_R g438 ( .A(n_51), .Y(n_438) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_52), .A2(n_462), .B1(n_463), .B2(n_472), .C1(n_752), .C2(n_756), .Y(n_461) );
INVx1_ASAP7_75t_L g219 ( .A(n_53), .Y(n_219) );
INVx1_ASAP7_75t_L g523 ( .A(n_54), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_55), .B(n_117), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_56), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_57), .Y(n_145) );
CKINVDCx14_ASAP7_75t_R g513 ( .A(n_58), .Y(n_513) );
INVx1_ASAP7_75t_L g123 ( .A(n_59), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_60), .B(n_117), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_61), .B(n_233), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_62), .A2(n_135), .B(n_158), .C(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g142 ( .A(n_63), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_64), .A2(n_102), .B1(n_468), .B2(n_469), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g469 ( .A(n_64), .Y(n_469) );
INVx1_ASAP7_75t_SL g577 ( .A(n_65), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_66), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_67), .B(n_161), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_68), .B(n_233), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_69), .B(n_162), .Y(n_207) );
INVx1_ASAP7_75t_L g567 ( .A(n_70), .Y(n_567) );
CKINVDCx16_ASAP7_75t_R g243 ( .A(n_71), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_72), .B(n_130), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_73), .A2(n_125), .B(n_156), .C(n_165), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_74), .Y(n_228) );
INVx1_ASAP7_75t_L g459 ( .A(n_75), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_76), .A2(n_117), .B(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_77), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_78), .A2(n_117), .B(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_79), .A2(n_116), .B(n_501), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_80), .Y(n_486) );
INVx1_ASAP7_75t_L g533 ( .A(n_81), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_82), .B(n_133), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_83), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_84), .A2(n_117), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g536 ( .A(n_85), .Y(n_536) );
INVx2_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
INVx1_ASAP7_75t_L g550 ( .A(n_87), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_88), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_89), .B(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g443 ( .A(n_90), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g475 ( .A(n_90), .B(n_445), .Y(n_475) );
INVx2_ASAP7_75t_L g477 ( .A(n_90), .Y(n_477) );
OAI22xp5_ASAP7_75t_SL g466 ( .A1(n_91), .A2(n_467), .B1(n_470), .B2(n_471), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_91), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_92), .A2(n_125), .B(n_165), .C(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_93), .B(n_117), .Y(n_172) );
INVx1_ASAP7_75t_L g177 ( .A(n_94), .Y(n_177) );
INVxp67_ASAP7_75t_L g231 ( .A(n_95), .Y(n_231) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_96), .A2(n_104), .B1(n_451), .B2(n_460), .C1(n_759), .C2(n_764), .Y(n_103) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_96), .B(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_96), .B(n_152), .Y(n_518) );
INVx1_ASAP7_75t_L g157 ( .A(n_97), .Y(n_157) );
INVx1_ASAP7_75t_L g203 ( .A(n_98), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_99), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g526 ( .A(n_100), .Y(n_526) );
AND2x2_ASAP7_75t_L g221 ( .A(n_101), .B(n_139), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_102), .Y(n_468) );
OAI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_440), .B(n_448), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g106 ( .A1(n_107), .A2(n_432), .B1(n_433), .B2(n_439), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_107), .A2(n_479), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g439 ( .A(n_108), .Y(n_439) );
AND3x1_ASAP7_75t_L g108 ( .A(n_109), .B(n_336), .C(n_393), .Y(n_108) );
NOR3xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_281), .C(n_317), .Y(n_109) );
OAI211xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_183), .B(n_235), .C(n_268), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_147), .Y(n_111) );
HB1xp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g238 ( .A(n_113), .B(n_239), .Y(n_238) );
INVx5_ASAP7_75t_L g267 ( .A(n_113), .Y(n_267) );
AND2x2_ASAP7_75t_L g340 ( .A(n_113), .B(n_256), .Y(n_340) );
AND2x2_ASAP7_75t_L g378 ( .A(n_113), .B(n_284), .Y(n_378) );
AND2x2_ASAP7_75t_L g398 ( .A(n_113), .B(n_240), .Y(n_398) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_144), .Y(n_113) );
AOI21xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_124), .B(n_137), .Y(n_114) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_118), .B(n_122), .Y(n_204) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_L g135 ( .A(n_119), .Y(n_135) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
INVx1_ASAP7_75t_L g198 ( .A(n_120), .Y(n_198) );
INVx1_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
INVx3_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
INVx1_ASAP7_75t_L g194 ( .A(n_121), .Y(n_194) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_121), .Y(n_209) );
BUFx3_ASAP7_75t_L g136 ( .A(n_122), .Y(n_136) );
INVx4_ASAP7_75t_SL g166 ( .A(n_122), .Y(n_166) );
INVx5_ASAP7_75t_L g175 ( .A(n_125), .Y(n_175) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
BUFx3_ASAP7_75t_L g180 ( .A(n_126), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B(n_134), .Y(n_128) );
INVx2_ASAP7_75t_L g133 ( .A(n_130), .Y(n_133) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx4_ASAP7_75t_L g159 ( .A(n_131), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_133), .A2(n_177), .B(n_178), .C(n_179), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g218 ( .A1(n_133), .A2(n_179), .B(n_219), .C(n_220), .Y(n_218) );
O2A1O1Ixp5_ASAP7_75t_L g549 ( .A1(n_133), .A2(n_550), .B(n_551), .C(n_552), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_133), .A2(n_552), .B(n_567), .C(n_568), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_134), .A2(n_161), .B(n_489), .C(n_490), .Y(n_488) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_135), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_138), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g146 ( .A(n_139), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_139), .A2(n_172), .B(n_173), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_139), .A2(n_216), .B(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_139), .A2(n_204), .B(n_486), .C(n_487), .Y(n_485) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_139), .A2(n_511), .B(n_518), .Y(n_510) );
AND2x2_ASAP7_75t_SL g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_L g153 ( .A(n_140), .B(n_141), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_146), .A2(n_546), .B(n_553), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_147), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_170), .Y(n_147) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_148), .Y(n_279) );
AND2x2_ASAP7_75t_L g293 ( .A(n_148), .B(n_239), .Y(n_293) );
INVx1_ASAP7_75t_L g316 ( .A(n_148), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_148), .B(n_267), .Y(n_355) );
OR2x2_ASAP7_75t_L g392 ( .A(n_148), .B(n_237), .Y(n_392) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_149), .Y(n_328) );
AND2x2_ASAP7_75t_L g335 ( .A(n_149), .B(n_240), .Y(n_335) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g256 ( .A(n_150), .B(n_240), .Y(n_256) );
BUFx2_ASAP7_75t_L g284 ( .A(n_150), .Y(n_284) );
AO21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_168), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_151), .B(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_151), .B(n_182), .Y(n_181) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_151), .A2(n_202), .B(n_210), .Y(n_201) );
INVx3_ASAP7_75t_L g233 ( .A(n_151), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_151), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_151), .B(n_554), .Y(n_553) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_151), .A2(n_563), .B(n_569), .Y(n_562) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_152), .A2(n_190), .B(n_191), .Y(n_189) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g212 ( .A(n_153), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_167), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B(n_160), .C(n_163), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp33_ASAP7_75t_L g504 ( .A1(n_159), .A2(n_161), .B1(n_505), .B2(n_506), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_159), .B(n_526), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_159), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_161), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g245 ( .A(n_161), .Y(n_245) );
INVx5_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_162), .B(n_517), .Y(n_516) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g578 ( .A(n_164), .Y(n_578) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_166), .A2(n_175), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_SL g242 ( .A1(n_166), .A2(n_175), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g501 ( .A1(n_166), .A2(n_175), .B(n_502), .C(n_503), .Y(n_501) );
O2A1O1Ixp33_ASAP7_75t_SL g512 ( .A1(n_166), .A2(n_175), .B(n_513), .C(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_166), .A2(n_175), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_166), .A2(n_175), .B(n_533), .C(n_534), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_L g573 ( .A1(n_166), .A2(n_175), .B(n_574), .C(n_575), .Y(n_573) );
INVx5_ASAP7_75t_L g237 ( .A(n_170), .Y(n_237) );
BUFx2_ASAP7_75t_L g260 ( .A(n_170), .Y(n_260) );
AND2x2_ASAP7_75t_L g417 ( .A(n_170), .B(n_271), .Y(n_417) );
OR2x6_ASAP7_75t_L g170 ( .A(n_171), .B(n_181), .Y(n_170) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g249 ( .A(n_180), .Y(n_249) );
INVx1_ASAP7_75t_L g537 ( .A(n_180), .Y(n_537) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NAND2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_222), .Y(n_184) );
OAI221xp5_ASAP7_75t_L g317 ( .A1(n_185), .A2(n_318), .B1(n_325), .B2(n_326), .C(n_329), .Y(n_317) );
OR2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_199), .Y(n_185) );
AND2x2_ASAP7_75t_L g223 ( .A(n_186), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_186), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g252 ( .A(n_187), .B(n_200), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_187), .B(n_201), .Y(n_262) );
OR2x2_ASAP7_75t_L g273 ( .A(n_187), .B(n_224), .Y(n_273) );
AND2x2_ASAP7_75t_L g276 ( .A(n_187), .B(n_264), .Y(n_276) );
AND2x2_ASAP7_75t_L g292 ( .A(n_187), .B(n_213), .Y(n_292) );
OR2x2_ASAP7_75t_L g308 ( .A(n_187), .B(n_201), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_187), .B(n_224), .Y(n_370) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_188), .B(n_213), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_188), .B(n_201), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_195), .B(n_196), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_196), .A2(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
OR2x2_ASAP7_75t_L g286 ( .A(n_199), .B(n_273), .Y(n_286) );
INVx2_ASAP7_75t_L g312 ( .A(n_199), .Y(n_312) );
OR2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
AND2x2_ASAP7_75t_L g234 ( .A(n_200), .B(n_214), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_200), .B(n_224), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_200), .B(n_214), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_200), .B(n_264), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_200), .A2(n_395), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_394) );
INVx5_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_201), .B(n_224), .Y(n_333) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_204), .A2(n_547), .B(n_548), .Y(n_546) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_204), .A2(n_564), .B(n_565), .Y(n_563) );
INVx4_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
INVx2_ASAP7_75t_L g515 ( .A(n_209), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx2_ASAP7_75t_L g498 ( .A(n_212), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_213), .B(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_213), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g280 ( .A(n_213), .B(n_252), .Y(n_280) );
OR2x2_ASAP7_75t_L g324 ( .A(n_213), .B(n_224), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_213), .B(n_276), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_213), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g389 ( .A(n_213), .B(n_390), .Y(n_389) );
INVx5_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_SL g253 ( .A(n_214), .B(n_223), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_214), .A2(n_258), .B(n_261), .C(n_265), .Y(n_257) );
OR2x2_ASAP7_75t_L g295 ( .A(n_214), .B(n_291), .Y(n_295) );
OR2x2_ASAP7_75t_L g331 ( .A(n_214), .B(n_273), .Y(n_331) );
OAI311xp33_ASAP7_75t_L g337 ( .A1(n_214), .A2(n_276), .A3(n_338), .B1(n_341), .C1(n_348), .Y(n_337) );
AND2x2_ASAP7_75t_L g388 ( .A(n_214), .B(n_224), .Y(n_388) );
AND2x2_ASAP7_75t_L g396 ( .A(n_214), .B(n_251), .Y(n_396) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_214), .Y(n_414) );
AND2x2_ASAP7_75t_L g431 ( .A(n_214), .B(n_252), .Y(n_431) );
OR2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_221), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
AND2x2_ASAP7_75t_L g259 ( .A(n_223), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g415 ( .A(n_223), .Y(n_415) );
AND2x2_ASAP7_75t_L g251 ( .A(n_224), .B(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g264 ( .A(n_224), .Y(n_264) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_224), .Y(n_307) );
INVxp67_ASAP7_75t_L g346 ( .A(n_224), .Y(n_346) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
OA21x2_ASAP7_75t_L g520 ( .A1(n_225), .A2(n_521), .B(n_527), .Y(n_520) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_225), .A2(n_531), .B(n_538), .Y(n_530) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_225), .A2(n_572), .B(n_579), .Y(n_571) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_233), .A2(n_241), .B(n_250), .Y(n_240) );
AND2x2_ASAP7_75t_L g424 ( .A(n_234), .B(n_272), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_251), .B1(n_253), .B2(n_254), .C(n_257), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_237), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g277 ( .A(n_237), .B(n_267), .Y(n_277) );
AND2x2_ASAP7_75t_L g285 ( .A(n_237), .B(n_239), .Y(n_285) );
OR2x2_ASAP7_75t_L g297 ( .A(n_237), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g315 ( .A(n_237), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g339 ( .A(n_237), .B(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_237), .Y(n_359) );
AND2x2_ASAP7_75t_L g411 ( .A(n_237), .B(n_335), .Y(n_411) );
OAI31xp33_ASAP7_75t_L g419 ( .A1(n_237), .A2(n_288), .A3(n_387), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_238), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_SL g383 ( .A(n_238), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_238), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g271 ( .A(n_239), .B(n_267), .Y(n_271) );
INVx1_ASAP7_75t_L g358 ( .A(n_239), .Y(n_358) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g408 ( .A(n_240), .B(n_267), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_248), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g552 ( .A(n_249), .Y(n_552) );
INVx1_ASAP7_75t_SL g418 ( .A(n_251), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_252), .B(n_323), .Y(n_322) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_253), .A2(n_365), .B1(n_403), .B2(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g266 ( .A(n_256), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g325 ( .A(n_256), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_256), .B(n_277), .Y(n_430) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g400 ( .A(n_259), .B(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_260), .A2(n_319), .B(n_321), .Y(n_318) );
OR2x2_ASAP7_75t_L g326 ( .A(n_260), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g347 ( .A(n_260), .B(n_335), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_260), .B(n_358), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_260), .B(n_398), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g374 ( .A1(n_261), .A2(n_375), .B1(n_380), .B2(n_383), .C(n_384), .Y(n_374) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
OR2x2_ASAP7_75t_L g351 ( .A(n_262), .B(n_324), .Y(n_351) );
INVx1_ASAP7_75t_L g390 ( .A(n_262), .Y(n_390) );
INVx2_ASAP7_75t_L g366 ( .A(n_263), .Y(n_366) );
INVx1_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
INVx1_ASAP7_75t_SL g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g305 ( .A(n_267), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_267), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g334 ( .A(n_267), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g422 ( .A(n_267), .B(n_392), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B1(n_274), .B2(n_277), .C1(n_278), .C2(n_280), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_271), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_271), .A2(n_321), .B1(n_349), .B2(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_271), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_SL g275 ( .A(n_276), .Y(n_275) );
OAI21xp33_ASAP7_75t_SL g309 ( .A1(n_280), .A2(n_310), .B(n_313), .Y(n_309) );
OAI211xp5_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_286), .B(n_287), .C(n_309), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AOI221xp5_ASAP7_75t_L g287 ( .A1(n_285), .A2(n_288), .B1(n_293), .B2(n_294), .C(n_296), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_285), .B(n_373), .Y(n_372) );
INVxp67_ASAP7_75t_L g379 ( .A(n_285), .Y(n_379) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AND2x2_ASAP7_75t_L g381 ( .A(n_290), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g298 ( .A(n_293), .Y(n_298) );
AND2x2_ASAP7_75t_L g304 ( .A(n_293), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .B1(n_303), .B2(n_306), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_300), .B(n_312), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_301), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g401 ( .A(n_305), .Y(n_401) );
AND2x2_ASAP7_75t_L g420 ( .A(n_305), .B(n_335), .Y(n_420) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_312), .B(n_369), .Y(n_428) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_315), .B(n_383), .Y(n_426) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g349 ( .A(n_327), .Y(n_349) );
BUFx2_ASAP7_75t_L g373 ( .A(n_328), .Y(n_373) );
OAI21xp5_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_332), .B(n_334), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_352), .C(n_374), .Y(n_336) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_356), .B(n_360), .C(n_363), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_353), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NOR2xp67_ASAP7_75t_SL g357 ( .A(n_358), .B(n_359), .Y(n_357) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_SL g382 ( .A(n_362), .Y(n_382) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B(n_371), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g387 ( .A(n_365), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B1(n_389), .B2(n_391), .Y(n_384) );
INVx2_ASAP7_75t_SL g405 ( .A(n_392), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_409), .C(n_421), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_405), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_412), .B1(n_416), .B2(n_418), .C(n_419), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g421 ( .A1(n_410), .A2(n_422), .B(n_423), .C(n_425), .Y(n_421) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_427), .B1(n_429), .B2(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_439), .A2(n_473), .B1(n_476), .B2(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_443), .Y(n_450) );
INVx1_ASAP7_75t_SL g763 ( .A(n_443), .Y(n_763) );
BUFx2_ASAP7_75t_L g766 ( .A(n_443), .Y(n_766) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_444), .B(n_477), .Y(n_758) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g476 ( .A(n_445), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
CKINVDCx6p67_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_SL g761 ( .A(n_456), .B(n_458), .Y(n_761) );
OA21x2_ASAP7_75t_L g765 ( .A1(n_456), .A2(n_457), .B(n_766), .Y(n_765) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVxp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g470 ( .A(n_467), .Y(n_470) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g753 ( .A(n_474), .Y(n_753) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g755 ( .A(n_476), .Y(n_755) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OR5x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_646), .C(n_710), .D(n_726), .E(n_741), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_481), .B(n_580), .C(n_607), .D(n_630), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_528), .B(n_539), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_493), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_SL g559 ( .A(n_484), .Y(n_559) );
AND2x4_ASAP7_75t_L g593 ( .A(n_484), .B(n_582), .Y(n_593) );
OR2x2_ASAP7_75t_L g603 ( .A(n_484), .B(n_561), .Y(n_603) );
OR2x2_ASAP7_75t_L g649 ( .A(n_484), .B(n_496), .Y(n_649) );
AND2x2_ASAP7_75t_L g663 ( .A(n_484), .B(n_560), .Y(n_663) );
AND2x2_ASAP7_75t_L g706 ( .A(n_484), .B(n_596), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_484), .B(n_571), .Y(n_713) );
AND2x2_ASAP7_75t_L g732 ( .A(n_484), .B(n_622), .Y(n_732) );
AND2x2_ASAP7_75t_L g750 ( .A(n_484), .B(n_592), .Y(n_750) );
OR2x6_ASAP7_75t_L g484 ( .A(n_485), .B(n_491), .Y(n_484) );
INVx1_ASAP7_75t_L g715 ( .A(n_493), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_509), .Y(n_493) );
AND2x2_ASAP7_75t_L g625 ( .A(n_494), .B(n_560), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_494), .B(n_645), .Y(n_644) );
AOI32xp33_ASAP7_75t_L g658 ( .A1(n_494), .A2(n_659), .A3(n_662), .B1(n_664), .B2(n_668), .Y(n_658) );
AND2x2_ASAP7_75t_L g728 ( .A(n_494), .B(n_622), .Y(n_728) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g592 ( .A(n_496), .B(n_561), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_496), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g634 ( .A(n_496), .B(n_581), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_496), .B(n_713), .Y(n_712) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_499), .B(n_507), .Y(n_496) );
INVx1_ASAP7_75t_L g597 ( .A(n_497), .Y(n_597) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OA21x2_ASAP7_75t_L g596 ( .A1(n_500), .A2(n_508), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g599 ( .A(n_509), .B(n_543), .Y(n_599) );
AND2x2_ASAP7_75t_L g675 ( .A(n_509), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g747 ( .A(n_509), .Y(n_747) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
OR2x2_ASAP7_75t_L g542 ( .A(n_510), .B(n_520), .Y(n_542) );
AND2x2_ASAP7_75t_L g556 ( .A(n_510), .B(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_510), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g606 ( .A(n_510), .Y(n_606) );
AND2x2_ASAP7_75t_L g633 ( .A(n_510), .B(n_520), .Y(n_633) );
BUFx3_ASAP7_75t_L g636 ( .A(n_510), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_510), .B(n_611), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_510), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g587 ( .A(n_519), .Y(n_587) );
AND2x2_ASAP7_75t_L g605 ( .A(n_519), .B(n_585), .Y(n_605) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x2_ASAP7_75t_L g616 ( .A(n_520), .B(n_530), .Y(n_616) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_520), .Y(n_629) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_529), .B(n_636), .Y(n_686) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_SL g557 ( .A(n_530), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_530), .B(n_605), .C(n_606), .Y(n_604) );
OR2x2_ASAP7_75t_L g612 ( .A(n_530), .B(n_585), .Y(n_612) );
AND2x2_ASAP7_75t_L g632 ( .A(n_530), .B(n_585), .Y(n_632) );
AND2x2_ASAP7_75t_L g676 ( .A(n_530), .B(n_545), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_555), .B(n_558), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x2_ASAP7_75t_L g751 ( .A(n_541), .B(n_676), .Y(n_751) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_542), .A2(n_649), .B1(n_691), .B2(n_693), .Y(n_690) );
OR2x2_ASAP7_75t_L g697 ( .A(n_542), .B(n_612), .Y(n_697) );
OR2x2_ASAP7_75t_L g721 ( .A(n_542), .B(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_542), .B(n_641), .Y(n_734) );
AND2x2_ASAP7_75t_L g627 ( .A(n_543), .B(n_628), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_543), .A2(n_700), .B(n_715), .Y(n_714) );
AOI32xp33_ASAP7_75t_L g735 ( .A1(n_543), .A2(n_625), .A3(n_736), .B1(n_738), .B2(n_739), .Y(n_735) );
OR2x2_ASAP7_75t_L g746 ( .A(n_543), .B(n_747), .Y(n_746) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g614 ( .A(n_544), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_544), .B(n_628), .Y(n_693) );
BUFx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g585 ( .A(n_545), .Y(n_585) );
AND2x2_ASAP7_75t_L g651 ( .A(n_545), .B(n_616), .Y(n_651) );
AND3x2_ASAP7_75t_L g660 ( .A(n_545), .B(n_556), .C(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g586 ( .A(n_557), .B(n_587), .Y(n_586) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_557), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_557), .B(n_585), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g581 ( .A(n_559), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g621 ( .A(n_559), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g639 ( .A(n_559), .B(n_571), .Y(n_639) );
AND2x2_ASAP7_75t_L g657 ( .A(n_559), .B(n_561), .Y(n_657) );
OR2x2_ASAP7_75t_L g671 ( .A(n_559), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g717 ( .A(n_559), .B(n_645), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_560), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_571), .Y(n_560) );
AND2x2_ASAP7_75t_L g618 ( .A(n_561), .B(n_596), .Y(n_618) );
OR2x2_ASAP7_75t_L g672 ( .A(n_561), .B(n_596), .Y(n_672) );
AND2x2_ASAP7_75t_L g725 ( .A(n_561), .B(n_582), .Y(n_725) );
INVx2_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g623 ( .A(n_562), .Y(n_623) );
AND2x2_ASAP7_75t_L g645 ( .A(n_562), .B(n_571), .Y(n_645) );
INVx2_ASAP7_75t_L g582 ( .A(n_571), .Y(n_582) );
INVx1_ASAP7_75t_L g602 ( .A(n_571), .Y(n_602) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .B(n_588), .C(n_600), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_581), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g744 ( .A(n_581), .Y(n_744) );
AND2x2_ASAP7_75t_L g622 ( .A(n_582), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_585), .B(n_586), .Y(n_594) );
INVx1_ASAP7_75t_L g679 ( .A(n_585), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_585), .B(n_606), .Y(n_703) );
AND2x2_ASAP7_75t_L g719 ( .A(n_585), .B(n_633), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_586), .B(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g610 ( .A(n_587), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_594), .B1(n_595), .B2(n_598), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_591), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_592), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g617 ( .A(n_593), .B(n_618), .Y(n_617) );
AOI221xp5_ASAP7_75t_SL g682 ( .A1(n_593), .A2(n_635), .B1(n_683), .B2(n_688), .C(n_690), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_593), .B(n_656), .Y(n_689) );
INVx1_ASAP7_75t_L g749 ( .A(n_595), .Y(n_749) );
BUFx3_ASAP7_75t_L g656 ( .A(n_596), .Y(n_656) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI21xp33_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_603), .B(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g665 ( .A(n_602), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_602), .B(n_656), .Y(n_709) );
INVx1_ASAP7_75t_L g666 ( .A(n_603), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_603), .B(n_656), .Y(n_667) );
INVxp67_ASAP7_75t_L g687 ( .A(n_605), .Y(n_687) );
AND2x2_ASAP7_75t_L g628 ( .A(n_606), .B(n_629), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_613), .B(n_617), .C(n_619), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
INVx1_ASAP7_75t_SL g642 ( .A(n_610), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_611), .B(n_642), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_611), .B(n_633), .Y(n_684) );
INVx2_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_614), .A2(n_620), .B1(n_624), .B2(n_626), .Y(n_619) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g635 ( .A(n_616), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g680 ( .A(n_616), .B(n_681), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_618), .A2(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_622), .A2(n_631), .B1(n_634), .B2(n_635), .C(n_637), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_622), .B(n_656), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_622), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g738 ( .A(n_628), .Y(n_738) );
INVxp67_ASAP7_75t_L g661 ( .A(n_629), .Y(n_661) );
INVx1_ASAP7_75t_L g668 ( .A(n_631), .Y(n_668) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_L g707 ( .A(n_632), .B(n_636), .Y(n_707) );
INVx1_ASAP7_75t_L g681 ( .A(n_636), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_636), .B(n_651), .Y(n_711) );
OAI32xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .A3(n_642), .B1(n_643), .B2(n_644), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_SL g650 ( .A(n_645), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_645), .B(n_677), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_645), .B(n_706), .Y(n_737) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_645), .B(n_656), .Y(n_745) );
NAND5xp2_ASAP7_75t_L g646 ( .A(n_647), .B(n_669), .C(n_682), .D(n_694), .E(n_695), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B1(n_652), .B2(n_654), .C(n_658), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND2xp33_ASAP7_75t_SL g673 ( .A(n_653), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_657), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_656), .B(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_657), .A2(n_670), .B1(n_673), .B2(n_677), .Y(n_669) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_660), .A2(n_665), .B(n_666), .C(n_667), .Y(n_664) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g692 ( .A(n_672), .Y(n_692) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_681), .B(n_730), .Y(n_740) );
OR2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI222xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_700), .B2(n_704), .C1(n_707), .C2(n_708), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_714), .B2(n_716), .C(n_718), .Y(n_710) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B(n_723), .Y(n_718) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g730 ( .A(n_722), .Y(n_730) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_729), .B1(n_731), .B2(n_733), .C(n_735), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_745), .B(n_746), .C(n_748), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI21xp33_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B(n_751), .Y(n_748) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
NAND2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
endmodule