module real_aes_6116_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_980;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_923;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_478;
wire n_356;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_976;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_931;
wire n_904;
wire n_780;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_909;
wire n_298;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_973;
wire n_960;
wire n_455;
wire n_671;
wire n_725;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_713;
wire n_288;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_749;
wire n_358;
wire n_275;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_915;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_823;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_0), .A2(n_62), .B1(n_394), .B2(n_403), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_1), .A2(n_235), .B1(n_545), .B2(n_549), .Y(n_668) );
AO22x2_ASAP7_75t_L g650 ( .A1(n_2), .A2(n_651), .B1(n_670), .B2(n_671), .Y(n_650) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_2), .Y(n_670) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_3), .Y(n_278) );
AND2x4_ASAP7_75t_L g734 ( .A(n_3), .B(n_735), .Y(n_734) );
AND2x4_ASAP7_75t_L g740 ( .A(n_3), .B(n_255), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g952 ( .A1(n_4), .A2(n_27), .B1(n_404), .B2(n_615), .Y(n_952) );
AO22x1_ASAP7_75t_L g738 ( .A1(n_5), .A2(n_7), .B1(n_739), .B2(n_741), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_6), .A2(n_121), .B1(n_457), .B2(n_459), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_8), .A2(n_185), .B1(n_731), .B2(n_746), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_9), .A2(n_200), .B1(n_403), .B2(n_404), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_10), .A2(n_227), .B1(n_397), .B2(n_399), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_11), .A2(n_175), .B1(n_404), .B2(n_472), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_12), .A2(n_96), .B1(n_545), .B2(n_549), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_13), .A2(n_17), .B1(n_334), .B2(n_336), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_14), .A2(n_45), .B1(n_527), .B2(n_560), .Y(n_953) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_15), .A2(n_19), .B1(n_387), .B2(n_389), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_16), .A2(n_206), .B1(n_387), .B2(n_462), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_18), .B(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_20), .A2(n_84), .B1(n_395), .B2(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g493 ( .A(n_21), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_22), .A2(n_132), .B1(n_549), .B2(n_550), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_23), .A2(n_125), .B1(n_489), .B2(n_511), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_24), .A2(n_195), .B1(n_509), .B2(n_677), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_25), .A2(n_122), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_26), .A2(n_127), .B1(n_409), .B2(n_447), .Y(n_961) );
INVx1_ASAP7_75t_L g607 ( .A(n_28), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_29), .A2(n_204), .B1(n_638), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_30), .A2(n_151), .B1(n_387), .B2(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g362 ( .A(n_31), .Y(n_362) );
AOI21x1_ASAP7_75t_L g486 ( .A1(n_32), .A2(n_487), .B(n_492), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_33), .A2(n_167), .B1(n_338), .B2(n_341), .Y(n_546) );
XOR2x2_ASAP7_75t_L g693 ( .A(n_34), .B(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_35), .A2(n_142), .B1(n_348), .B2(n_364), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_36), .A2(n_217), .B1(n_495), .B2(n_964), .Y(n_963) );
XNOR2x1_ASAP7_75t_L g600 ( .A(n_37), .B(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_38), .A2(n_78), .B1(n_397), .B2(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g517 ( .A(n_39), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_40), .B(n_194), .Y(n_276) );
INVx1_ASAP7_75t_L g311 ( .A(n_40), .Y(n_311) );
INVxp67_ASAP7_75t_L g358 ( .A(n_40), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_41), .A2(n_130), .B1(n_334), .B2(n_348), .Y(n_547) );
INVx1_ASAP7_75t_L g452 ( .A(n_42), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_43), .B(n_679), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_44), .A2(n_104), .B1(n_394), .B2(n_395), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_46), .A2(n_155), .B1(n_419), .B2(n_483), .Y(n_962) );
OAI22xp33_ASAP7_75t_R g970 ( .A1(n_47), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_970) );
CKINVDCx5p33_ASAP7_75t_R g972 ( .A(n_47), .Y(n_972) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_48), .A2(n_77), .B1(n_536), .B2(n_550), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_49), .B(n_295), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_50), .A2(n_119), .B1(n_444), .B2(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_51), .A2(n_89), .B1(n_478), .B2(n_562), .Y(n_561) );
AOI21xp33_ASAP7_75t_SL g653 ( .A1(n_52), .A2(n_654), .B(n_655), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_53), .A2(n_241), .B1(n_462), .B2(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_54), .A2(n_181), .B1(n_289), .B2(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g634 ( .A(n_55), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_56), .A2(n_246), .B1(n_364), .B2(n_538), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_57), .A2(n_216), .B1(n_361), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_58), .A2(n_168), .B1(n_445), .B2(n_572), .Y(n_571) );
BUFx2_ASAP7_75t_L g660 ( .A(n_59), .Y(n_660) );
XNOR2x1_ASAP7_75t_L g440 ( .A(n_60), .B(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_61), .A2(n_103), .B1(n_334), .B2(n_336), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_63), .A2(n_163), .B1(n_741), .B2(n_757), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_64), .A2(n_190), .B1(n_334), .B2(n_336), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_65), .A2(n_252), .B1(n_289), .B2(n_314), .Y(n_288) );
INVx2_ASAP7_75t_L g273 ( .A(n_66), .Y(n_273) );
INVx1_ASAP7_75t_L g702 ( .A(n_67), .Y(n_702) );
INVx1_ASAP7_75t_L g733 ( .A(n_68), .Y(n_733) );
AND2x4_ASAP7_75t_L g737 ( .A(n_68), .B(n_273), .Y(n_737) );
INVx1_ASAP7_75t_SL g745 ( .A(n_68), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_69), .A2(n_199), .B1(n_338), .B2(n_341), .Y(n_337) );
INVx1_ASAP7_75t_L g704 ( .A(n_70), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_71), .A2(n_154), .B1(n_445), .B2(n_511), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_72), .A2(n_179), .B1(n_457), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_73), .A2(n_231), .B1(n_711), .B2(n_713), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_74), .B(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_75), .A2(n_165), .B1(n_409), .B2(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_76), .A2(n_160), .B1(n_314), .B2(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_79), .A2(n_173), .B1(n_739), .B2(n_758), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_80), .A2(n_224), .B1(n_394), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g402 ( .A1(n_81), .A2(n_239), .B1(n_403), .B2(n_404), .Y(n_402) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_82), .Y(n_295) );
XNOR2x2_ASAP7_75t_SL g285 ( .A(n_83), .B(n_286), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_85), .A2(n_196), .B1(n_338), .B2(n_341), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_86), .A2(n_262), .B1(n_336), .B2(n_545), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_87), .A2(n_176), .B1(n_476), .B2(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g625 ( .A(n_88), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_90), .A2(n_513), .B(n_516), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_91), .A2(n_157), .B1(n_731), .B2(n_736), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_92), .A2(n_93), .B1(n_364), .B2(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_94), .A2(n_210), .B1(n_416), .B2(n_419), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_95), .A2(n_150), .B1(n_507), .B2(n_509), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_97), .A2(n_184), .B1(n_741), .B2(n_757), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_98), .A2(n_266), .B1(n_409), .B2(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g296 ( .A(n_99), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_99), .B(n_193), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_100), .A2(n_170), .B1(n_739), .B2(n_741), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_101), .A2(n_247), .B1(n_314), .B2(n_464), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_102), .A2(n_166), .B1(n_447), .B2(n_448), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_105), .A2(n_162), .B1(n_731), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_106), .A2(n_207), .B1(n_348), .B2(n_361), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_107), .A2(n_152), .B1(n_445), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_108), .A2(n_113), .B1(n_731), .B2(n_746), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_109), .A2(n_232), .B1(n_367), .B2(n_369), .C(n_371), .Y(n_366) );
XNOR2x1_ASAP7_75t_L g531 ( .A(n_110), .B(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_111), .A2(n_174), .B1(n_427), .B2(n_430), .Y(n_426) );
INVx1_ASAP7_75t_L g719 ( .A(n_112), .Y(n_719) );
INVx1_ASAP7_75t_L g383 ( .A(n_114), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_115), .A2(n_202), .B1(n_399), .B2(n_404), .Y(n_523) );
INVx1_ASAP7_75t_L g707 ( .A(n_116), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_117), .A2(n_153), .B1(n_397), .B2(n_399), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_118), .A2(n_197), .B1(n_754), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_120), .A2(n_261), .B1(n_536), .B2(n_550), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_123), .A2(n_221), .B1(n_564), .B2(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_124), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g372 ( .A(n_126), .Y(n_372) );
INVx1_ASAP7_75t_L g656 ( .A(n_128), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_129), .A2(n_245), .B1(n_731), .B2(n_746), .Y(n_773) );
AOI21xp33_ASAP7_75t_L g539 ( .A1(n_131), .A2(n_370), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_133), .Y(n_541) );
INVx1_ASAP7_75t_L g609 ( .A(n_134), .Y(n_609) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_135), .B(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_136), .A2(n_225), .B1(n_364), .B2(n_444), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g449 ( .A1(n_137), .A2(n_450), .B(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_138), .A2(n_147), .B1(n_325), .B2(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_139), .A2(n_409), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g346 ( .A(n_140), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_141), .A2(n_198), .B1(n_461), .B2(n_462), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_143), .A2(n_145), .B1(n_314), .B2(n_527), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_144), .A2(n_226), .B1(n_399), .B2(n_697), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_146), .A2(n_244), .B1(n_744), .B2(n_746), .Y(n_743) );
INVx1_ASAP7_75t_L g673 ( .A(n_148), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_149), .B(n_491), .Y(n_534) );
INVx1_ASAP7_75t_L g706 ( .A(n_156), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_158), .B(n_498), .Y(n_573) );
INVx1_ASAP7_75t_L g577 ( .A(n_159), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_159), .A2(n_211), .B1(n_749), .B2(n_757), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_161), .A2(n_209), .B1(n_289), .B2(n_615), .Y(n_614) );
XOR2xp5_ASAP7_75t_L g503 ( .A(n_164), .B(n_504), .Y(n_503) );
AO221x2_ASAP7_75t_L g730 ( .A1(n_169), .A2(n_220), .B1(n_731), .B2(n_736), .C(n_738), .Y(n_730) );
OA22x2_ASAP7_75t_L g301 ( .A1(n_171), .A2(n_194), .B1(n_295), .B2(n_299), .Y(n_301) );
INVx1_ASAP7_75t_L g321 ( .A(n_171), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_172), .A2(n_264), .B1(n_404), .B2(n_620), .Y(n_619) );
XOR2x2_ASAP7_75t_L g555 ( .A(n_173), .B(n_556), .Y(n_555) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_177), .A2(n_180), .B1(n_338), .B2(n_341), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_178), .A2(n_249), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI222xp33_ASAP7_75t_L g948 ( .A1(n_178), .A2(n_949), .B1(n_966), .B2(n_970), .C1(n_974), .C2(n_976), .Y(n_948) );
INVx1_ASAP7_75t_SL g965 ( .A(n_178), .Y(n_965) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_182), .A2(n_251), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_183), .A2(n_243), .B1(n_545), .B2(n_549), .Y(n_636) );
XOR2x2_ASAP7_75t_L g468 ( .A(n_186), .B(n_469), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_187), .A2(n_215), .B1(n_361), .B2(n_538), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_188), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_189), .B(n_514), .Y(n_580) );
BUFx2_ASAP7_75t_L g662 ( .A(n_191), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_192), .A2(n_222), .B1(n_338), .B2(n_341), .Y(n_669) );
INVx1_ASAP7_75t_L g313 ( .A(n_193), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_193), .B(n_319), .Y(n_378) );
OAI21xp33_ASAP7_75t_L g322 ( .A1(n_194), .A2(n_213), .B(n_323), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_201), .A2(n_223), .B1(n_325), .B2(n_329), .Y(n_324) );
INVx1_ASAP7_75t_L g605 ( .A(n_203), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_205), .A2(n_242), .B1(n_536), .B2(n_550), .Y(n_587) );
INVx1_ASAP7_75t_L g412 ( .A(n_208), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_212), .A2(n_260), .B1(n_369), .B2(n_423), .C(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_213), .B(n_248), .Y(n_277) );
INVx1_ASAP7_75t_L g298 ( .A(n_213), .Y(n_298) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_214), .A2(n_409), .B(n_411), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_218), .A2(n_229), .B1(n_612), .B2(n_627), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_219), .A2(n_250), .B1(n_483), .B2(n_622), .C(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g684 ( .A(n_228), .Y(n_684) );
INVx1_ASAP7_75t_L g585 ( .A(n_230), .Y(n_585) );
AOI21xp33_ASAP7_75t_L g583 ( .A1(n_233), .A2(n_370), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_234), .A2(n_238), .B1(n_397), .B2(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_236), .A2(n_256), .B1(n_403), .B2(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_237), .A2(n_491), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_240), .B(n_960), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_248), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g496 ( .A(n_253), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_254), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g735 ( .A(n_255), .Y(n_735) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_255), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_257), .A2(n_258), .B1(n_461), .B2(n_462), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_259), .A2(n_263), .B1(n_387), .B2(n_462), .Y(n_618) );
INVx1_ASAP7_75t_L g365 ( .A(n_265), .Y(n_365) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_279), .B(n_724), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx4_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_274), .C(n_278), .Y(n_270) );
AND2x2_ASAP7_75t_L g967 ( .A(n_271), .B(n_968), .Y(n_967) );
AND2x2_ASAP7_75t_L g975 ( .A(n_271), .B(n_969), .Y(n_975) );
AOI21xp5_ASAP7_75t_L g980 ( .A1(n_271), .A2(n_278), .B(n_745), .Y(n_980) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AO21x1_ASAP7_75t_L g977 ( .A1(n_272), .A2(n_978), .B(n_980), .Y(n_977) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g732 ( .A(n_273), .B(n_733), .Y(n_732) );
AND3x4_ASAP7_75t_L g744 ( .A(n_273), .B(n_734), .C(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_274), .B(n_969), .Y(n_968) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AO21x2_ASAP7_75t_L g375 ( .A1(n_275), .A2(n_376), .B(n_377), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g969 ( .A(n_278), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B1(n_595), .B2(n_597), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
XNOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_500), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B1(n_436), .B2(n_499), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AO22x2_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_379), .B1(n_434), .B2(n_435), .Y(n_284) );
INVx2_ASAP7_75t_L g434 ( .A(n_285), .Y(n_434) );
NAND4xp75_ASAP7_75t_L g286 ( .A(n_287), .B(n_332), .C(n_344), .D(n_366), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_324), .Y(n_287) );
BUFx12f_ASAP7_75t_L g562 ( .A(n_289), .Y(n_562) );
INVx1_ASAP7_75t_L g712 ( .A(n_289), .Y(n_712) );
BUFx12f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_290), .Y(n_394) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_290), .Y(n_464) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_302), .Y(n_290) );
AND2x4_ASAP7_75t_L g326 ( .A(n_291), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g338 ( .A(n_291), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g341 ( .A(n_291), .B(n_342), .Y(n_341) );
AND2x4_ASAP7_75t_L g388 ( .A(n_291), .B(n_339), .Y(n_388) );
AND2x2_ASAP7_75t_L g392 ( .A(n_291), .B(n_342), .Y(n_392) );
AND2x4_ASAP7_75t_L g536 ( .A(n_291), .B(n_401), .Y(n_536) );
AND2x4_ASAP7_75t_L g545 ( .A(n_291), .B(n_302), .Y(n_545) );
AND2x4_ASAP7_75t_L g291 ( .A(n_292), .B(n_300), .Y(n_291) );
AND2x2_ASAP7_75t_L g349 ( .A(n_292), .B(n_301), .Y(n_349) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g335 ( .A(n_293), .B(n_301), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
NAND2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
INVx2_ASAP7_75t_L g299 ( .A(n_295), .Y(n_299) );
INVx3_ASAP7_75t_L g305 ( .A(n_295), .Y(n_305) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_295), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g323 ( .A(n_295), .Y(n_323) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_295), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_296), .B(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_298), .A2(n_323), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g356 ( .A(n_301), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g316 ( .A(n_302), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g334 ( .A(n_302), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g398 ( .A(n_302), .B(n_335), .Y(n_398) );
AND2x2_ASAP7_75t_L g458 ( .A(n_302), .B(n_335), .Y(n_458) );
AND2x4_ASAP7_75t_L g549 ( .A(n_302), .B(n_317), .Y(n_549) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_307), .Y(n_302) );
OR2x2_ASAP7_75t_L g328 ( .A(n_303), .B(n_308), .Y(n_328) );
AND2x4_ASAP7_75t_L g339 ( .A(n_303), .B(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
AND2x2_ASAP7_75t_L g352 ( .A(n_303), .B(n_353), .Y(n_352) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_305), .B(n_311), .Y(n_310) );
INVxp67_ASAP7_75t_L g319 ( .A(n_305), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g377 ( .A(n_306), .B(n_318), .C(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
AND2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx4_ASAP7_75t_L g395 ( .A(n_315), .Y(n_395) );
INVx1_ASAP7_75t_L g478 ( .A(n_315), .Y(n_478) );
INVx1_ASAP7_75t_L g699 ( .A(n_315), .Y(n_699) );
INVx2_ASAP7_75t_L g957 ( .A(n_315), .Y(n_957) );
INVx8_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g331 ( .A(n_317), .B(n_327), .Y(n_331) );
AND2x4_ASAP7_75t_L g364 ( .A(n_317), .B(n_342), .Y(n_364) );
AND2x4_ASAP7_75t_L g420 ( .A(n_317), .B(n_342), .Y(n_420) );
AND2x4_ASAP7_75t_L g550 ( .A(n_317), .B(n_327), .Y(n_550) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_322), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
BUFx3_ASAP7_75t_L g713 ( .A(n_325), .Y(n_713) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_326), .Y(n_403) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_326), .Y(n_472) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_326), .Y(n_615) );
AND2x4_ASAP7_75t_L g336 ( .A(n_327), .B(n_335), .Y(n_336) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g401 ( .A(n_328), .Y(n_401) );
INVx3_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx5_ASAP7_75t_L g466 ( .A(n_330), .Y(n_466) );
INVx2_ASAP7_75t_L g687 ( .A(n_330), .Y(n_687) );
INVx6_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx12f_ASAP7_75t_L g404 ( .A(n_331), .Y(n_404) );
AND2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .Y(n_332) );
AND2x4_ASAP7_75t_L g361 ( .A(n_335), .B(n_339), .Y(n_361) );
AND2x2_ASAP7_75t_L g368 ( .A(n_335), .B(n_342), .Y(n_368) );
AND2x4_ASAP7_75t_L g400 ( .A(n_335), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g425 ( .A(n_335), .B(n_342), .Y(n_425) );
AND2x2_ASAP7_75t_L g433 ( .A(n_335), .B(n_339), .Y(n_433) );
AND2x4_ASAP7_75t_L g348 ( .A(n_339), .B(n_349), .Y(n_348) );
AND2x4_ASAP7_75t_L g410 ( .A(n_339), .B(n_349), .Y(n_410) );
AND2x4_ASAP7_75t_L g342 ( .A(n_340), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g370 ( .A(n_342), .B(n_349), .Y(n_370) );
AND2x4_ASAP7_75t_L g418 ( .A(n_342), .B(n_349), .Y(n_418) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_359), .Y(n_344) );
OAI21xp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B(n_350), .Y(n_345) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g518 ( .A(n_351), .Y(n_518) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_356), .Y(n_351) );
AND2x4_ASAP7_75t_L g429 ( .A(n_352), .B(n_356), .Y(n_429) );
AND2x2_ASAP7_75t_L g538 ( .A(n_352), .B(n_356), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g376 ( .A(n_354), .Y(n_376) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B1(n_363), .B2(n_365), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g663 ( .A(n_361), .Y(n_663) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g498 ( .A(n_374), .Y(n_498) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_374), .Y(n_521) );
INVx1_ASAP7_75t_L g964 ( .A(n_374), .Y(n_964) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g414 ( .A(n_375), .Y(n_414) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
XNOR2x1_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_385), .B(n_405), .Y(n_384) );
NAND4xp25_ASAP7_75t_L g385 ( .A(n_386), .B(n_393), .C(n_396), .D(n_402), .Y(n_385) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx12f_ASAP7_75t_L g461 ( .A(n_388), .Y(n_461) );
INVx3_ASAP7_75t_L g566 ( .A(n_388), .Y(n_566) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_392), .Y(n_462) );
BUFx5_ASAP7_75t_L g476 ( .A(n_392), .Y(n_476) );
BUFx3_ASAP7_75t_L g716 ( .A(n_392), .Y(n_716) );
BUFx8_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_398), .Y(n_527) );
BUFx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_400), .Y(n_459) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_400), .Y(n_560) );
BUFx12f_ASAP7_75t_L g620 ( .A(n_400), .Y(n_620) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_400), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_421), .C(n_426), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_415), .Y(n_407) );
INVx4_ASAP7_75t_L g610 ( .A(n_409), .Y(n_610) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
INVx1_ASAP7_75t_L g508 ( .A(n_410), .Y(n_508) );
BUFx3_ASAP7_75t_L g654 ( .A(n_410), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_413), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_413), .B(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_413), .B(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx4_ASAP7_75t_L g542 ( .A(n_414), .Y(n_542) );
INVx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g511 ( .A(n_417), .Y(n_511) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_418), .Y(n_444) );
BUFx3_ASAP7_75t_L g483 ( .A(n_418), .Y(n_483) );
BUFx6f_ASAP7_75t_L g681 ( .A(n_418), .Y(n_681) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_420), .Y(n_445) );
INVx3_ASAP7_75t_L g485 ( .A(n_420), .Y(n_485) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g454 ( .A(n_424), .Y(n_454) );
INVx2_ASAP7_75t_L g679 ( .A(n_424), .Y(n_679) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
BUFx3_ASAP7_75t_L g491 ( .A(n_425), .Y(n_491) );
INVx2_ASAP7_75t_L g515 ( .A(n_425), .Y(n_515) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx4_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
INVx3_ASAP7_75t_L g569 ( .A(n_428), .Y(n_569) );
INVx2_ASAP7_75t_L g677 ( .A(n_428), .Y(n_677) );
INVx5_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g448 ( .A(n_429), .Y(n_448) );
BUFx4f_ASAP7_75t_L g612 ( .A(n_429), .Y(n_612) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g572 ( .A(n_431), .Y(n_572) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_431), .Y(n_708) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_433), .Y(n_447) );
BUFx3_ASAP7_75t_L g509 ( .A(n_433), .Y(n_509) );
INVx1_ASAP7_75t_L g499 ( .A(n_436), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_467), .B2(n_468), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_455), .Y(n_441) );
NAND4xp25_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .C(n_449), .D(n_453), .Y(n_442) );
INVx2_ASAP7_75t_L g703 ( .A(n_444), .Y(n_703) );
INVx3_ASAP7_75t_L g606 ( .A(n_445), .Y(n_606) );
INVx3_ASAP7_75t_L g604 ( .A(n_447), .Y(n_604) );
NAND4xp25_ASAP7_75t_SL g455 ( .A(n_456), .B(n_460), .C(n_463), .D(n_465), .Y(n_455) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx4f_ASAP7_75t_L g689 ( .A(n_458), .Y(n_689) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
NAND4xp75_ASAP7_75t_SL g469 ( .A(n_470), .B(n_474), .C(n_479), .D(n_486), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_482), .Y(n_479) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g722 ( .A(n_491), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_496), .B2(n_497), .Y(n_492) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_553), .B1(n_593), .B2(n_594), .Y(n_500) );
INVx1_ASAP7_75t_L g593 ( .A(n_501), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_528), .B1(n_551), .B2(n_552), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g551 ( .A(n_503), .Y(n_551) );
NOR2x1_ASAP7_75t_SL g504 ( .A(n_505), .B(n_522), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .C(n_512), .Y(n_505) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_515), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_519), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_518), .A2(n_659), .B1(n_661), .B2(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_521), .B(n_684), .Y(n_683) );
NAND4xp25_ASAP7_75t_SL g522 ( .A(n_523), .B(n_524), .C(n_525), .D(n_526), .Y(n_522) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_530), .Y(n_552) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_543), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .C(n_537), .D(n_539), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_542), .B(n_585), .Y(n_584) );
INVx4_ASAP7_75t_L g627 ( .A(n_542), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_542), .B(n_634), .Y(n_633) );
NAND4xp25_ASAP7_75t_L g543 ( .A(n_544), .B(n_546), .C(n_547), .D(n_548), .Y(n_543) );
INVx1_ASAP7_75t_L g594 ( .A(n_553), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_574), .B2(n_591), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
NOR2x1_ASAP7_75t_L g556 ( .A(n_557), .B(n_567), .Y(n_556) );
NAND4xp25_ASAP7_75t_SL g557 ( .A(n_558), .B(n_559), .C(n_561), .D(n_563), .Y(n_557) );
BUFx4f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g955 ( .A(n_566), .Y(n_955) );
NAND4xp25_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .C(n_571), .D(n_573), .Y(n_567) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
BUFx3_ASAP7_75t_L g592 ( .A(n_576), .Y(n_592) );
XNOR2x1_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_586), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .C(n_582), .D(n_583), .Y(n_579) );
NAND4xp25_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .C(n_589), .D(n_590), .Y(n_586) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
XNOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_647), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_628), .B1(n_644), .B2(n_645), .Y(n_598) );
INVx1_ASAP7_75t_L g644 ( .A(n_599), .Y(n_644) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND4xp75_ASAP7_75t_L g601 ( .A(n_602), .B(n_613), .C(n_617), .D(n_621), .Y(n_601) );
NOR2xp67_ASAP7_75t_L g602 ( .A(n_603), .B(n_608), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_605), .B1(n_606), .B2(n_607), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_606), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_610), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g960 ( .A(n_623), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVxp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_630), .Y(n_646) );
NAND3x1_ASAP7_75t_L g631 ( .A(n_632), .B(n_635), .C(n_639), .Y(n_631) );
AND2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND4x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .C(n_642), .D(n_643), .Y(n_639) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AO22x2_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_692), .B2(n_693), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
XOR2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_672), .Y(n_649) );
INVx1_ASAP7_75t_L g671 ( .A(n_651), .Y(n_671) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_665), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_657), .C(n_664), .Y(n_652) );
CKINVDCx16_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
CKINVDCx9p33_ASAP7_75t_R g661 ( .A(n_662), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .C(n_668), .D(n_669), .Y(n_665) );
XNOR2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_675), .B(n_685), .Y(n_674) );
NAND4xp25_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .C(n_680), .D(n_682), .Y(n_675) );
NAND4xp25_ASAP7_75t_SL g685 ( .A(n_686), .B(n_688), .C(n_690), .D(n_691), .Y(n_685) );
BUFx2_ASAP7_75t_L g697 ( .A(n_687), .Y(n_697) );
INVx2_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND4xp75_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .C(n_709), .D(n_717), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_705), .Y(n_700) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B(n_723), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_946), .B(n_948), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_873), .C(n_911), .Y(n_725) );
OAI221xp5_ASAP7_75t_SL g726 ( .A1(n_727), .A2(n_831), .B1(n_832), .B2(n_837), .C(n_857), .Y(n_726) );
NOR4xp25_ASAP7_75t_L g727 ( .A(n_728), .B(n_802), .C(n_816), .D(n_824), .Y(n_727) );
OAI211xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_750), .B(n_768), .C(n_795), .Y(n_728) );
INVx1_ASAP7_75t_L g800 ( .A(n_729), .Y(n_800) );
NOR2x1_ASAP7_75t_L g899 ( .A(n_729), .B(n_805), .Y(n_899) );
OR2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_742), .Y(n_729) );
INVx1_ASAP7_75t_L g786 ( .A(n_730), .Y(n_786) );
AND2x2_ASAP7_75t_L g815 ( .A(n_730), .B(n_779), .Y(n_815) );
AND2x2_ASAP7_75t_L g821 ( .A(n_730), .B(n_742), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_730), .B(n_776), .Y(n_909) );
OAI321xp33_ASAP7_75t_L g930 ( .A1(n_730), .A2(n_813), .A3(n_905), .B1(n_931), .B2(n_932), .C(n_934), .Y(n_930) );
AND2x2_ASAP7_75t_L g944 ( .A(n_730), .B(n_775), .Y(n_944) );
INVx3_ASAP7_75t_L g835 ( .A(n_731), .Y(n_835) );
AND2x4_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
AND2x4_ASAP7_75t_L g739 ( .A(n_732), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g748 ( .A(n_732), .B(n_740), .Y(n_748) );
AND2x2_ASAP7_75t_L g757 ( .A(n_732), .B(n_740), .Y(n_757) );
AND2x4_ASAP7_75t_L g736 ( .A(n_734), .B(n_737), .Y(n_736) );
AND2x4_ASAP7_75t_L g746 ( .A(n_734), .B(n_737), .Y(n_746) );
AND2x2_ASAP7_75t_L g741 ( .A(n_737), .B(n_740), .Y(n_741) );
AND2x2_ASAP7_75t_L g749 ( .A(n_737), .B(n_740), .Y(n_749) );
AND2x4_ASAP7_75t_L g758 ( .A(n_737), .B(n_740), .Y(n_758) );
BUFx2_ASAP7_75t_L g947 ( .A(n_739), .Y(n_947) );
INVx1_ASAP7_75t_L g779 ( .A(n_742), .Y(n_779) );
AND2x2_ASAP7_75t_L g791 ( .A(n_742), .B(n_776), .Y(n_791) );
AND2x2_ASAP7_75t_L g810 ( .A(n_742), .B(n_786), .Y(n_810) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_747), .Y(n_742) );
INVx2_ASAP7_75t_SL g755 ( .A(n_746), .Y(n_755) );
INVx1_ASAP7_75t_L g927 ( .A(n_750), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_751), .B(n_759), .Y(n_750) );
AND2x2_ASAP7_75t_L g787 ( .A(n_751), .B(n_764), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_751), .B(n_789), .Y(n_811) );
AND2x2_ASAP7_75t_L g823 ( .A(n_751), .B(n_813), .Y(n_823) );
OR2x2_ASAP7_75t_L g849 ( .A(n_751), .B(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_751), .B(n_771), .Y(n_905) );
NOR2xp33_ASAP7_75t_L g925 ( .A(n_751), .B(n_831), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_751), .B(n_830), .Y(n_941) );
INVx4_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g840 ( .A(n_752), .B(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g846 ( .A(n_752), .B(n_765), .Y(n_846) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_752), .B(n_810), .C(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g863 ( .A(n_752), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_752), .B(n_832), .Y(n_885) );
AND2x2_ASAP7_75t_L g888 ( .A(n_752), .B(n_813), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_752), .B(n_842), .Y(n_933) );
NOR3xp33_ASAP7_75t_SL g935 ( .A(n_752), .B(n_866), .C(n_902), .Y(n_935) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .Y(n_752) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI332xp33_ASAP7_75t_L g900 ( .A1(n_760), .A2(n_845), .A3(n_901), .B1(n_904), .B2(n_905), .B3(n_906), .C1(n_907), .C2(n_910), .Y(n_900) );
OAI222xp33_ASAP7_75t_SL g917 ( .A1(n_760), .A2(n_775), .B1(n_830), .B2(n_918), .C1(n_922), .C2(n_923), .Y(n_917) );
OR2x2_ASAP7_75t_L g760 ( .A(n_761), .B(n_764), .Y(n_760) );
INVx4_ASAP7_75t_L g784 ( .A(n_761), .Y(n_784) );
OR2x2_ASAP7_75t_L g830 ( .A(n_761), .B(n_765), .Y(n_830) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_761), .B(n_794), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_761), .B(n_771), .Y(n_852) );
AND2x2_ASAP7_75t_L g855 ( .A(n_761), .B(n_764), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_761), .B(n_794), .Y(n_866) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx2_ASAP7_75t_L g789 ( .A(n_764), .Y(n_789) );
OR2x2_ASAP7_75t_L g842 ( .A(n_764), .B(n_784), .Y(n_842) );
INVxp67_ASAP7_75t_L g850 ( .A(n_764), .Y(n_850) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_780), .B(n_787), .C(n_788), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_774), .Y(n_769) );
AND2x2_ASAP7_75t_L g818 ( .A(n_770), .B(n_814), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_770), .B(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_770), .B(n_809), .Y(n_892) );
AND2x2_ASAP7_75t_L g945 ( .A(n_770), .B(n_841), .Y(n_945) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g794 ( .A(n_771), .Y(n_794) );
AND2x2_ASAP7_75t_L g801 ( .A(n_771), .B(n_775), .Y(n_801) );
INVx3_ASAP7_75t_L g806 ( .A(n_771), .Y(n_806) );
AOI211xp5_ASAP7_75t_L g837 ( .A1(n_771), .A2(n_838), .B(n_843), .C(n_853), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g908 ( .A(n_771), .B(n_909), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_771), .B(n_855), .Y(n_922) );
AND2x2_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g879 ( .A(n_774), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_779), .Y(n_774) );
AND2x2_ASAP7_75t_L g808 ( .A(n_775), .B(n_800), .Y(n_808) );
AND2x2_ASAP7_75t_L g820 ( .A(n_775), .B(n_821), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_775), .B(n_810), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_775), .B(n_861), .Y(n_860) );
AND2x2_ASAP7_75t_L g867 ( .A(n_775), .B(n_815), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_775), .B(n_899), .Y(n_898) );
CKINVDCx6p67_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_776), .B(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g809 ( .A(n_776), .B(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g814 ( .A(n_776), .B(n_815), .Y(n_814) );
AND2x2_ASAP7_75t_L g829 ( .A(n_776), .B(n_800), .Y(n_829) );
AND2x2_ASAP7_75t_L g871 ( .A(n_776), .B(n_805), .Y(n_871) );
AND2x2_ASAP7_75t_L g915 ( .A(n_776), .B(n_861), .Y(n_915) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_776), .B(n_779), .Y(n_921) );
AND2x2_ASAP7_75t_L g928 ( .A(n_776), .B(n_779), .Y(n_928) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_779), .B(n_848), .Y(n_847) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_785), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_781), .B(n_870), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g912 ( .A1(n_781), .A2(n_913), .B1(n_915), .B2(n_916), .C(n_917), .Y(n_912) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_782), .Y(n_916) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g793 ( .A(n_783), .Y(n_793) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g813 ( .A(n_784), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_786), .A2(n_804), .B1(n_875), .B2(n_877), .C(n_880), .Y(n_874) );
AOI221xp5_ASAP7_75t_L g893 ( .A1(n_787), .A2(n_894), .B1(n_895), .B2(n_897), .C(n_900), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_787), .B(n_891), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx3_ASAP7_75t_SL g804 ( .A(n_789), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_789), .B(n_831), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_789), .B(n_832), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_792), .Y(n_790) );
INVx1_ASAP7_75t_L g906 ( .A(n_791), .Y(n_906) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx1_ASAP7_75t_L g798 ( .A(n_793), .Y(n_798) );
NOR2xp33_ASAP7_75t_L g919 ( .A(n_794), .B(n_920), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_799), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_796), .B(n_898), .Y(n_897) );
HB1xp67_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g891 ( .A(n_798), .Y(n_891) );
AND2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
AND2x2_ASAP7_75t_L g870 ( .A(n_800), .B(n_871), .Y(n_870) );
INVxp67_ASAP7_75t_L g904 ( .A(n_801), .Y(n_904) );
OAI22xp33_ASAP7_75t_SL g802 ( .A1(n_803), .A2(n_807), .B1(n_811), .B2(n_812), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_805), .Y(n_803) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_804), .A2(n_927), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_926) );
NOR2x1_ASAP7_75t_L g826 ( .A(n_805), .B(n_827), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_805), .B(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g894 ( .A(n_805), .B(n_856), .Y(n_894) );
INVx3_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
AND2x2_ASAP7_75t_L g861 ( .A(n_806), .B(n_821), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_L g942 ( .A(n_808), .Y(n_942) );
INVx1_ASAP7_75t_L g844 ( .A(n_809), .Y(n_844) );
OAI21xp5_ASAP7_75t_L g943 ( .A1(n_809), .A2(n_944), .B(n_945), .Y(n_943) );
INVx1_ASAP7_75t_L g902 ( .A(n_810), .Y(n_902) );
INVx1_ASAP7_75t_L g858 ( .A(n_811), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
O2A1O1Ixp33_ASAP7_75t_L g868 ( .A1(n_813), .A2(n_819), .B(n_869), .C(n_872), .Y(n_868) );
INVx1_ASAP7_75t_L g923 ( .A(n_814), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_815), .B(n_840), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_815), .B(n_871), .Y(n_883) );
INVx1_ASAP7_75t_L g903 ( .A(n_815), .Y(n_903) );
AOI21xp5_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_819), .B(n_822), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_821), .B(n_871), .Y(n_914) );
INVx1_ASAP7_75t_L g931 ( .A(n_821), .Y(n_931) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
AOI21xp33_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_828), .B(n_830), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g856 ( .A(n_827), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_828), .B(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
CKINVDCx5p33_ASAP7_75t_R g831 ( .A(n_832), .Y(n_831) );
OAI221xp5_ASAP7_75t_SL g873 ( .A1(n_832), .A2(n_874), .B1(n_884), .B2(n_886), .C(n_893), .Y(n_873) );
OAI221xp5_ASAP7_75t_SL g911 ( .A1(n_832), .A2(n_912), .B1(n_924), .B2(n_926), .C(n_936), .Y(n_911) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_836), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVxp67_ASAP7_75t_SL g838 ( .A(n_839), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_840), .A2(n_877), .B1(n_937), .B2(n_938), .C(n_939), .Y(n_936) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B1(n_847), .B2(n_849), .C(n_851), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVxp67_ASAP7_75t_SL g853 ( .A(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g876 ( .A(n_855), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_855), .B(n_882), .Y(n_881) );
AOI211xp5_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_859), .B(n_862), .C(n_868), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_859), .A2(n_887), .B(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVxp67_ASAP7_75t_SL g938 ( .A(n_872), .Y(n_938) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVxp67_ASAP7_75t_SL g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .Y(n_889) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g937 ( .A(n_892), .Y(n_937) );
INVxp67_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g929 ( .A(n_898), .Y(n_929) );
AND2x2_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVxp67_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVxp67_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
OAI21xp5_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_942), .B(n_943), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_947), .Y(n_946) );
XOR2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_965), .Y(n_949) );
INVxp33_ASAP7_75t_L g971 ( .A(n_950), .Y(n_971) );
NOR2x1_ASAP7_75t_L g950 ( .A(n_951), .B(n_958), .Y(n_950) );
NAND4xp25_ASAP7_75t_L g951 ( .A(n_952), .B(n_953), .C(n_954), .D(n_956), .Y(n_951) );
NAND4xp25_ASAP7_75t_L g958 ( .A(n_959), .B(n_961), .C(n_962), .D(n_963), .Y(n_958) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_SL g973 ( .A(n_971), .Y(n_973) );
BUFx2_ASAP7_75t_SL g974 ( .A(n_975), .Y(n_974) );
BUFx2_ASAP7_75t_L g976 ( .A(n_977), .Y(n_976) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_979), .Y(n_978) );
endmodule