module real_jpeg_17747_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_556;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_0),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B(n_581),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_1),
.B(n_582),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_61)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_2),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_67),
.B1(n_172),
.B2(n_178),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_2),
.A2(n_67),
.B1(n_202),
.B2(n_205),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_2),
.A2(n_67),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_4),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g432 ( 
.A(n_4),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_5),
.A2(n_237),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_5),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_5),
.A2(n_244),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_5),
.A2(n_244),
.B1(n_450),
.B2(n_452),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_SL g506 ( 
.A1(n_5),
.A2(n_244),
.B1(n_507),
.B2(n_512),
.Y(n_506)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_6),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_6),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_7),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_7),
.Y(n_145)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_7),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_7),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g227 ( 
.A(n_7),
.Y(n_227)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_7),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_7),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_7),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_8),
.A2(n_39),
.B1(n_103),
.B2(n_106),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_39),
.B1(n_152),
.B2(n_156),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_8),
.A2(n_39),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_9),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_10),
.A2(n_123),
.B1(n_286),
.B2(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_10),
.A2(n_316),
.B1(n_360),
.B2(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_10),
.A2(n_316),
.B1(n_440),
.B2(n_445),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_10),
.A2(n_316),
.B1(n_482),
.B2(n_483),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_12),
.A2(n_281),
.A3(n_285),
.B1(n_287),
.B2(n_292),
.Y(n_280)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_12),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_12),
.A2(n_69),
.B1(n_291),
.B2(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_12),
.B(n_24),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_12),
.B(n_73),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_12),
.B(n_491),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_12),
.B(n_132),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g514 ( 
.A1(n_12),
.A2(n_174),
.B1(n_291),
.B2(n_515),
.Y(n_514)
);

OAI32xp33_ASAP7_75t_L g518 ( 
.A1(n_12),
.A2(n_519),
.A3(n_521),
.B1(n_522),
.B2(n_526),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_14),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_122)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_14),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_14),
.A2(n_128),
.B1(n_224),
.B2(n_228),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_14),
.A2(n_128),
.B1(n_299),
.B2(n_305),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_14),
.A2(n_128),
.B1(n_333),
.B2(n_337),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_15),
.Y(n_134)
);

BUFx4f_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_15),
.Y(n_198)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_15),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_16),
.A2(n_49),
.B1(n_112),
.B2(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_16),
.A2(n_49),
.B1(n_215),
.B2(n_218),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_16),
.A2(n_49),
.B1(n_226),
.B2(n_232),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_161),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_159),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_22),
.B(n_59),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_44),
.Y(n_22)
);

OAI21x1_ASAP7_75t_SL g338 ( 
.A1(n_23),
.A2(n_51),
.B(n_243),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

OR2x6_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_24),
.B(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_24),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_24),
.A2(n_50),
.B1(n_314),
.B2(n_317),
.Y(n_313)
);

AO22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_30),
.Y(n_177)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_30),
.Y(n_373)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_33),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_34),
.Y(n_181)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_38),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_41),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_41),
.Y(n_245)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21x1_ASAP7_75t_SL g168 ( 
.A1(n_44),
.A2(n_122),
.B(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_61),
.B(n_71),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_51),
.A2(n_61),
.B1(n_122),
.B2(n_129),
.Y(n_121)
);

OAI22x1_ASAP7_75t_SL g235 ( 
.A1(n_51),
.A2(n_129),
.B1(n_236),
.B2(n_243),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_51),
.A2(n_129),
.B1(n_315),
.B2(n_352),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_51),
.A2(n_71),
.B(n_403),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_56),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_58),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_59),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_59),
.B(n_164),
.Y(n_580)
);

FAx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_72),
.CI(n_108),
.CON(n_59),
.SN(n_59)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_85),
.B(n_101),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_73),
.B(n_111),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_73),
.A2(n_85),
.B1(n_171),
.B2(n_394),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_78),
.B2(n_81),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_76),
.Y(n_438)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_77),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_78),
.Y(n_459)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_79),
.Y(n_263)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_83),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g110 ( 
.A1(n_85),
.A2(n_111),
.B(n_118),
.Y(n_110)
);

AOI21x1_ASAP7_75t_L g170 ( 
.A1(n_85),
.A2(n_171),
.B(n_182),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_85),
.A2(n_118),
.B(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_86),
.A2(n_102),
.B(n_183),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_86),
.A2(n_119),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_86),
.A2(n_119),
.B1(n_272),
.B2(n_356),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g369 ( 
.A1(n_86),
.A2(n_119),
.B1(n_356),
.B2(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_86),
.A2(n_119),
.B1(n_370),
.B2(n_514),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_92),
.Y(n_273)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_102),
.B(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_104),
.Y(n_529)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_105),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_120),
.C(n_130),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_109),
.A2(n_110),
.B1(n_130),
.B2(n_131),
.Y(n_167)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_111),
.Y(n_331)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_125),
.Y(n_294)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_126),
.Y(n_286)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_168),
.C(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_131),
.B(n_170),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_141),
.B(n_150),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_132),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_132),
.B(n_231),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_132),
.A2(n_141),
.B1(n_437),
.B2(n_439),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_132),
.A2(n_141),
.B1(n_439),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_133),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_133),
.B(n_151),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_133),
.A2(n_260),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

OA22x2_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_133)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_134),
.Y(n_451)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_134),
.Y(n_489)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_135),
.Y(n_426)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_137),
.Y(n_255)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_138),
.Y(n_256)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_138),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_141),
.B(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_141),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_141),
.A2(n_397),
.B(n_542),
.Y(n_541)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_144),
.Y(n_233)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_145),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_149),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_151),
.A2(n_260),
.B(n_326),
.Y(n_350)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_184),
.B(n_579),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_166),
.A2(n_168),
.B1(n_560),
.B2(n_561),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_166),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_168),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_168),
.A2(n_561),
.B1(n_564),
.B2(n_565),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_169),
.B(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_178),
.Y(n_360)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_181),
.Y(n_520)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_556),
.B(n_576),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_408),
.Y(n_185)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_343),
.B(n_384),
.C(n_385),
.D(n_407),
.Y(n_186)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_187),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_318),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_188),
.B(n_318),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_247),
.C(n_268),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_189),
.A2(n_190),
.B1(n_247),
.B2(n_248),
.Y(n_345)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_234),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_191),
.B(n_235),
.C(n_246),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_221),
.Y(n_191)
);

XOR2x2_ASAP7_75t_L g361 ( 
.A(n_192),
.B(n_221),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_201),
.B(n_208),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_193),
.A2(n_201),
.B1(n_298),
.B2(n_309),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_193),
.A2(n_467),
.B1(n_472),
.B2(n_473),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_193),
.A2(n_208),
.B(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_194),
.B(n_214),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_194),
.A2(n_254),
.B(n_322),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_194),
.A2(n_449),
.B(n_455),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_194),
.A2(n_291),
.B1(n_480),
.B2(n_481),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_194),
.A2(n_468),
.B1(n_481),
.B2(n_495),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_196),
.Y(n_483)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_197),
.Y(n_454)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_198),
.Y(n_424)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_213),
.Y(n_492)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_230),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_233),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_240),
.B2(n_242),
.Y(n_236)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_238),
.Y(n_354)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_239),
.A2(n_242),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_239),
.A2(n_242),
.B1(n_459),
.B2(n_460),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_239),
.A2(n_242),
.B1(n_433),
.B2(n_469),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_258),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_249),
.B(n_258),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_250),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_254),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_257),
.A2(n_298),
.B(n_378),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_260),
.A2(n_261),
.B(n_326),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_267),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_268),
.B(n_345),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_279),
.C(n_313),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_270),
.B(n_313),
.Y(n_348)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_276),
.Y(n_516)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_278),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_279),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_297),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_280),
.B(n_297),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_291),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_291),
.B(n_428),
.Y(n_427)
);

OAI21xp33_ASAP7_75t_SL g437 ( 
.A1(n_291),
.A2(n_427),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_291),
.B(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_304),
.Y(n_308)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_312),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_328),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_320),
.B(n_328),
.C(n_340),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_324),
.B1(n_325),
.B2(n_327),
.Y(n_320)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_SL g400 ( 
.A(n_321),
.B(n_325),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_321),
.A2(n_327),
.B1(n_402),
.B2(n_404),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

AOI21xp33_ASAP7_75t_L g568 ( 
.A1(n_327),
.A2(n_404),
.B(n_569),
.Y(n_568)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_339),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_338),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g394 ( 
.A(n_332),
.Y(n_394)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_339),
.C(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_346),
.C(n_362),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_346),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.C(n_361),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_361),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.C(n_355),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_355),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx2_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_382),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_363),
.B(n_382),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.C(n_368),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_364),
.B(n_553),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_366),
.A2(n_367),
.B1(n_368),
.B2(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_368),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_374),
.C(n_376),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_369),
.B(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_374),
.A2(n_375),
.B1(n_377),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_377),
.Y(n_546)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_378),
.Y(n_495)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_381),
.Y(n_474)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_410),
.C(n_413),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_388),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_389),
.B(n_399),
.C(n_405),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_399),
.B1(n_405),
.B2(n_406),
.Y(n_391)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_392),
.Y(n_405)
);

OAI21xp33_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_395),
.B(n_398),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_395),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_398),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_398),
.A2(n_563),
.B1(n_566),
.B2(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_399),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_400),
.Y(n_569)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_402),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_414),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_549),
.B(n_555),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_536),
.B(n_548),
.Y(n_415)
);

OAI21x1_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_500),
.B(n_535),
.Y(n_416)
);

AOI21x1_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_464),
.B(n_499),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_447),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_419),
.B(n_447),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_435),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_420),
.A2(n_435),
.B1(n_436),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_420),
.Y(n_476)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.A3(n_425),
.B1(n_427),
.B2(n_430),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_424),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_429),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_444),
.Y(n_525)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_456),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_457),
.C(n_463),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_463),
.Y(n_456)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_458),
.Y(n_505)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_465),
.A2(n_477),
.B(n_498),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_475),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_475),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_493),
.B(n_497),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_484),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_490),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_494),
.B(n_496),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_502),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_501),
.B(n_502),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_517),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_513),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_504),
.B(n_513),
.C(n_517),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_506),
.Y(n_542)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_510),
.Y(n_521)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_533),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_518),
.B(n_533),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_530),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_538),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_537),
.B(n_538),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_539),
.A2(n_543),
.B1(n_544),
.B2(n_547),
.Y(n_538)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_539),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_540),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_541),
.B(n_543),
.C(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_552),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_550),
.B(n_552),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_570),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_557),
.A2(n_577),
.B(n_578),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_562),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g578 ( 
.A(n_558),
.B(n_562),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_566),
.C(n_567),
.Y(n_562)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_563),
.Y(n_575)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_564),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_567),
.A2(n_568),
.B1(n_573),
.B2(n_574),
.Y(n_572)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

NOR2xp67_ASAP7_75t_SL g570 ( 
.A(n_571),
.B(n_572),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_571),
.B(n_572),
.Y(n_577)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);


endmodule