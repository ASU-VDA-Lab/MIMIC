module real_jpeg_4978_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_0),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_0),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_0),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_0),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_0),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_0),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_0),
.B(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_1),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_2),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_2),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_2),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_2),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_3),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_121),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_3),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_139),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_3),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_4),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_4),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_4),
.B(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_4),
.B(n_319),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_4),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_4),
.B(n_131),
.Y(n_419)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_5),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g409 ( 
.A(n_5),
.Y(n_409)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_6),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_7),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_7),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_7),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_7),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_8),
.Y(n_70)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_8),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_8),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_8),
.Y(n_358)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_12),
.B(n_45),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_12),
.B(n_31),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_12),
.B(n_310),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_12),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_12),
.B(n_349),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_12),
.B(n_391),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_12),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_13),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_13),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_13),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_13),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_13),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_13),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_14),
.B(n_106),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_14),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_14),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_14),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_14),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_14),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_14),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_14),
.B(n_415),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_15),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_106),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_16),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_16),
.B(n_121),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_188),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_16),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_16),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_16),
.B(n_424),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_17),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_17),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_17),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_17),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_17),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_17),
.B(n_319),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_17),
.B(n_376),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_17),
.B(n_417),
.Y(n_416)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_19),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_19),
.B(n_224),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_19),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_19),
.B(n_73),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_19),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_19),
.B(n_388),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_19),
.B(n_407),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_517),
.B(n_520),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_169),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_168),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_110),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_25),
.B(n_110),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_89),
.B1(n_90),
.B2(n_109),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_26),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_58),
.C(n_77),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_27),
.A2(n_28),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_41),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_30),
.B(n_34),
.C(n_41),
.Y(n_108)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_40),
.Y(n_136)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_40),
.Y(n_158)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_40),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.C(n_54),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_42),
.B(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_45),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_46),
.A2(n_47),
.B1(n_54),
.B2(n_55),
.Y(n_143)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_52),
.Y(n_192)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_53),
.Y(n_356)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_53),
.Y(n_393)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_53),
.Y(n_415)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_57),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_58),
.A2(n_77),
.B1(n_78),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.C(n_71),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_59),
.B(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_64),
.A2(n_65),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_64),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_161)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_65),
.B(n_134),
.C(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_70),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_71),
.A2(n_72),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_84),
.C(n_88),
.Y(n_99)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_76),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_76),
.Y(n_352)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_76),
.Y(n_385)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B1(n_83),
.B2(n_88),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_85),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_86),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_108),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_99),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_159),
.C(n_164),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_111),
.A2(n_112),
.B1(n_499),
.B2(n_500),
.Y(n_498)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_142),
.C(n_144),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_113),
.B(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_125),
.C(n_133),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_114),
.A2(n_115),
.B1(n_125),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_118),
.C(n_122),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_125),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.C(n_130),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_126),
.B(n_130),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_127),
.B(n_248),
.Y(n_247)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_129),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_133),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_147),
.C(n_149),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_138),
.A2(n_141),
.B1(n_149),
.B2(n_150),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_140),
.Y(n_311)
);

BUFx8_ASAP7_75t_L g328 ( 
.A(n_140),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_142),
.Y(n_505)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_152),
.C(n_156),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_146),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_147),
.B(n_245),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_149),
.A2(n_150),
.B1(n_199),
.B2(n_203),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_150),
.B(n_194),
.C(n_199),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_242)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_157),
.B1(n_206),
.B2(n_210),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_157),
.B(n_210),
.C(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_158),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_159),
.B(n_164),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_160),
.B(n_507),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_162),
.B(n_163),
.Y(n_507)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_496),
.B(n_514),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_298),
.B(n_495),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_249),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_173),
.B(n_249),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_233),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_174),
.B(n_234),
.C(n_237),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_204),
.C(n_212),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_175),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_184),
.C(n_193),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_176),
.B(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_180),
.C(n_181),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_184),
.A2(n_185),
.B1(n_193),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.C(n_189),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_186),
.B(n_189),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_187),
.B(n_471),
.Y(n_470)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_193),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_212),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.Y(n_204)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.C(n_228),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_213),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.C(n_220),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_214),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_220),
.Y(n_261)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_219),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_219),
.Y(n_376)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_222),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_222),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_228),
.Y(n_278)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_227),
.Y(n_286)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_232),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_232),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_243),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_239),
.B(n_241),
.C(n_243),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_251),
.B(n_254),
.Y(n_491)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_256),
.B(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_276),
.C(n_279),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_258),
.B(n_484),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_268),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_259),
.A2(n_260),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_262),
.A2(n_263),
.B(n_265),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_262),
.B(n_268),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.C(n_273),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_439)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_273),
.B(n_439),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_275),
.B(n_369),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_279),
.Y(n_485)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.C(n_295),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_281),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_281),
.B(n_473),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_287),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_282),
.B(n_451),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_284),
.A2(n_287),
.B1(n_288),
.B2(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_284),
.Y(n_452)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_291),
.B(n_295),
.Y(n_473)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_489),
.B(n_494),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_476),
.B(n_488),
.Y(n_299)
);

AOI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_458),
.B(n_475),
.Y(n_300)
);

OAI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_432),
.B(n_457),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_397),
.B(n_431),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_361),
.B(n_396),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_338),
.B(n_360),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_322),
.B(n_337),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_317),
.B(n_321),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_316),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_316),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_312),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_312),
.Y(n_323)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_311),
.Y(n_425)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx8_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_324),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_330),
.B2(n_331),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_325),
.B(n_333),
.C(n_335),
.Y(n_359)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_329),
.Y(n_346)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_359),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_359),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_347),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_341),
.B(n_346),
.C(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_342),
.B(n_345),
.Y(n_366)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_347),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_380),
.C(n_381),
.Y(n_379)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_357),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx6_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_364),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_362),
.B(n_364),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_378),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_379),
.C(n_382),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_366),
.B(n_368),
.C(n_371),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_374),
.B1(n_375),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_372),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_373),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_377),
.Y(n_410)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_382),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

MAJx2_ASAP7_75t_L g429 ( 
.A(n_383),
.B(n_390),
.C(n_394),
.Y(n_429)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_387),
.A2(n_390),
.B1(n_394),
.B2(n_395),
.Y(n_386)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_387),
.Y(n_394)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_390),
.Y(n_395)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_430),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_398),
.B(n_430),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_412),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_411),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_400),
.B(n_411),
.C(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_410),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_406),
.Y(n_401)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_402),
.Y(n_446)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_406),
.Y(n_447)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_446),
.C(n_447),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_412),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_420),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_422),
.C(n_428),
.Y(n_435)
);

BUFx24_ASAP7_75t_SL g523 ( 
.A(n_413),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.CI(n_419),
.CON(n_413),
.SN(n_413)
);

MAJx2_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_416),
.C(n_419),
.Y(n_443)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B1(n_428),
.B2(n_429),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_423),
.B(n_426),
.Y(n_442)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_455),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_455),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_444),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_436),
.C(n_444),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_437),
.A2(n_438),
.B1(n_440),
.B2(n_441),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_467),
.C(n_468),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_443),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_448),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_449),
.C(n_454),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_453),
.B2(n_454),
.Y(n_448)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_449),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_450),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_474),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_474),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_465),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_461),
.B(n_464),
.C(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_462),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_470),
.C(n_472),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_486),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_486),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_478),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_483),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_483),
.C(n_493),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_490),
.B(n_492),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_509),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_L g514 ( 
.A1(n_497),
.A2(n_515),
.B(n_516),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_498),
.B(n_501),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_501),
.Y(n_516)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_499),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_506),
.C(n_508),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_502),
.A2(n_503),
.B1(n_506),
.B2(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_506),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_508),
.B(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_510),
.B(n_513),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_513),
.Y(n_515)
);

BUFx12f_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_518),
.Y(n_521)
);

INVx13_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_522),
.Y(n_520)
);


endmodule