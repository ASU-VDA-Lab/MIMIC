module fake_jpeg_10209_n_257 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_19),
.B1(n_18),
.B2(n_34),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_61),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_49),
.B1(n_63),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_20),
.B1(n_29),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_20),
.B1(n_29),
.B2(n_21),
.Y(n_49)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_29),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_20),
.B1(n_32),
.B2(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_38),
.A2(n_26),
.B1(n_32),
.B2(n_21),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_27),
.B1(n_30),
.B2(n_33),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_43),
.B(n_26),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_65),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g66 ( 
.A1(n_53),
.A2(n_43),
.B(n_3),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_26),
.B(n_32),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_77),
.Y(n_116)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_74),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_73),
.B1(n_71),
.B2(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_27),
.B1(n_30),
.B2(n_24),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_17),
.B1(n_22),
.B2(n_58),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_59),
.A2(n_36),
.B(n_17),
.C(n_24),
.Y(n_72)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_80),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_2),
.B(n_4),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_79),
.B(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_86),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_57),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_96),
.B(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_112),
.B1(n_80),
.B2(n_76),
.Y(n_118)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_23),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_111),
.Y(n_131)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_64),
.B1(n_56),
.B2(n_60),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_115),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_117),
.B(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_113),
.A2(n_95),
.B1(n_92),
.B2(n_105),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_122),
.B1(n_128),
.B2(n_132),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_115),
.B(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_116),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_87),
.B1(n_91),
.B2(n_60),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_129),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_81),
.B1(n_73),
.B2(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_134),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_83),
.B1(n_72),
.B2(n_82),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_64),
.B1(n_56),
.B2(n_89),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_136),
.B1(n_99),
.B2(n_54),
.Y(n_160)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_84),
.B(n_78),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_135),
.A2(n_111),
.B(n_102),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_106),
.A2(n_54),
.B1(n_90),
.B2(n_44),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_138),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_130),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_141),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_110),
.B1(n_106),
.B2(n_90),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_129),
.B1(n_139),
.B2(n_120),
.Y(n_168)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_148),
.A2(n_165),
.B1(n_124),
.B2(n_52),
.C(n_5),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_116),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_153),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_108),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_150),
.B(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_134),
.B(n_99),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_42),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_2),
.C(n_4),
.Y(n_178)
);

OAI22x1_ASAP7_75t_L g156 ( 
.A1(n_122),
.A2(n_67),
.B1(n_94),
.B2(n_114),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_163),
.B(n_122),
.C(n_57),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_158),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_140),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_167),
.B1(n_94),
.B2(n_52),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_44),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_44),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_169),
.B1(n_149),
.B2(n_157),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_122),
.B1(n_135),
.B2(n_123),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_152),
.B1(n_9),
.B2(n_10),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_42),
.C(n_124),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_178),
.C(n_183),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NAND2x1_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_5),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_6),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_144),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_16),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_147),
.C(n_143),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_159),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_145),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_187),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_205)
);

AOI221xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_15),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_153),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_151),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_158),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_197),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_196),
.A2(n_202),
.B1(n_171),
.B2(n_172),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_203),
.C(n_207),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_166),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_149),
.B1(n_160),
.B2(n_152),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_162),
.C(n_161),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_204),
.A2(n_205),
.B1(n_187),
.B2(n_179),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_178),
.B(n_168),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_12),
.C(n_13),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_182),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_209),
.A2(n_206),
.B(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_210),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_188),
.C(n_185),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_174),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_171),
.B(n_170),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_200),
.B(n_191),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_171),
.C(n_180),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_220),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_12),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_190),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_231),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_216),
.C(n_217),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_227),
.B(n_228),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_191),
.C(n_204),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_222),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_233),
.Y(n_246)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_237),
.B(n_233),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_239),
.C(n_213),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_230),
.B(n_211),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_218),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_208),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_207),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_245),
.C(n_212),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_243),
.B(n_244),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_246),
.A2(n_212),
.B1(n_227),
.B2(n_238),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_250),
.C(n_223),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_249),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_12),
.B(n_13),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_253),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_255),
.A2(n_248),
.B(n_13),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_254),
.Y(n_257)
);


endmodule