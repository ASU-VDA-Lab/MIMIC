module fake_jpeg_29454_n_12 (n_3, n_2, n_1, n_0, n_4, n_12);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_12;

wire n_11;
wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx1_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

AND2x6_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_0),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_SL g7 ( 
.A(n_4),
.B(n_3),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_5),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_8),
.B(n_9),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_L g9 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_8),
.B(n_7),
.C(n_1),
.Y(n_11)
);

A2O1A1O1Ixp25_ASAP7_75t_L g12 ( 
.A1(n_11),
.A2(n_0),
.B(n_1),
.C(n_3),
.D(n_10),
.Y(n_12)
);


endmodule