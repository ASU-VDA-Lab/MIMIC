module fake_aes_12741_n_505 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_505);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_505;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_486;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_295;
wire n_143;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g69 ( .A(n_66), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_37), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_12), .Y(n_71) );
BUFx2_ASAP7_75t_SL g72 ( .A(n_6), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_42), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_45), .Y(n_74) );
BUFx6f_ASAP7_75t_L g75 ( .A(n_49), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_22), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_36), .Y(n_77) );
INVx1_ASAP7_75t_SL g78 ( .A(n_29), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_16), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_8), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_28), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_31), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_35), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_34), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_13), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_61), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_19), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_30), .Y(n_89) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_58), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_67), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_51), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_48), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_21), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_62), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_23), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_24), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_39), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_68), .Y(n_101) );
INVxp33_ASAP7_75t_L g102 ( .A(n_10), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_54), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_46), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_6), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_55), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_104), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_75), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_70), .Y(n_110) );
AND2x2_ASAP7_75t_L g111 ( .A(n_102), .B(n_0), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_75), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_96), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_70), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_73), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_96), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_90), .B(n_0), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_105), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_75), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_84), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_75), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_75), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_79), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_94), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_80), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_75), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_71), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_95), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_69), .Y(n_130) );
INVx2_ASAP7_75t_SL g131 ( .A(n_110), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_108), .B(n_104), .Y(n_132) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_111), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_128), .B(n_71), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_130), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_121), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_128), .B(n_76), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_110), .B(n_69), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_114), .B(n_74), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_130), .Y(n_141) );
NOR2xp33_ASAP7_75t_SL g142 ( .A(n_114), .B(n_85), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_130), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_128), .B(n_76), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_130), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_130), .Y(n_147) );
BUFx4f_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_118), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_119), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_119), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_108), .B(n_74), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_113), .Y(n_153) );
INVxp67_ASAP7_75t_L g154 ( .A(n_111), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_109), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_131), .B(n_126), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_150), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_131), .B(n_126), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_150), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
NOR2xp33_ASAP7_75t_R g165 ( .A(n_153), .B(n_116), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_131), .B(n_119), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_154), .B(n_129), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_148), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
NAND2xp33_ASAP7_75t_SL g171 ( .A(n_133), .B(n_111), .Y(n_171) );
BUFx2_ASAP7_75t_L g172 ( .A(n_137), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_155), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
CKINVDCx8_ASAP7_75t_R g175 ( .A(n_136), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_148), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_148), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
NOR2xp33_ASAP7_75t_SL g181 ( .A(n_142), .B(n_115), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_133), .B(n_154), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_137), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_142), .B(n_115), .Y(n_185) );
NOR3xp33_ASAP7_75t_SL g186 ( .A(n_153), .B(n_125), .C(n_124), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
NOR3xp33_ASAP7_75t_SL g189 ( .A(n_149), .B(n_125), .C(n_117), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_166), .A2(n_137), .B(n_132), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_157), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_183), .B(n_137), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_166), .A2(n_137), .B(n_132), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_184), .B(n_134), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_188), .A2(n_140), .B1(n_152), .B2(n_145), .Y(n_196) );
BUFx12f_ASAP7_75t_L g197 ( .A(n_172), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_165), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_158), .A2(n_152), .B(n_145), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_184), .B(n_134), .Y(n_202) );
NAND2xp33_ASAP7_75t_L g203 ( .A(n_157), .B(n_134), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_183), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_183), .B(n_145), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_167), .B(n_118), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_159), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g209 ( .A1(n_188), .A2(n_72), .B1(n_117), .B2(n_83), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_159), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_159), .Y(n_211) );
BUFx12f_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_157), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_159), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_169), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_187), .B(n_108), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_187), .B(n_83), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_181), .B(n_89), .Y(n_219) );
AOI22xp33_ASAP7_75t_L g220 ( .A1(n_172), .A2(n_72), .B1(n_97), .B2(n_88), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_157), .Y(n_221) );
NOR2xp33_ASAP7_75t_R g222 ( .A(n_175), .B(n_91), .Y(n_222) );
INVx1_ASAP7_75t_SL g223 ( .A(n_157), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_182), .B(n_86), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_216), .Y(n_225) );
OR2x2_ASAP7_75t_L g226 ( .A(n_195), .B(n_158), .Y(n_226) );
AOI221xp5_ASAP7_75t_L g227 ( .A1(n_206), .A2(n_171), .B1(n_167), .B2(n_182), .C(n_189), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_208), .Y(n_228) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_216), .A2(n_185), .B(n_169), .Y(n_229) );
OR2x2_ASAP7_75t_L g230 ( .A(n_195), .B(n_161), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_205), .A2(n_171), .B1(n_182), .B2(n_161), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_198), .Y(n_232) );
INVx3_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
NAND3xp33_ASAP7_75t_SL g234 ( .A(n_222), .B(n_175), .C(n_199), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_191), .A2(n_181), .B(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_198), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_202), .A2(n_189), .B1(n_174), .B2(n_164), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_201), .B(n_164), .Y(n_238) );
NAND4xp25_ASAP7_75t_L g239 ( .A(n_209), .B(n_86), .C(n_97), .D(n_88), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_196), .A2(n_174), .B1(n_164), .B2(n_170), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g241 ( .A1(n_197), .A2(n_175), .B1(n_164), .B2(n_174), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_197), .B(n_160), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_214), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_207), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_202), .B(n_170), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_205), .A2(n_162), .B1(n_163), .B2(n_174), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_205), .B(n_170), .Y(n_247) );
BUFx2_ASAP7_75t_L g248 ( .A(n_197), .Y(n_248) );
NAND2xp33_ASAP7_75t_R g249 ( .A(n_193), .B(n_186), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_205), .B(n_173), .Y(n_250) );
AOI21xp33_ASAP7_75t_L g251 ( .A1(n_196), .A2(n_164), .B(n_174), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_193), .A2(n_162), .B1(n_163), .B2(n_173), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_225), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g254 ( .A1(n_235), .A2(n_194), .B(n_191), .Y(n_254) );
AOI22xp33_ASAP7_75t_SL g255 ( .A1(n_248), .A2(n_212), .B1(n_224), .B2(n_203), .Y(n_255) );
INVxp67_ASAP7_75t_SL g256 ( .A(n_245), .Y(n_256) );
INVx3_ASAP7_75t_L g257 ( .A(n_238), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_245), .B(n_217), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_227), .A2(n_209), .B1(n_224), .B2(n_217), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_251), .A2(n_200), .B(n_194), .C(n_218), .Y(n_260) );
BUFx12f_ASAP7_75t_L g261 ( .A(n_248), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_226), .B(n_230), .Y(n_262) );
AOI222xp33_ASAP7_75t_L g263 ( .A1(n_231), .A2(n_224), .B1(n_218), .B2(n_212), .C1(n_220), .C2(n_193), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_225), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_226), .B(n_201), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_228), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_230), .B(n_201), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g269 ( .A1(n_239), .A2(n_224), .B1(n_200), .B2(n_212), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_247), .A2(n_193), .B1(n_204), .B2(n_215), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_232), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_232), .Y(n_272) );
OAI22xp33_ASAP7_75t_L g273 ( .A1(n_237), .A2(n_223), .B1(n_213), .B2(n_208), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_236), .Y(n_274) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_229), .A2(n_219), .B(n_192), .Y(n_275) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_241), .A2(n_186), .B1(n_93), .B2(n_77), .C(n_81), .Y(n_276) );
OAI33xp33_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_77), .A3(n_81), .B1(n_107), .B2(n_82), .B3(n_106), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_257), .B(n_233), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_269), .A2(n_234), .B1(n_250), .B2(n_247), .C(n_236), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_265), .Y(n_281) );
NAND4xp25_ASAP7_75t_L g282 ( .A(n_269), .B(n_249), .C(n_87), .D(n_107), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_265), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_271), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_271), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_257), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_272), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g289 ( .A(n_257), .B(n_233), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_272), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_262), .B(n_250), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_256), .B(n_242), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_263), .A2(n_240), .B1(n_246), .B2(n_233), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_262), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_262), .Y(n_296) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_276), .A2(n_243), .B(n_101), .C(n_106), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_274), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_284), .B(n_256), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_292), .B(n_261), .Y(n_303) );
AOI21xp33_ASAP7_75t_L g304 ( .A1(n_292), .A2(n_263), .B(n_273), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_294), .B(n_266), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_296), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_284), .Y(n_308) );
NOR3xp33_ASAP7_75t_L g309 ( .A(n_282), .B(n_276), .C(n_255), .Y(n_309) );
INVx1_ASAP7_75t_SL g310 ( .A(n_278), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_285), .B(n_258), .Y(n_311) );
NOR3xp33_ASAP7_75t_SL g312 ( .A(n_297), .B(n_243), .C(n_260), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_285), .B(n_258), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_291), .B(n_266), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_291), .B(n_266), .Y(n_316) );
OAI31xp33_ASAP7_75t_L g317 ( .A1(n_293), .A2(n_268), .A3(n_258), .B(n_273), .Y(n_317) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_283), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_280), .B(n_255), .C(n_259), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g321 ( .A1(n_277), .A2(n_259), .B1(n_254), .B2(n_100), .C(n_98), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_286), .B(n_268), .Y(n_322) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_287), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_268), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_288), .B(n_265), .Y(n_326) );
AOI211x1_ASAP7_75t_L g327 ( .A1(n_290), .A2(n_82), .B(n_99), .C(n_254), .Y(n_327) );
OAI33xp33_ASAP7_75t_L g328 ( .A1(n_290), .A2(n_123), .A3(n_112), .B1(n_127), .B2(n_120), .B3(n_109), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_299), .B(n_298), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_307), .B(n_295), .Y(n_331) );
OAI332xp33_ASAP7_75t_L g332 ( .A1(n_311), .A2(n_298), .A3(n_295), .B1(n_78), .B2(n_127), .B3(n_123), .C1(n_122), .C2(n_120), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_315), .B(n_287), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_299), .B(n_300), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_308), .B(n_287), .Y(n_336) );
CKINVDCx8_ASAP7_75t_R g337 ( .A(n_309), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_318), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_316), .B(n_278), .Y(n_339) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_320), .A2(n_270), .B1(n_278), .B2(n_244), .C(n_127), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_303), .B(n_257), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_324), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_306), .B(n_278), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_325), .B(n_267), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_317), .A2(n_261), .B1(n_270), .B2(n_244), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_301), .Y(n_349) );
NAND2xp33_ASAP7_75t_R g350 ( .A(n_312), .B(n_267), .Y(n_350) );
NAND2xp33_ASAP7_75t_SL g351 ( .A(n_322), .B(n_267), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_322), .Y(n_352) );
NOR4xp25_ASAP7_75t_SL g353 ( .A(n_304), .B(n_261), .C(n_103), .D(n_92), .Y(n_353) );
OAI31xp33_ASAP7_75t_L g354 ( .A1(n_317), .A2(n_289), .A3(n_238), .B(n_252), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_325), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_321), .B(n_109), .C(n_112), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_311), .B(n_289), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_314), .B(n_289), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_314), .B(n_1), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_326), .B(n_2), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_302), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_304), .B(n_305), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_310), .B(n_305), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_305), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_319), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_310), .B(n_2), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_319), .B(n_275), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_319), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_323), .A2(n_238), .B1(n_120), .B2(n_122), .C(n_123), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_347), .A2(n_313), .B1(n_328), .B2(n_275), .Y(n_371) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_350), .A2(n_313), .B1(n_327), .B2(n_223), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_338), .B(n_313), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_338), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_347), .A2(n_327), .B1(n_221), .B2(n_192), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_337), .A2(n_341), .B1(n_340), .B2(n_359), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_341), .A2(n_192), .B1(n_221), .B2(n_208), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_355), .B(n_3), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_331), .B(n_3), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_360), .A2(n_135), .B1(n_143), .B2(n_141), .C(n_144), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_352), .B(n_356), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_330), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_348), .B(n_4), .Y(n_385) );
NOR2xp33_ASAP7_75t_SL g386 ( .A(n_354), .B(n_213), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_349), .B(n_4), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_351), .B(n_275), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_345), .Y(n_389) );
OAI322xp33_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_135), .A3(n_143), .B1(n_141), .B2(n_144), .C1(n_146), .C2(n_147), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_332), .A2(n_229), .B(n_213), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_329), .B(n_5), .Y(n_392) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_361), .A2(n_141), .B1(n_144), .B2(n_146), .C(n_147), .Y(n_393) );
INVxp67_ASAP7_75t_SL g394 ( .A(n_369), .Y(n_394) );
OAI32xp33_ASAP7_75t_L g395 ( .A1(n_350), .A2(n_5), .A3(n_7), .B1(n_9), .B2(n_10), .Y(n_395) );
AOI221x1_ASAP7_75t_L g396 ( .A1(n_335), .A2(n_146), .B1(n_147), .B2(n_11), .C(n_12), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_364), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_346), .B(n_7), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_358), .A2(n_339), .B1(n_333), .B2(n_367), .Y(n_399) );
NAND2xp33_ASAP7_75t_L g400 ( .A(n_336), .B(n_9), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_329), .B(n_11), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_343), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_344), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_336), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_370), .A2(n_13), .B(n_14), .C(n_15), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_362), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_366), .B(n_14), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_364), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_342), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_365), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_365), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_368), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g413 ( .A1(n_357), .A2(n_147), .B1(n_138), .B2(n_210), .C(n_211), .Y(n_413) );
OAI31xp33_ASAP7_75t_L g414 ( .A1(n_368), .A2(n_15), .A3(n_16), .B(n_17), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_353), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_355), .B(n_17), .Y(n_416) );
XNOR2x1_ASAP7_75t_L g417 ( .A(n_339), .B(n_18), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
AOI311xp33_ASAP7_75t_L g419 ( .A1(n_399), .A2(n_18), .A3(n_19), .B(n_20), .C(n_21), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_412), .B(n_22), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_375), .B(n_156), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_383), .B(n_404), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_397), .B(n_138), .Y(n_423) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_394), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_397), .B(n_138), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_402), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_403), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_389), .B(n_138), .Y(n_430) );
HAxp5_ASAP7_75t_SL g431 ( .A(n_415), .B(n_25), .CON(n_431), .SN(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_412), .B(n_26), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_401), .B(n_138), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_374), .Y(n_435) );
OAI22xp33_ASAP7_75t_L g436 ( .A1(n_386), .A2(n_221), .B1(n_177), .B2(n_179), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_400), .A2(n_372), .B(n_388), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_384), .B(n_409), .Y(n_438) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_417), .A2(n_177), .B(n_176), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_392), .B(n_27), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_373), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_378), .A2(n_173), .B1(n_176), .B2(n_190), .Y(n_442) );
AOI211x1_ASAP7_75t_L g443 ( .A1(n_395), .A2(n_32), .B(n_33), .C(n_38), .Y(n_443) );
AOI21xp33_ASAP7_75t_L g444 ( .A1(n_381), .A2(n_40), .B(n_41), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_411), .Y(n_446) );
NOR2xp33_ASAP7_75t_R g447 ( .A(n_398), .B(n_416), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_407), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_385), .B(n_43), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_387), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_372), .A2(n_190), .B1(n_180), .B2(n_178), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_437), .A2(n_380), .B1(n_376), .B2(n_379), .Y(n_452) );
NOR2x1p5_ASAP7_75t_L g453 ( .A(n_424), .B(n_414), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_439), .A2(n_371), .B1(n_405), .B2(n_391), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_424), .B(n_396), .Y(n_455) );
OAI21xp5_ASAP7_75t_L g456 ( .A1(n_420), .A2(n_451), .B(n_442), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g457 ( .A1(n_420), .A2(n_413), .B1(n_382), .B2(n_393), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_429), .Y(n_458) );
XNOR2xp5_ASAP7_75t_L g459 ( .A(n_422), .B(n_44), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_433), .B(n_47), .Y(n_460) );
OAI22xp33_ASAP7_75t_SL g461 ( .A1(n_450), .A2(n_390), .B1(n_52), .B2(n_53), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_448), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_441), .A2(n_177), .B1(n_179), .B2(n_168), .Y(n_463) );
OAI21xp33_ASAP7_75t_L g464 ( .A1(n_447), .A2(n_179), .B(n_57), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_428), .A2(n_177), .B1(n_168), .B2(n_60), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_418), .B(n_56), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_432), .B(n_168), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_438), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_449), .A2(n_63), .B(n_64), .C(n_65), .Y(n_472) );
INVxp67_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
AOI322xp5_ASAP7_75t_L g474 ( .A1(n_452), .A2(n_419), .A3(n_432), .B1(n_445), .B2(n_446), .C1(n_435), .C2(n_447), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_471), .A2(n_443), .B1(n_444), .B2(n_430), .C(n_434), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_470), .Y(n_476) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_454), .B(n_440), .C(n_421), .Y(n_477) );
NOR2xp33_ASAP7_75t_R g478 ( .A(n_459), .B(n_431), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_453), .A2(n_432), .B1(n_436), .B2(n_431), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_455), .B(n_436), .Y(n_480) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_467), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_458), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_466), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_454), .B(n_163), .C(n_168), .D(n_160), .Y(n_484) );
NAND3xp33_ASAP7_75t_SL g485 ( .A(n_472), .B(n_168), .C(n_160), .Y(n_485) );
OAI31xp33_ASAP7_75t_L g486 ( .A1(n_461), .A2(n_160), .A3(n_455), .B(n_469), .Y(n_486) );
NAND4xp25_ASAP7_75t_L g487 ( .A(n_456), .B(n_160), .C(n_457), .D(n_468), .Y(n_487) );
NAND4xp25_ASAP7_75t_L g488 ( .A(n_462), .B(n_160), .C(n_465), .D(n_460), .Y(n_488) );
NOR4xp25_ASAP7_75t_L g489 ( .A(n_463), .B(n_419), .C(n_450), .D(n_454), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_471), .A2(n_473), .B1(n_454), .B2(n_450), .C(n_467), .Y(n_490) );
OAI311xp33_ASAP7_75t_L g491 ( .A1(n_464), .A2(n_439), .A3(n_456), .B1(n_381), .C1(n_347), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_485), .Y(n_492) );
XNOR2xp5_ASAP7_75t_L g493 ( .A(n_479), .B(n_489), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_481), .B(n_490), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_480), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_482), .Y(n_496) );
NOR4xp25_ASAP7_75t_L g497 ( .A(n_493), .B(n_491), .C(n_487), .D(n_479), .Y(n_497) );
OAI211xp5_ASAP7_75t_L g498 ( .A1(n_495), .A2(n_478), .B(n_474), .C(n_486), .Y(n_498) );
OR3x2_ASAP7_75t_L g499 ( .A(n_493), .B(n_484), .C(n_488), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_498), .A2(n_494), .B1(n_477), .B2(n_492), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_499), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_501), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_500), .B(n_497), .Y(n_503) );
AOI322xp5_ASAP7_75t_L g504 ( .A1(n_502), .A2(n_494), .A3(n_492), .B1(n_496), .B2(n_483), .C1(n_475), .C2(n_476), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_504), .A2(n_503), .B(n_492), .Y(n_505) );
endmodule