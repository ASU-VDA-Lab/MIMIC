module fake_netlist_6_3682_n_1647 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1647);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1647;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx10_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_57),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_19),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_79),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_19),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_103),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_37),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_96),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_109),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_45),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_81),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_51),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_10),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_56),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_87),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_36),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_69),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_77),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_37),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_21),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_52),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_3),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_84),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_53),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_68),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_46),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_66),
.Y(n_191)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_107),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_15),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_31),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_127),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_58),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_62),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_36),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_7),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_48),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_92),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_49),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_60),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_90),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_9),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_31),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_22),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_35),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_137),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_78),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_153),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_88),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_123),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_102),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_130),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_9),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_113),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_8),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_59),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_141),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_145),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_41),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_65),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_116),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_89),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_148),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_95),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_63),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_5),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_122),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_40),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_26),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_124),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_16),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_149),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_39),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_93),
.Y(n_245)
);

CKINVDCx11_ASAP7_75t_R g246 ( 
.A(n_34),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_117),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_14),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_67),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_146),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_43),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_111),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_15),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_71),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_1),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_50),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_4),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_73),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_82),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_133),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

BUFx8_ASAP7_75t_SL g263 ( 
.A(n_150),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_132),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_125),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_112),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_97),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_39),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_47),
.Y(n_270)
);

BUFx2_ASAP7_75t_SL g271 ( 
.A(n_20),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_131),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_24),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_100),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_75),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_42),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_33),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_76),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_3),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_26),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_54),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_21),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_6),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_144),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_104),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_64),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_0),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_83),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_94),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_22),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_147),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_129),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_25),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_139),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_29),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_55),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_86),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_140),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_101),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_17),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_5),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

INVxp33_ASAP7_75t_SL g307 ( 
.A(n_200),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_293),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_157),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_263),
.Y(n_313)
);

INVx4_ASAP7_75t_R g314 ( 
.A(n_226),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_246),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_267),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_199),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_194),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_203),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_183),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_186),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_188),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_194),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_242),
.Y(n_326)
);

INVxp33_ASAP7_75t_SL g327 ( 
.A(n_158),
.Y(n_327)
);

INVxp33_ASAP7_75t_SL g328 ( 
.A(n_158),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_242),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g330 ( 
.A(n_226),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_302),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_189),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_163),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_288),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_191),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_175),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_163),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_195),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_196),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_197),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_202),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_257),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_175),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_206),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_155),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_257),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_209),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_214),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

INVxp33_ASAP7_75t_SL g353 ( 
.A(n_172),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_216),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_302),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_182),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_218),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_217),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_235),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_172),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_219),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_220),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_229),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_253),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_221),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_235),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_279),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_212),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_295),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_254),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_227),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_181),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_175),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_228),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_181),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_254),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_321),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_235),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_306),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_222),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_367),
.B(n_222),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_308),
.B(n_275),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_310),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_330),
.B(n_156),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_346),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_331),
.B(n_165),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_311),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_346),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_336),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_311),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_375),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_L g406 ( 
.A(n_322),
.B(n_284),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_375),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_R g408 ( 
.A(n_307),
.B(n_304),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_355),
.B(n_315),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_370),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_375),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_315),
.B(n_159),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_352),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_333),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_249),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_372),
.A2(n_169),
.B(n_168),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_379),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_378),
.B(n_159),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_378),
.B(n_171),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_324),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

INVx6_ASAP7_75t_L g428 ( 
.A(n_375),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_342),
.B(n_161),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_319),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_161),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_319),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_325),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_325),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_326),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_374),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_326),
.B(n_178),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_318),
.A2(n_283),
.B1(n_177),
.B2(n_239),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_320),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_329),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_329),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_332),
.B(n_154),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_348),
.B(n_162),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_337),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_337),
.B(n_185),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_356),
.Y(n_448)
);

OR2x6_ASAP7_75t_L g449 ( 
.A(n_409),
.B(n_192),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_409),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_385),
.B(n_335),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_405),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_385),
.B(n_340),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_SL g458 ( 
.A1(n_410),
.A2(n_317),
.B1(n_291),
.B2(n_334),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_410),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_341),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_394),
.B(n_343),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_444),
.B(n_344),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_385),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g471 ( 
.A(n_440),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_381),
.B(n_347),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_400),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_383),
.Y(n_476)
);

AO22x2_ASAP7_75t_L g477 ( 
.A1(n_385),
.A2(n_309),
.B1(n_271),
.B2(n_269),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_426),
.B(n_350),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_386),
.B(n_338),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_430),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_391),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_415),
.B(n_276),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_430),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_387),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_430),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_386),
.B(n_338),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_386),
.B(n_351),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_430),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_382),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

NAND3xp33_ASAP7_75t_L g497 ( 
.A(n_396),
.B(n_357),
.C(n_356),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_415),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_430),
.Y(n_499)
);

INVx8_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_441),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_387),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_387),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_427),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_444),
.B(n_354),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_387),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_427),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_387),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_432),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_432),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_425),
.Y(n_513)
);

NAND3xp33_ASAP7_75t_L g514 ( 
.A(n_396),
.B(n_358),
.C(n_357),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_432),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_425),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_448),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_448),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_R g519 ( 
.A(n_437),
.B(n_327),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_L g520 ( 
.A(n_396),
.B(n_364),
.C(n_358),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_420),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

AND3x2_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_349),
.C(n_345),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_383),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_424),
.B(n_359),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_433),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_424),
.B(n_362),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_383),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_383),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_433),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_388),
.Y(n_536)
);

CKINVDCx6p67_ASAP7_75t_R g537 ( 
.A(n_440),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_423),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_412),
.B(n_363),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_408),
.B(n_316),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_438),
.Y(n_544)
);

INVxp33_ASAP7_75t_SL g545 ( 
.A(n_439),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_412),
.B(n_366),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_434),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_438),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_438),
.Y(n_549)
);

OR2x6_ASAP7_75t_L g550 ( 
.A(n_421),
.B(n_190),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_198),
.Y(n_551)
);

INVx11_ASAP7_75t_L g552 ( 
.A(n_382),
.Y(n_552)
);

CKINVDCx6p67_ASAP7_75t_R g553 ( 
.A(n_434),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_406),
.B(n_373),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_422),
.Y(n_557)
);

OA22x2_ASAP7_75t_L g558 ( 
.A1(n_422),
.A2(n_345),
.B1(n_349),
.B2(n_369),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_433),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_442),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_421),
.B(n_376),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_SL g562 ( 
.A(n_429),
.B(n_284),
.C(n_296),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_388),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_429),
.B(n_328),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_442),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_439),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_431),
.B(n_353),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_442),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_431),
.B(n_313),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_445),
.B(n_154),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_445),
.B(n_364),
.Y(n_573)
);

AND3x2_ASAP7_75t_L g574 ( 
.A(n_436),
.B(n_213),
.C(n_303),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_393),
.B(n_238),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_388),
.Y(n_576)
);

INVx4_ASAP7_75t_L g577 ( 
.A(n_382),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_388),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_442),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_442),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_419),
.A2(n_175),
.B1(n_369),
.B2(n_368),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_389),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_389),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_419),
.A2(n_371),
.B1(n_368),
.B2(n_365),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_389),
.Y(n_587)
);

HB1xp67_ASAP7_75t_L g588 ( 
.A(n_408),
.Y(n_588)
);

INVxp67_ASAP7_75t_SL g589 ( 
.A(n_393),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_435),
.B(n_371),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_SL g591 ( 
.A1(n_419),
.A2(n_160),
.B1(n_294),
.B2(n_301),
.Y(n_591)
);

CKINVDCx6p67_ASAP7_75t_R g592 ( 
.A(n_382),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_392),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_392),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_392),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_399),
.Y(n_596)
);

NAND2xp33_ASAP7_75t_SL g597 ( 
.A(n_454),
.B(n_285),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_505),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_513),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_454),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_162),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_469),
.B(n_435),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_584),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_467),
.B(n_164),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_469),
.B(n_435),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_544),
.A2(n_234),
.B1(n_205),
.B2(n_207),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_505),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_493),
.B(n_164),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_451),
.A2(n_417),
.B1(n_252),
.B2(n_256),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_573),
.B(n_435),
.Y(n_610)
);

INVxp67_ASAP7_75t_SL g611 ( 
.A(n_536),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_573),
.B(n_443),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_584),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_452),
.A2(n_417),
.B1(n_245),
.B2(n_274),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_544),
.B(n_443),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_548),
.B(n_443),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_457),
.B(n_215),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_562),
.B(n_365),
.C(n_225),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_548),
.B(n_443),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_486),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_557),
.B(n_224),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_516),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_549),
.B(n_393),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_555),
.B(n_166),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_488),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_471),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_465),
.B(n_154),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_588),
.B(n_232),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_549),
.B(n_393),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_L g633 ( 
.A1(n_557),
.A2(n_418),
.B(n_399),
.Y(n_633)
);

NOR2x1p5_ASAP7_75t_L g634 ( 
.A(n_537),
.B(n_285),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_498),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_554),
.B(n_395),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_585),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_561),
.B(n_166),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_554),
.B(n_395),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_537),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_556),
.B(n_395),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_564),
.A2(n_260),
.B1(n_241),
.B2(n_243),
.Y(n_642)
);

AND2x2_ASAP7_75t_SL g643 ( 
.A(n_542),
.B(n_230),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_565),
.B(n_231),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_517),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_546),
.B(n_167),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_556),
.B(n_395),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_517),
.Y(n_648)
);

NAND2xp33_ASAP7_75t_SL g649 ( 
.A(n_498),
.B(n_289),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_518),
.B(n_236),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_553),
.B(n_289),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_547),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_518),
.Y(n_653)
);

O2A1O1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_497),
.A2(n_261),
.B(n_259),
.C(n_258),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_568),
.B(n_167),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_483),
.B(n_398),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_486),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_485),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_483),
.B(n_398),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_565),
.B(n_266),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_571),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_532),
.B(n_204),
.C(n_184),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_593),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_571),
.B(n_287),
.Y(n_664)
);

NOR3xp33_ASAP7_75t_L g665 ( 
.A(n_458),
.B(n_208),
.C(n_262),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_501),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_500),
.B(n_247),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_450),
.B(n_495),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_491),
.B(n_522),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_503),
.Y(n_670)
);

NAND2x1p5_ASAP7_75t_L g671 ( 
.A(n_450),
.B(n_290),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_491),
.B(n_398),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_522),
.B(n_398),
.Y(n_673)
);

A2O1A1Ixp33_ASAP7_75t_L g674 ( 
.A1(n_503),
.A2(n_446),
.B(n_436),
.C(n_416),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_558),
.A2(n_382),
.B1(n_304),
.B2(n_292),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_526),
.B(n_403),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_593),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_526),
.B(n_403),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_558),
.A2(n_382),
.B1(n_292),
.B2(n_299),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_466),
.B(n_170),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_529),
.B(n_403),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_529),
.B(n_403),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_527),
.B(n_170),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_547),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_558),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_596),
.Y(n_686)
);

O2A1O1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_497),
.A2(n_446),
.B(n_436),
.C(n_416),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_SL g688 ( 
.A(n_460),
.B(n_388),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_540),
.B(n_507),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_540),
.B(n_411),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_510),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_SL g692 ( 
.A(n_506),
.B(n_296),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_572),
.B(n_173),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_551),
.A2(n_418),
.B(n_411),
.C(n_414),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_L g695 ( 
.A(n_500),
.B(n_250),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_453),
.B(n_411),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_453),
.B(n_418),
.Y(n_697)
);

BUFx6f_ASAP7_75t_SL g698 ( 
.A(n_449),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_519),
.Y(n_699)
);

NOR2x1p5_ASAP7_75t_L g700 ( 
.A(n_553),
.B(n_297),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_455),
.B(n_446),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_500),
.B(n_251),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_551),
.B(n_173),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_550),
.B(n_174),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_587),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_455),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_514),
.B(n_174),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_456),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_587),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_504),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_464),
.Y(n_711)
);

NAND2x1p5_ASAP7_75t_L g712 ( 
.A(n_450),
.B(n_388),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_464),
.B(n_399),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_550),
.B(n_176),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_550),
.B(n_176),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_514),
.B(n_237),
.C(n_281),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_500),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_449),
.Y(n_718)
);

INVx3_ASAP7_75t_L g719 ( 
.A(n_456),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_509),
.B(n_297),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_468),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_468),
.Y(n_722)
);

O2A1O1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_520),
.A2(n_414),
.B(n_413),
.C(n_314),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_543),
.B(n_193),
.C(n_201),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_550),
.B(n_179),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_495),
.B(n_264),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_495),
.B(n_265),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_470),
.B(n_413),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_477),
.A2(n_299),
.B1(n_160),
.B2(n_244),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_R g730 ( 
.A(n_524),
.B(n_592),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_577),
.B(n_270),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_550),
.A2(n_233),
.B1(n_223),
.B2(n_280),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_577),
.B(n_272),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_577),
.B(n_278),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_475),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_594),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_500),
.B(n_298),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_594),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_475),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_536),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_595),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_551),
.B(n_179),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_520),
.B(n_298),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_478),
.B(n_414),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_595),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_478),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_551),
.B(n_180),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_460),
.B(n_180),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_460),
.B(n_300),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_SL g750 ( 
.A(n_570),
.B(n_240),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_461),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_482),
.B(n_407),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_449),
.B(n_286),
.Y(n_753)
);

OAI221xp5_ASAP7_75t_L g754 ( 
.A1(n_591),
.A2(n_248),
.B1(n_273),
.B2(n_300),
.C(n_282),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_474),
.B(n_282),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_567),
.B(n_286),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_601),
.B(n_449),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_658),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_618),
.Y(n_759)
);

INVx5_ASAP7_75t_L g760 ( 
.A(n_717),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_710),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_626),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_607),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_601),
.B(n_449),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_600),
.Y(n_765)
);

INVx2_ASAP7_75t_SL g766 ( 
.A(n_635),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_R g767 ( 
.A(n_699),
.B(n_592),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_626),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_685),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_628),
.Y(n_770)
);

A2O1A1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_638),
.A2(n_590),
.B(n_582),
.C(n_575),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_638),
.B(n_590),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_643),
.A2(n_481),
.B1(n_589),
.B2(n_477),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_607),
.Y(n_774)
);

AND2x4_ASAP7_75t_SL g775 ( 
.A(n_666),
.B(n_607),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_628),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_621),
.B(n_545),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_646),
.B(n_461),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_652),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_646),
.B(n_473),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_730),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_708),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_SL g783 ( 
.A1(n_657),
.A2(n_545),
.B1(n_729),
.B2(n_655),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_661),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_643),
.B(n_473),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_653),
.B(n_479),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_685),
.A2(n_477),
.B1(n_586),
.B2(n_479),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_670),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_756),
.B(n_480),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_610),
.B(n_480),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_691),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_684),
.B(n_462),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_598),
.B(n_484),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_720),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_717),
.B(n_460),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_627),
.B(n_462),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_640),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_607),
.B(n_477),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_612),
.A2(n_583),
.B(n_581),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_598),
.B(n_484),
.Y(n_800)
);

CKINVDCx8_ASAP7_75t_R g801 ( 
.A(n_703),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_655),
.B(n_187),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_599),
.B(n_487),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_669),
.B(n_462),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_717),
.B(n_460),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_719),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_751),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_623),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_603),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_613),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_683),
.B(n_574),
.C(n_581),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_630),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_604),
.B(n_472),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_645),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_606),
.A2(n_301),
.B1(n_294),
.B2(n_187),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_648),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_650),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_650),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_706),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_637),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_680),
.A2(n_583),
.B1(n_580),
.B2(n_579),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_656),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_703),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_711),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_663),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_721),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_722),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_717),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_735),
.B(n_487),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_677),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_739),
.B(n_476),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_730),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_606),
.A2(n_301),
.B1(n_294),
.B2(n_187),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_686),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_729),
.A2(n_580),
.B1(n_579),
.B2(n_489),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_671),
.B(n_460),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_680),
.A2(n_531),
.B1(n_492),
.B2(n_569),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_742),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_740),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_671),
.B(n_536),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_746),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_659),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_705),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_675),
.A2(n_492),
.B1(n_494),
.B2(n_569),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_718),
.B(n_489),
.Y(n_845)
);

CKINVDCx16_ASAP7_75t_R g846 ( 
.A(n_698),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_689),
.B(n_476),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_672),
.B(n_496),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_624),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_615),
.B(n_496),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_632),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_683),
.B(n_496),
.Y(n_852)
);

AOI22x1_ASAP7_75t_L g853 ( 
.A1(n_709),
.A2(n_528),
.B1(n_511),
.B2(n_566),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_704),
.A2(n_528),
.B1(n_511),
.B2(n_566),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_616),
.B(n_525),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_620),
.B(n_525),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_631),
.B(n_525),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_736),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_636),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_738),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_639),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_742),
.B(n_490),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_741),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_675),
.A2(n_531),
.B1(n_508),
.B2(n_512),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_718),
.B(n_490),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_747),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_641),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_745),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_732),
.B(n_499),
.C(n_494),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_647),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_740),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_617),
.B(n_679),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_697),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_679),
.B(n_539),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_R g875 ( 
.A(n_750),
.B(n_120),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_747),
.B(n_629),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_694),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_740),
.Y(n_878)
);

AND2x6_ASAP7_75t_SL g879 ( 
.A(n_753),
.B(n_2),
.Y(n_879)
);

AND2x4_ASAP7_75t_L g880 ( 
.A(n_716),
.B(n_535),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_692),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_732),
.B(n_704),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_625),
.B(n_533),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_714),
.B(n_576),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_701),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_714),
.B(n_576),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_688),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_715),
.B(n_563),
.Y(n_888)
);

BUFx4f_ASAP7_75t_L g889 ( 
.A(n_698),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_634),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_673),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_715),
.B(n_563),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_725),
.B(n_563),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_676),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_602),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_678),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_725),
.B(n_534),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_753),
.B(n_534),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_611),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_608),
.B(n_499),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_665),
.B(n_508),
.Y(n_901)
);

BUFx12f_ASAP7_75t_SL g902 ( 
.A(n_597),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_681),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_605),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_622),
.B(n_578),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_622),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_644),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_712),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_649),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_609),
.B(n_530),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_752),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_754),
.A2(n_530),
.B1(n_560),
.B2(n_559),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_682),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_690),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_651),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_723),
.B(n_614),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_660),
.B(n_578),
.Y(n_917)
);

NOR2x1_ASAP7_75t_L g918 ( 
.A(n_662),
.B(n_755),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_619),
.A2(n_664),
.B1(n_707),
.B2(n_743),
.Y(n_919)
);

NAND2x1p5_ASAP7_75t_L g920 ( 
.A(n_668),
.B(n_535),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_696),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_693),
.B(n_578),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_712),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_664),
.B(n_578),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_713),
.B(n_578),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_724),
.B(n_4),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_668),
.B(n_521),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_882),
.A2(n_733),
.B1(n_726),
.B2(n_727),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_882),
.A2(n_734),
.B1(n_726),
.B2(n_731),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_762),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_761),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_785),
.A2(n_757),
.B(n_764),
.C(n_872),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_763),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_769),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_836),
.A2(n_695),
.B(n_702),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_758),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_772),
.A2(n_731),
.B1(n_727),
.B2(n_734),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_R g938 ( 
.A(n_781),
.B(n_737),
.Y(n_938)
);

INVx6_ASAP7_75t_L g939 ( 
.A(n_797),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_899),
.A2(n_733),
.B1(n_633),
.B2(n_642),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_779),
.Y(n_941)
);

INVx4_ASAP7_75t_L g942 ( 
.A(n_763),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_802),
.A2(n_926),
.B(n_777),
.C(n_785),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_803),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_840),
.A2(n_667),
.B(n_536),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_777),
.B(n_749),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_763),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_916),
.A2(n_674),
.B(n_749),
.C(n_748),
.Y(n_948)
);

O2A1O1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_906),
.A2(n_907),
.B(n_778),
.C(n_780),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_760),
.A2(n_536),
.B(n_728),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_R g951 ( 
.A(n_832),
.B(n_744),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_774),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_822),
.B(n_654),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_842),
.B(n_687),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_842),
.B(n_885),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_760),
.A2(n_388),
.B(n_402),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_773),
.A2(n_919),
.B(n_888),
.C(n_852),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_760),
.A2(n_790),
.B(n_899),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_774),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_852),
.A2(n_552),
.B1(n_700),
.B2(n_541),
.Y(n_960)
);

BUFx2_ASAP7_75t_L g961 ( 
.A(n_759),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_775),
.Y(n_962)
);

OAI22x1_ASAP7_75t_L g963 ( 
.A1(n_866),
.A2(n_6),
.B1(n_7),
.B2(n_10),
.Y(n_963)
);

AOI33xp33_ASAP7_75t_L g964 ( 
.A1(n_815),
.A2(n_515),
.A3(n_523),
.B1(n_538),
.B2(n_539),
.B3(n_17),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_873),
.B(n_515),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_760),
.A2(n_771),
.B(n_847),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_888),
.A2(n_538),
.B1(n_314),
.B2(n_428),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_803),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_829),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_769),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_783),
.B(n_11),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_794),
.B(n_11),
.Y(n_972)
);

INVx1_ASAP7_75t_SL g973 ( 
.A(n_765),
.Y(n_973)
);

AO21x1_ASAP7_75t_L g974 ( 
.A1(n_916),
.A2(n_13),
.B(n_14),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_798),
.B(n_428),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_887),
.A2(n_407),
.B(n_402),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_910),
.A2(n_152),
.B(n_151),
.C(n_142),
.Y(n_977)
);

AO22x1_ASAP7_75t_L g978 ( 
.A1(n_876),
.A2(n_13),
.B1(n_16),
.B2(n_20),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_784),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_849),
.B(n_23),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_851),
.B(n_23),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_887),
.A2(n_407),
.B(n_402),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_887),
.A2(n_407),
.B(n_402),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_923),
.A2(n_428),
.B1(n_407),
.B2(n_402),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_887),
.A2(n_925),
.B(n_923),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_829),
.Y(n_986)
);

CKINVDCx8_ASAP7_75t_R g987 ( 
.A(n_846),
.Y(n_987)
);

AND2x2_ASAP7_75t_SL g988 ( 
.A(n_815),
.B(n_24),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_923),
.A2(n_402),
.B(n_428),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_SL g990 ( 
.A(n_801),
.B(n_428),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_789),
.B(n_135),
.Y(n_991)
);

O2A1O1Ixp5_ASAP7_75t_L g992 ( 
.A1(n_910),
.A2(n_126),
.B(n_114),
.C(n_110),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_890),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_866),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_859),
.B(n_25),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_L g996 ( 
.A1(n_874),
.A2(n_106),
.B(n_99),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_857),
.A2(n_91),
.B(n_72),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_861),
.B(n_27),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_898),
.A2(n_61),
.B1(n_28),
.B2(n_29),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_774),
.Y(n_1000)
);

OR2x6_ASAP7_75t_SL g1001 ( 
.A(n_915),
.B(n_27),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_774),
.Y(n_1002)
);

NOR2xp67_ASAP7_75t_L g1003 ( 
.A(n_811),
.B(n_28),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_838),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_788),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_767),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_902),
.B(n_42),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_826),
.B(n_30),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_867),
.B(n_870),
.Y(n_1009)
);

O2A1O1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_906),
.A2(n_30),
.B(n_32),
.C(n_33),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_898),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_786),
.B(n_38),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_786),
.B(n_841),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_907),
.A2(n_41),
.B1(n_919),
.B2(n_893),
.Y(n_1014)
);

OAI22x1_ASAP7_75t_L g1015 ( 
.A1(n_909),
.A2(n_823),
.B1(n_817),
.B2(n_918),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_848),
.A2(n_927),
.B(n_804),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_901),
.A2(n_798),
.B1(n_862),
.B2(n_880),
.Y(n_1017)
);

INVx3_ASAP7_75t_SL g1018 ( 
.A(n_881),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_767),
.B(n_766),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_791),
.B(n_808),
.Y(n_1020)
);

INVx8_ASAP7_75t_L g1021 ( 
.A(n_880),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_818),
.B(n_796),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_814),
.B(n_816),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_798),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_796),
.B(n_819),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_824),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_884),
.A2(n_897),
.B1(n_892),
.B2(n_886),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_828),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_827),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_862),
.B(n_895),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_843),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_839),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_833),
.A2(n_869),
.B(n_874),
.C(n_913),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_891),
.B(n_894),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_858),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_869),
.A2(n_833),
.B1(n_900),
.B2(n_787),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_860),
.B(n_863),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_813),
.A2(n_922),
.B(n_896),
.C(n_914),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_SL g1039 ( 
.A1(n_813),
.A2(n_922),
.B(n_792),
.C(n_912),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_927),
.A2(n_805),
.B(n_795),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_768),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_795),
.A2(n_805),
.B(n_855),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_SL g1043 ( 
.A1(n_879),
.A2(n_787),
.B1(n_776),
.B2(n_770),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_889),
.B(n_868),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_839),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_807),
.B(n_825),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_875),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_903),
.A2(n_865),
.B(n_845),
.C(n_921),
.Y(n_1048)
);

NOR3xp33_ASAP7_75t_L g1049 ( 
.A(n_845),
.B(n_865),
.C(n_883),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_911),
.B(n_895),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_908),
.A2(n_904),
.B1(n_895),
.B2(n_920),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_839),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_839),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_878),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_SL g1055 ( 
.A1(n_792),
.A2(n_912),
.B(n_877),
.C(n_908),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_878),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_895),
.A2(n_904),
.B1(n_782),
.B2(n_806),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_809),
.Y(n_1058)
);

INVx5_ASAP7_75t_L g1059 ( 
.A(n_878),
.Y(n_1059)
);

OAI22x1_ASAP7_75t_L g1060 ( 
.A1(n_854),
.A2(n_821),
.B1(n_837),
.B2(n_889),
.Y(n_1060)
);

NAND2x1p5_ASAP7_75t_L g1061 ( 
.A(n_871),
.B(n_793),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_793),
.B(n_800),
.Y(n_1062)
);

OAI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_835),
.A2(n_875),
.B(n_844),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_850),
.A2(n_856),
.B(n_924),
.Y(n_1064)
);

OAI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_957),
.A2(n_799),
.B(n_844),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1046),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_1044),
.B(n_800),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_931),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_946),
.A2(n_920),
.B1(n_917),
.B2(n_905),
.Y(n_1069)
);

OAI21x1_ASAP7_75t_SL g1070 ( 
.A1(n_974),
.A2(n_835),
.B(n_799),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_979),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1022),
.B(n_810),
.Y(n_1072)
);

AO31x2_ASAP7_75t_L g1073 ( 
.A1(n_937),
.A2(n_831),
.A3(n_820),
.B(n_830),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_955),
.B(n_812),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_1040),
.A2(n_853),
.B(n_864),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_1032),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1009),
.B(n_834),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_1027),
.B(n_940),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1034),
.B(n_1025),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_941),
.Y(n_1080)
);

OAI21x1_ASAP7_75t_L g1081 ( 
.A1(n_1042),
.A2(n_1016),
.B(n_1064),
.Y(n_1081)
);

AO22x2_ASAP7_75t_L g1082 ( 
.A1(n_1014),
.A2(n_1011),
.B1(n_999),
.B2(n_988),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_1021),
.B(n_962),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_985),
.A2(n_1051),
.B(n_950),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_L g1085 ( 
.A1(n_971),
.A2(n_1024),
.B1(n_1012),
.B2(n_1008),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1038),
.A2(n_1039),
.B(n_932),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_1060),
.A2(n_967),
.A3(n_1015),
.B(n_960),
.Y(n_1087)
);

AOI21x1_ASAP7_75t_L g1088 ( 
.A1(n_958),
.A2(n_953),
.B(n_954),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_1004),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_956),
.A2(n_989),
.B(n_965),
.Y(n_1090)
);

OR2x6_ASAP7_75t_L g1091 ( 
.A(n_1021),
.B(n_939),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1036),
.B(n_1026),
.Y(n_1092)
);

OA22x2_ASAP7_75t_L g1093 ( 
.A1(n_963),
.A2(n_1043),
.B1(n_970),
.B2(n_934),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1033),
.A2(n_928),
.B(n_929),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1047),
.B(n_994),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_1006),
.Y(n_1096)
);

NOR4xp25_ASAP7_75t_L g1097 ( 
.A(n_1010),
.B(n_1063),
.C(n_949),
.D(n_964),
.Y(n_1097)
);

AO22x2_ASAP7_75t_L g1098 ( 
.A1(n_996),
.A2(n_981),
.B1(n_980),
.B2(n_995),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1020),
.B(n_1023),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_SL g1100 ( 
.A1(n_972),
.A2(n_1017),
.B(n_1013),
.Y(n_1100)
);

OA21x2_ASAP7_75t_L g1101 ( 
.A1(n_977),
.A2(n_992),
.B(n_1049),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1050),
.B(n_1005),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_1062),
.Y(n_1103)
);

INVxp67_ASAP7_75t_L g1104 ( 
.A(n_961),
.Y(n_1104)
);

INVx3_ASAP7_75t_SL g1105 ( 
.A(n_939),
.Y(n_1105)
);

BUFx12f_ASAP7_75t_L g1106 ( 
.A(n_936),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_951),
.B(n_973),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_1059),
.Y(n_1108)
);

AO22x1_ASAP7_75t_L g1109 ( 
.A1(n_1018),
.A2(n_1029),
.B1(n_998),
.B2(n_1031),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1055),
.A2(n_948),
.B(n_1030),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_991),
.A2(n_997),
.B(n_1003),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_944),
.B(n_986),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_968),
.B(n_969),
.Y(n_1113)
);

BUFx3_ASAP7_75t_L g1114 ( 
.A(n_993),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1037),
.B(n_1019),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1035),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_976),
.A2(n_982),
.B(n_983),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1003),
.B(n_1058),
.Y(n_1118)
);

NOR2x1_ASAP7_75t_R g1119 ( 
.A(n_1059),
.B(n_942),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1059),
.A2(n_1057),
.B(n_1028),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_1037),
.B(n_975),
.Y(n_1121)
);

AO32x2_ASAP7_75t_L g1122 ( 
.A1(n_933),
.A2(n_1000),
.A3(n_942),
.B1(n_1054),
.B2(n_984),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_930),
.B(n_1041),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_SL g1124 ( 
.A(n_1007),
.B(n_938),
.C(n_990),
.Y(n_1124)
);

AO31x2_ASAP7_75t_L g1125 ( 
.A1(n_933),
.A2(n_1000),
.A3(n_1054),
.B(n_978),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_975),
.A2(n_1061),
.B1(n_1028),
.B2(n_959),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_947),
.A2(n_952),
.B(n_1002),
.Y(n_1127)
);

OR2x2_ASAP7_75t_L g1128 ( 
.A(n_952),
.B(n_1002),
.Y(n_1128)
);

NAND3xp33_ASAP7_75t_L g1129 ( 
.A(n_987),
.B(n_952),
.C(n_1002),
.Y(n_1129)
);

AO21x2_ASAP7_75t_L g1130 ( 
.A1(n_1032),
.A2(n_1045),
.B(n_1052),
.Y(n_1130)
);

AOI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1045),
.A2(n_1052),
.B(n_1053),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1056),
.A2(n_993),
.B(n_1001),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1056),
.B(n_955),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_L g1134 ( 
.A(n_1059),
.B(n_811),
.Y(n_1134)
);

AOI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_971),
.A2(n_882),
.B1(n_783),
.B2(n_405),
.C(n_307),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_L g1136 ( 
.A1(n_957),
.A2(n_601),
.B(n_604),
.C(n_882),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1046),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_935),
.A2(n_836),
.B(n_840),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_957),
.A2(n_932),
.B(n_1033),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_946),
.B(n_310),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_955),
.B(n_1009),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_988),
.A2(n_882),
.B1(n_783),
.B2(n_971),
.Y(n_1142)
);

AOI21x1_ASAP7_75t_L g1143 ( 
.A1(n_966),
.A2(n_916),
.B(n_1027),
.Y(n_1143)
);

AOI221xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1011),
.A2(n_882),
.B1(n_1014),
.B2(n_754),
.C(n_957),
.Y(n_1144)
);

CKINVDCx8_ASAP7_75t_R g1145 ( 
.A(n_931),
.Y(n_1145)
);

AO32x2_ASAP7_75t_L g1146 ( 
.A1(n_1014),
.A2(n_1011),
.A3(n_1043),
.B1(n_1027),
.B2(n_783),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_SL g1147 ( 
.A1(n_1014),
.A2(n_604),
.B(n_1011),
.C(n_999),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_988),
.A2(n_882),
.B1(n_783),
.B2(n_971),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_931),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_957),
.A2(n_932),
.B(n_1033),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1028),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_935),
.A2(n_836),
.B(n_840),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1046),
.Y(n_1153)
);

INVxp67_ASAP7_75t_SL g1154 ( 
.A(n_1050),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_931),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_957),
.A2(n_932),
.B(n_601),
.Y(n_1156)
);

AO32x2_ASAP7_75t_L g1157 ( 
.A1(n_1014),
.A2(n_1011),
.A3(n_1043),
.B1(n_1027),
.B2(n_783),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_955),
.B(n_1009),
.Y(n_1158)
);

INVx6_ASAP7_75t_L g1159 ( 
.A(n_939),
.Y(n_1159)
);

O2A1O1Ixp5_ASAP7_75t_SL g1160 ( 
.A1(n_1014),
.A2(n_604),
.B(n_1011),
.C(n_999),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_SL g1161 ( 
.A1(n_974),
.A2(n_1048),
.B(n_996),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1046),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1040),
.A2(n_799),
.B(n_1042),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_SL g1164 ( 
.A1(n_957),
.A2(n_1063),
.B(n_923),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_957),
.A2(n_1063),
.B(n_923),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_935),
.A2(n_836),
.B(n_840),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1040),
.A2(n_799),
.B(n_1042),
.Y(n_1167)
);

INVx3_ASAP7_75t_SL g1168 ( 
.A(n_939),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_939),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_935),
.A2(n_836),
.B(n_840),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1046),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_988),
.A2(n_882),
.B1(n_783),
.B2(n_971),
.Y(n_1172)
);

OAI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_946),
.A2(n_882),
.B1(n_601),
.B2(n_957),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1040),
.A2(n_799),
.B(n_1042),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_955),
.B(n_1009),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1040),
.A2(n_799),
.B(n_1042),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_955),
.B(n_1009),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_946),
.A2(n_882),
.B(n_601),
.C(n_943),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_931),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_935),
.A2(n_836),
.B(n_840),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1040),
.A2(n_799),
.B(n_1042),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_SL g1182 ( 
.A1(n_957),
.A2(n_1063),
.B(n_923),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_931),
.B(n_459),
.Y(n_1183)
);

BUFx8_ASAP7_75t_L g1184 ( 
.A(n_931),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_957),
.A2(n_932),
.B(n_966),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_939),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1040),
.A2(n_799),
.B(n_1042),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_931),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_957),
.A2(n_932),
.B(n_601),
.Y(n_1189)
);

BUFx2_ASAP7_75t_L g1190 ( 
.A(n_931),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_955),
.B(n_1009),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_1108),
.B(n_1151),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1173),
.A2(n_1136),
.B(n_1178),
.Y(n_1193)
);

AO21x2_ASAP7_75t_L g1194 ( 
.A1(n_1094),
.A2(n_1078),
.B(n_1156),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1142),
.B(n_1148),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1186),
.Y(n_1196)
);

OA21x2_ASAP7_75t_L g1197 ( 
.A1(n_1086),
.A2(n_1094),
.B(n_1139),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1183),
.Y(n_1198)
);

CKINVDCx14_ASAP7_75t_R g1199 ( 
.A(n_1096),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1135),
.A2(n_1148),
.B1(n_1142),
.B2(n_1172),
.Y(n_1200)
);

BUFx4f_ASAP7_75t_L g1201 ( 
.A(n_1105),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1188),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1168),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1138),
.A2(n_1166),
.B(n_1152),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1163),
.A2(n_1187),
.B(n_1176),
.Y(n_1205)
);

AO21x2_ASAP7_75t_L g1206 ( 
.A1(n_1189),
.A2(n_1161),
.B(n_1065),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1172),
.B(n_1140),
.Y(n_1207)
);

OA21x2_ASAP7_75t_L g1208 ( 
.A1(n_1139),
.A2(n_1150),
.B(n_1110),
.Y(n_1208)
);

AO21x2_ASAP7_75t_L g1209 ( 
.A1(n_1065),
.A2(n_1143),
.B(n_1150),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1167),
.A2(n_1174),
.B(n_1181),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1170),
.A2(n_1180),
.A3(n_1069),
.B(n_1085),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1158),
.B(n_1175),
.Y(n_1212)
);

AO21x2_ASAP7_75t_L g1213 ( 
.A1(n_1070),
.A2(n_1081),
.B(n_1088),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1159),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1164),
.A2(n_1165),
.B(n_1182),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1072),
.B(n_1066),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1137),
.B(n_1153),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1117),
.A2(n_1090),
.B(n_1075),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1162),
.B(n_1171),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1084),
.A2(n_1111),
.B(n_1144),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1177),
.B(n_1191),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1093),
.A2(n_1092),
.B1(n_1099),
.B2(n_1100),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1100),
.B(n_1068),
.Y(n_1223)
);

OR2x6_ASAP7_75t_L g1224 ( 
.A(n_1109),
.B(n_1091),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1097),
.A2(n_1144),
.B1(n_1082),
.B2(n_1098),
.C(n_1111),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1154),
.B(n_1097),
.Y(n_1226)
);

NAND2x1p5_ASAP7_75t_L g1227 ( 
.A(n_1151),
.B(n_1115),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1159),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1190),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1123),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1118),
.A2(n_1077),
.B(n_1102),
.C(n_1133),
.Y(n_1231)
);

BUFx2_ASAP7_75t_L g1232 ( 
.A(n_1080),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1068),
.B(n_1149),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1082),
.A2(n_1098),
.B1(n_1185),
.B2(n_1116),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1074),
.A2(n_1121),
.B1(n_1129),
.B2(n_1091),
.Y(n_1235)
);

AOI221x1_ASAP7_75t_L g1236 ( 
.A1(n_1120),
.A2(n_1129),
.B1(n_1126),
.B2(n_1160),
.C(n_1147),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1103),
.A2(n_1134),
.B(n_1067),
.C(n_1113),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1112),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1101),
.A2(n_1131),
.B(n_1127),
.Y(n_1239)
);

CKINVDCx16_ASAP7_75t_R g1240 ( 
.A(n_1106),
.Y(n_1240)
);

BUFx2_ASAP7_75t_SL g1241 ( 
.A(n_1169),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1184),
.Y(n_1242)
);

BUFx3_ASAP7_75t_L g1243 ( 
.A(n_1184),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1128),
.Y(n_1244)
);

BUFx3_ASAP7_75t_L g1245 ( 
.A(n_1169),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1114),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_SL g1247 ( 
.A1(n_1146),
.A2(n_1157),
.B1(n_1132),
.B2(n_1155),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1146),
.A2(n_1157),
.B1(n_1179),
.B2(n_1095),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1089),
.A2(n_1104),
.B1(n_1107),
.B2(n_1157),
.C(n_1146),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1083),
.A2(n_1145),
.B1(n_1124),
.B2(n_1076),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1119),
.A2(n_1130),
.B(n_1073),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1119),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1122),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1087),
.A2(n_1122),
.B(n_1125),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1121),
.B(n_1067),
.Y(n_1255)
);

BUFx10_ASAP7_75t_L g1256 ( 
.A(n_1159),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1188),
.Y(n_1257)
);

AO31x2_ASAP7_75t_L g1258 ( 
.A1(n_1173),
.A2(n_1078),
.A3(n_957),
.B(n_1086),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1159),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1094),
.A2(n_882),
.B(n_1173),
.C(n_943),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1186),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_SL g1262 ( 
.A1(n_1178),
.A2(n_1173),
.B(n_957),
.C(n_882),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1094),
.A2(n_1078),
.B(n_1189),
.Y(n_1263)
);

AND2x6_ASAP7_75t_L g1264 ( 
.A(n_1142),
.B(n_882),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1071),
.Y(n_1265)
);

BUFx8_ASAP7_75t_L g1266 ( 
.A(n_1186),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1148),
.B2(n_988),
.Y(n_1267)
);

BUFx8_ASAP7_75t_L g1268 ( 
.A(n_1186),
.Y(n_1268)
);

AOI221x1_ASAP7_75t_L g1269 ( 
.A1(n_1173),
.A2(n_1178),
.B1(n_1094),
.B2(n_1098),
.C(n_1156),
.Y(n_1269)
);

INVx3_ASAP7_75t_L g1270 ( 
.A(n_1151),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1094),
.A2(n_1152),
.B(n_1138),
.Y(n_1271)
);

NOR2x1_ASAP7_75t_L g1272 ( 
.A(n_1079),
.B(n_1141),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1096),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1173),
.B(n_1142),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1105),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1105),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1173),
.A2(n_882),
.B1(n_988),
.B2(n_1135),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1135),
.B(n_1178),
.C(n_1148),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1178),
.A2(n_1173),
.B(n_882),
.C(n_1094),
.Y(n_1279)
);

CKINVDCx6p67_ASAP7_75t_R g1280 ( 
.A(n_1105),
.Y(n_1280)
);

AO21x2_ASAP7_75t_L g1281 ( 
.A1(n_1094),
.A2(n_1078),
.B(n_1189),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1094),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_1186),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1148),
.B2(n_988),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1173),
.B(n_1142),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1173),
.A2(n_1136),
.B(n_1178),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1173),
.A2(n_1078),
.A3(n_957),
.B(n_1086),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1071),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1188),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1094),
.A2(n_1078),
.B(n_1189),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1198),
.B(n_1246),
.Y(n_1291)
);

OA21x2_ASAP7_75t_L g1292 ( 
.A1(n_1269),
.A2(n_1236),
.B(n_1193),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1244),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1201),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1216),
.B(n_1223),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1223),
.B(n_1217),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1198),
.B(n_1228),
.Y(n_1297)
);

BUFx10_ASAP7_75t_L g1298 ( 
.A(n_1203),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1219),
.B(n_1226),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1226),
.B(n_1230),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1221),
.B(n_1272),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1215),
.A2(n_1260),
.B(n_1237),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1256),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1215),
.A2(n_1271),
.B(n_1279),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_SL g1305 ( 
.A1(n_1279),
.A2(n_1212),
.B(n_1278),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1212),
.B(n_1207),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1278),
.A2(n_1284),
.B(n_1267),
.C(n_1207),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1195),
.B(n_1255),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1238),
.B(n_1222),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1265),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1274),
.A2(n_1285),
.B(n_1282),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1222),
.B(n_1274),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1285),
.B(n_1282),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1200),
.B(n_1264),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1202),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1248),
.B(n_1249),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1200),
.B(n_1264),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1264),
.B(n_1277),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1277),
.A2(n_1284),
.B(n_1267),
.C(n_1193),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1276),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1224),
.A2(n_1248),
.B1(n_1247),
.B2(n_1235),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1288),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1271),
.A2(n_1262),
.B(n_1204),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1286),
.A2(n_1231),
.B(n_1250),
.C(n_1235),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1286),
.A2(n_1250),
.B(n_1224),
.C(n_1225),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1201),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1273),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1264),
.B(n_1233),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1224),
.A2(n_1225),
.B(n_1197),
.C(n_1233),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1264),
.B(n_1229),
.Y(n_1330)
);

OR2x2_ASAP7_75t_L g1331 ( 
.A(n_1257),
.B(n_1289),
.Y(n_1331)
);

O2A1O1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1197),
.A2(n_1290),
.B(n_1263),
.C(n_1194),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1256),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1232),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1247),
.B(n_1227),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1208),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1208),
.B(n_1194),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1270),
.B(n_1234),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1234),
.B(n_1192),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1192),
.B(n_1199),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1281),
.A2(n_1211),
.B(n_1287),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1245),
.Y(n_1342)
);

OAI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1252),
.A2(n_1241),
.B1(n_1275),
.B2(n_1280),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1252),
.A2(n_1206),
.B(n_1209),
.C(n_1251),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1242),
.A2(n_1243),
.B1(n_1240),
.B2(n_1261),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1258),
.B(n_1220),
.Y(n_1346)
);

OA21x2_ASAP7_75t_L g1347 ( 
.A1(n_1218),
.A2(n_1254),
.B(n_1205),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1253),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1214),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_1266),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1259),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1196),
.B(n_1261),
.Y(n_1352)
);

AND2x2_ASAP7_75t_SL g1353 ( 
.A(n_1196),
.B(n_1261),
.Y(n_1353)
);

INVx3_ASAP7_75t_SL g1354 ( 
.A(n_1283),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1213),
.A2(n_1239),
.B(n_1210),
.C(n_1266),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1196),
.B(n_1268),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1268),
.Y(n_1357)
);

CKINVDCx14_ASAP7_75t_R g1358 ( 
.A(n_1199),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1219),
.B(n_1244),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1216),
.B(n_1244),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1216),
.B(n_1244),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1269),
.A2(n_1236),
.B(n_1193),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1215),
.A2(n_1094),
.B(n_1138),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1221),
.B(n_1272),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1200),
.A2(n_1148),
.B1(n_1172),
.B2(n_1142),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1216),
.B(n_1244),
.Y(n_1366)
);

BUFx12f_ASAP7_75t_L g1367 ( 
.A(n_1276),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1269),
.A2(n_1236),
.B(n_1193),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1336),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1346),
.B(n_1337),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1348),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1304),
.B(n_1323),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1347),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1313),
.B(n_1306),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1347),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1299),
.B(n_1300),
.Y(n_1376)
);

INVx5_ASAP7_75t_L g1377 ( 
.A(n_1302),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1332),
.B(n_1335),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1316),
.B(n_1292),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1363),
.B(n_1322),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1310),
.Y(n_1381)
);

AO21x2_ASAP7_75t_L g1382 ( 
.A1(n_1319),
.A2(n_1344),
.B(n_1311),
.Y(n_1382)
);

INVx11_ASAP7_75t_L g1383 ( 
.A(n_1367),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1368),
.B(n_1362),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1344),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1312),
.B(n_1307),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1339),
.Y(n_1387)
);

INVx4_ASAP7_75t_L g1388 ( 
.A(n_1362),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1355),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1338),
.B(n_1296),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1330),
.B(n_1321),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1295),
.B(n_1328),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1318),
.B(n_1305),
.Y(n_1393)
);

INVxp67_ASAP7_75t_SL g1394 ( 
.A(n_1324),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1355),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1315),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1293),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1301),
.B(n_1364),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1366),
.B(n_1361),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1329),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1340),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1309),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1329),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1359),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1342),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1314),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1369),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1402),
.B(n_1307),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1370),
.B(n_1360),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1370),
.B(n_1380),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1377),
.A2(n_1324),
.B(n_1325),
.C(n_1394),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1370),
.B(n_1380),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1386),
.B(n_1365),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1377),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1380),
.B(n_1308),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1369),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1381),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1371),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1380),
.B(n_1325),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1373),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1378),
.B(n_1334),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1405),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1381),
.Y(n_1424)
);

OAI33xp33_ASAP7_75t_L g1425 ( 
.A1(n_1385),
.A2(n_1317),
.A3(n_1343),
.B1(n_1345),
.B2(n_1331),
.B3(n_1357),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_1385),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1378),
.B(n_1341),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1377),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1378),
.B(n_1372),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1397),
.Y(n_1430)
);

AOI221xp5_ASAP7_75t_L g1431 ( 
.A1(n_1413),
.A2(n_1386),
.B1(n_1394),
.B2(n_1400),
.C(n_1403),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1407),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1413),
.A2(n_1377),
.B1(n_1382),
.B2(n_1403),
.Y(n_1433)
);

NAND3xp33_ASAP7_75t_L g1434 ( 
.A(n_1411),
.B(n_1393),
.C(n_1403),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_R g1435 ( 
.A(n_1408),
.B(n_1320),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1411),
.B(n_1393),
.C(n_1400),
.Y(n_1436)
);

OAI322xp33_ASAP7_75t_L g1437 ( 
.A1(n_1408),
.A2(n_1398),
.A3(n_1400),
.B1(n_1374),
.B2(n_1391),
.C1(n_1376),
.C2(n_1402),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1428),
.A2(n_1377),
.B1(n_1391),
.B2(n_1374),
.Y(n_1438)
);

OAI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1421),
.A2(n_1377),
.B1(n_1391),
.B2(n_1393),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1425),
.B(n_1358),
.Y(n_1440)
);

NOR2x1_ASAP7_75t_L g1441 ( 
.A(n_1428),
.B(n_1382),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1409),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1414),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1418),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1412),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1407),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1415),
.B(n_1377),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1425),
.A2(n_1377),
.B1(n_1382),
.B2(n_1406),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1417),
.B(n_1388),
.Y(n_1450)
);

OAI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1426),
.A2(n_1376),
.B1(n_1406),
.B2(n_1402),
.C(n_1297),
.Y(n_1451)
);

NAND4xp25_ASAP7_75t_SL g1452 ( 
.A(n_1427),
.B(n_1379),
.C(n_1356),
.D(n_1352),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1421),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1454)
);

OAI211xp5_ASAP7_75t_L g1455 ( 
.A1(n_1427),
.A2(n_1379),
.B(n_1388),
.C(n_1384),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1422),
.Y(n_1456)
);

OAI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1426),
.A2(n_1406),
.B1(n_1402),
.B2(n_1351),
.C(n_1401),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1415),
.B(n_1404),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1419),
.A2(n_1382),
.B1(n_1406),
.B2(n_1379),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1416),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1431),
.B(n_1409),
.Y(n_1461)
);

INVx5_ASAP7_75t_L g1462 ( 
.A(n_1444),
.Y(n_1462)
);

AND2x4_ASAP7_75t_SL g1463 ( 
.A(n_1442),
.B(n_1415),
.Y(n_1463)
);

INVx4_ASAP7_75t_SL g1464 ( 
.A(n_1444),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1432),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1432),
.Y(n_1466)
);

CKINVDCx16_ASAP7_75t_R g1467 ( 
.A(n_1435),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1447),
.Y(n_1468)
);

NAND3xp33_ASAP7_75t_L g1469 ( 
.A(n_1434),
.B(n_1389),
.C(n_1395),
.Y(n_1469)
);

BUFx3_ASAP7_75t_L g1470 ( 
.A(n_1444),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1446),
.B(n_1429),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1449),
.B(n_1392),
.Y(n_1472)
);

INVx5_ASAP7_75t_L g1473 ( 
.A(n_1444),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1436),
.B(n_1389),
.C(n_1395),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1460),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1456),
.A2(n_1420),
.B(n_1423),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1445),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1433),
.A2(n_1419),
.B(n_1427),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1453),
.B(n_1412),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1450),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1444),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1440),
.A2(n_1429),
.B(n_1419),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1450),
.Y(n_1483)
);

INVx4_ASAP7_75t_L g1484 ( 
.A(n_1456),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1458),
.B(n_1424),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1461),
.B(n_1412),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1464),
.B(n_1471),
.Y(n_1487)
);

INVx1_ASAP7_75t_SL g1488 ( 
.A(n_1467),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1482),
.B(n_1459),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1477),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1464),
.B(n_1471),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1464),
.B(n_1446),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1476),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1472),
.B(n_1390),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1473),
.B(n_1443),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1469),
.A2(n_1382),
.B1(n_1452),
.B2(n_1372),
.Y(n_1499)
);

OAI321xp33_ASAP7_75t_L g1500 ( 
.A1(n_1474),
.A2(n_1438),
.A3(n_1451),
.B1(n_1439),
.B2(n_1457),
.C(n_1455),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1477),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1473),
.B(n_1454),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1462),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1465),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1465),
.Y(n_1505)
);

NAND4xp25_ASAP7_75t_L g1506 ( 
.A(n_1478),
.B(n_1441),
.C(n_1291),
.D(n_1396),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1466),
.Y(n_1507)
);

NOR2x1_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_1437),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1454),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1462),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1462),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1485),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1462),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1485),
.B(n_1399),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1488),
.B(n_1508),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1493),
.B(n_1481),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1490),
.Y(n_1519)
);

AOI211x1_ASAP7_75t_L g1520 ( 
.A1(n_1506),
.A2(n_1479),
.B(n_1468),
.C(n_1475),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1510),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1501),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1508),
.B(n_1467),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1501),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1510),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1493),
.B(n_1481),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1487),
.B(n_1481),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1528)
);

INVx2_ASAP7_75t_SL g1529 ( 
.A(n_1487),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1492),
.B(n_1496),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1511),
.B(n_1473),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1504),
.Y(n_1532)
);

NAND2x1_ASAP7_75t_L g1533 ( 
.A(n_1503),
.B(n_1484),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1514),
.B(n_1462),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1504),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1491),
.B(n_1462),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1505),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1507),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1491),
.Y(n_1541)
);

NOR2x1_ASAP7_75t_L g1542 ( 
.A(n_1511),
.B(n_1484),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1507),
.Y(n_1543)
);

INVxp67_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1494),
.Y(n_1545)
);

INVxp67_ASAP7_75t_L g1546 ( 
.A(n_1498),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1494),
.B(n_1502),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1500),
.B(n_1484),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1486),
.B(n_1442),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1511),
.B(n_1463),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1543),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1543),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1516),
.B(n_1489),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1532),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1523),
.B(n_1497),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1535),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1541),
.B(n_1383),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1536),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1547),
.B(n_1515),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1521),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1536),
.B(n_1502),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1521),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1533),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1544),
.B(n_1509),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1546),
.B(n_1509),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1545),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1537),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1527),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1527),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_SL g1571 ( 
.A(n_1531),
.B(n_1511),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1539),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1540),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1517),
.B(n_1503),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1525),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1562),
.B(n_1529),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1561),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1559),
.Y(n_1578)
);

OAI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1553),
.A2(n_1548),
.B1(n_1529),
.B2(n_1499),
.C(n_1528),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1561),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1561),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1559),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1567),
.B(n_1569),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1570),
.B(n_1548),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1563),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1525),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1563),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1556),
.A2(n_1542),
.B(n_1526),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1556),
.B(n_1517),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1560),
.B(n_1520),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1560),
.B(n_1526),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1555),
.A2(n_1531),
.B1(n_1534),
.B2(n_1533),
.C(n_1530),
.Y(n_1592)
);

NAND3xp33_ASAP7_75t_L g1593 ( 
.A(n_1571),
.B(n_1538),
.C(n_1519),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1565),
.B(n_1549),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1578),
.B(n_1563),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1579),
.A2(n_1566),
.B1(n_1571),
.B2(n_1558),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1589),
.B(n_1574),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1577),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1580),
.Y(n_1599)
);

NOR2xp33_ASAP7_75t_L g1600 ( 
.A(n_1582),
.B(n_1383),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1576),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1582),
.B(n_1575),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1576),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1581),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1585),
.Y(n_1605)
);

NOR4xp25_ASAP7_75t_L g1606 ( 
.A(n_1602),
.B(n_1583),
.C(n_1584),
.D(n_1593),
.Y(n_1606)
);

NAND4xp75_ASAP7_75t_L g1607 ( 
.A(n_1595),
.B(n_1588),
.C(n_1587),
.D(n_1586),
.Y(n_1607)
);

AOI221xp5_ASAP7_75t_L g1608 ( 
.A1(n_1596),
.A2(n_1590),
.B1(n_1592),
.B2(n_1594),
.C(n_1591),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1596),
.A2(n_1575),
.B(n_1589),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1600),
.A2(n_1550),
.B1(n_1574),
.B2(n_1564),
.Y(n_1610)
);

NAND4xp25_ASAP7_75t_L g1611 ( 
.A(n_1600),
.B(n_1575),
.C(n_1573),
.D(n_1572),
.Y(n_1611)
);

AO21x1_ASAP7_75t_L g1612 ( 
.A1(n_1603),
.A2(n_1531),
.B(n_1551),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1601),
.A2(n_1564),
.B(n_1538),
.Y(n_1613)
);

NOR3x1_ASAP7_75t_L g1614 ( 
.A(n_1598),
.B(n_1557),
.C(n_1554),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_SL g1615 ( 
.A1(n_1609),
.A2(n_1603),
.B1(n_1604),
.B2(n_1599),
.C(n_1597),
.Y(n_1615)
);

AOI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1606),
.A2(n_1605),
.B1(n_1573),
.B2(n_1572),
.C(n_1568),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1607),
.A2(n_1564),
.B(n_1550),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1614),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_L g1619 ( 
.A1(n_1608),
.A2(n_1564),
.B(n_1550),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1619),
.A2(n_1610),
.B1(n_1611),
.B2(n_1613),
.C(n_1554),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1617),
.Y(n_1621)
);

NAND3xp33_ASAP7_75t_L g1622 ( 
.A(n_1616),
.B(n_1568),
.C(n_1557),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1618),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1615),
.B(n_1612),
.Y(n_1624)
);

NOR3xp33_ASAP7_75t_L g1625 ( 
.A(n_1619),
.B(n_1294),
.C(n_1350),
.Y(n_1625)
);

INVx1_ASAP7_75t_SL g1626 ( 
.A(n_1623),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1625),
.A2(n_1551),
.B1(n_1552),
.B2(n_1513),
.Y(n_1627)
);

XNOR2xp5_ASAP7_75t_L g1628 ( 
.A(n_1620),
.B(n_1353),
.Y(n_1628)
);

OAI321xp33_ASAP7_75t_L g1629 ( 
.A1(n_1624),
.A2(n_1552),
.A3(n_1530),
.B1(n_1524),
.B2(n_1522),
.C(n_1518),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1622),
.Y(n_1630)
);

INVxp33_ASAP7_75t_SL g1631 ( 
.A(n_1626),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1628),
.Y(n_1632)
);

BUFx12f_ASAP7_75t_L g1633 ( 
.A(n_1630),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1631),
.B(n_1621),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1634),
.A2(n_1632),
.B(n_1627),
.C(n_1631),
.Y(n_1635)
);

INVxp67_ASAP7_75t_L g1636 ( 
.A(n_1635),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1635),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1637),
.Y(n_1638)
);

AOI21xp33_ASAP7_75t_L g1639 ( 
.A1(n_1636),
.A2(n_1633),
.B(n_1629),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1638),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1639),
.B(n_1513),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1640),
.A2(n_1327),
.B(n_1303),
.Y(n_1642)
);

AOI21xp5_ASAP7_75t_L g1643 ( 
.A1(n_1642),
.A2(n_1641),
.B(n_1383),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1643),
.B(n_1354),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1644),
.A2(n_1326),
.B(n_1513),
.Y(n_1645)
);

AOI22xp5_ASAP7_75t_L g1646 ( 
.A1(n_1645),
.A2(n_1298),
.B1(n_1333),
.B2(n_1349),
.Y(n_1646)
);

AOI211xp5_ASAP7_75t_L g1647 ( 
.A1(n_1646),
.A2(n_1333),
.B(n_1298),
.C(n_1495),
.Y(n_1647)
);


endmodule