module fake_jpeg_14484_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_8),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_53),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_54),
.B1(n_47),
.B2(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_14),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_43),
.B1(n_35),
.B2(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_4),
.Y(n_62)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_47),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_48),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_40),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_4),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_56),
.B1(n_57),
.B2(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_40),
.B1(n_6),
.B2(n_7),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_80),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g81 ( 
.A1(n_62),
.A2(n_40),
.A3(n_19),
.B1(n_22),
.B2(n_33),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_18),
.C(n_30),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_94),
.B1(n_5),
.B2(n_8),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_93),
.B1(n_12),
.B2(n_23),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_78),
.C(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_9),
.C(n_10),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_68),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_96),
.C(n_93),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_89),
.B1(n_86),
.B2(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_100),
.C(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_105),
.B(n_96),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_84),
.C(n_97),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_101),
.A3(n_87),
.B1(n_91),
.B2(n_29),
.C1(n_25),
.C2(n_27),
.Y(n_110)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_110),
.Y(n_111)
);


endmodule