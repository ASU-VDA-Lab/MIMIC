module fake_netlist_6_3570_n_4426 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_442, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_443, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_433, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4426);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_433;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4426;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3813;
wire n_3660;
wire n_801;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_700;
wire n_3773;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2534;
wire n_2353;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_4285;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_461;
wire n_1371;
wire n_1285;
wire n_873;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_522;
wire n_2919;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_2356;
wire n_1143;
wire n_1511;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_616;
wire n_658;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_2739;
wire n_1300;
wire n_641;
wire n_2480;
wire n_1541;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4071;
wire n_4255;
wire n_4403;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_551;
wire n_699;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_451;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_2190;
wire n_1918;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4366;
wire n_3446;
wire n_4158;
wire n_4377;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_966;
wire n_3888;
wire n_2908;
wire n_3168;
wire n_764;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3092;
wire n_3055;
wire n_3492;
wire n_3895;
wire n_4369;
wire n_3966;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_882;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1950;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2749;
wire n_2008;
wire n_3298;
wire n_2192;
wire n_3281;
wire n_2254;
wire n_2345;
wire n_3346;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4386;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_4072;
wire n_3940;
wire n_4220;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_3917;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2519;
wire n_2319;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_696;
wire n_1515;
wire n_961;
wire n_4356;
wire n_3510;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2972;
wire n_2194;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3696;
wire n_3780;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3450;
wire n_3337;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_2750;
wire n_2558;
wire n_2893;
wire n_2775;
wire n_1208;
wire n_1523;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_2767;
wire n_794;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_1139;
wire n_1714;
wire n_872;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_2747;
wire n_1513;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2643;
wire n_2590;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_765;
wire n_1492;
wire n_987;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_4058;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3229;
wire n_3348;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_2335;
wire n_1529;
wire n_2473;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2667;
wire n_2539;
wire n_2698;
wire n_4096;
wire n_1431;
wire n_4123;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2958;
wire n_1577;
wire n_2948;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_2857;
wire n_446;
wire n_3693;
wire n_3788;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3203;
wire n_3325;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_1284;
wire n_745;
wire n_2424;
wire n_2296;
wire n_1604;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1398;
wire n_1201;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_2442;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3540;
wire n_3577;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3226;
wire n_3364;
wire n_4176;
wire n_4020;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_4261;
wire n_4204;
wire n_3894;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_4237;
wire n_3986;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1892;
wire n_1459;
wire n_1614;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4034;
wire n_1617;
wire n_4056;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3284;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_3205;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4132;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_3360;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2993;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4126;
wire n_1129;
wire n_3870;
wire n_4003;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_2181;
wire n_1594;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4067;
wire n_4252;
wire n_4357;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3250;
wire n_1934;
wire n_3276;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_4420;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4234;
wire n_4304;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1397;
wire n_1037;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4189;
wire n_4270;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_1320;
wire n_2716;
wire n_3249;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3238;
wire n_2235;
wire n_3529;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4109;
wire n_4192;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_4038;
wire n_4131;
wire n_2790;
wire n_3957;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2373;
wire n_2050;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4174;
wire n_1870;
wire n_2964;
wire n_4144;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3475;
wire n_662;
wire n_3501;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_450;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2970;
wire n_2084;
wire n_2167;
wire n_3676;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_4122;
wire n_3988;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_482;
wire n_934;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_3588;
wire n_4209;
wire n_2871;
wire n_4135;
wire n_4279;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4183;
wire n_1489;
wire n_4321;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_3292;
wire n_1271;
wire n_1496;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_2258;
wire n_1485;
wire n_1640;
wire n_4040;
wire n_804;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_799;
wire n_1548;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_3007;
wire n_2809;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4084;
wire n_3558;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_2695;
wire n_4269;
wire n_3818;
wire n_4035;
wire n_743;
wire n_766;
wire n_3124;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2888;
wire n_2715;
wire n_2793;
wire n_1804;
wire n_2923;
wire n_3711;
wire n_3776;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_3308;
wire n_1113;
wire n_2833;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_1742;
wire n_3190;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4173;
wire n_3135;
wire n_4324;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2186;
wire n_2163;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_2020;
wire n_1643;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3701;
wire n_3154;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_452;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_1303;
wire n_761;
wire n_2769;
wire n_4342;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3551;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4027;
wire n_4373;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_445;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_3584;
wire n_3486;
wire n_4086;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2743;
wire n_2437;
wire n_3962;
wire n_708;
wire n_1973;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_1058;
wire n_854;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3802;
wire n_3868;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2111;
wire n_2466;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3697;
wire n_3643;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3408;
wire n_3461;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4089;
wire n_4351;
wire n_4346;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2723;
wire n_2440;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2478;
wire n_1619;
wire n_2303;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_635;
wire n_1194;
wire n_3374;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4051;
wire n_1051;
wire n_3976;
wire n_4254;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_3147;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_633;
wire n_1170;
wire n_665;
wire n_2221;
wire n_1629;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_2280;
wire n_1557;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_3274;
wire n_2899;
wire n_3333;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3431;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_4030;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_236),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_416),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_419),
.Y(n_447)
);

BUFx10_ASAP7_75t_L g448 ( 
.A(n_206),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_277),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_385),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_22),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_62),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_209),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_16),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_263),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_175),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_181),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_39),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_330),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_259),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_369),
.Y(n_461)
);

BUFx10_ASAP7_75t_L g462 ( 
.A(n_54),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_353),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_165),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_0),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_273),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_429),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_30),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_388),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_32),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_113),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_185),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_179),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_213),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_351),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_62),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_383),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_182),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_282),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_307),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_343),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_279),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_404),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_224),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_389),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_284),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_298),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_193),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_148),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_390),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_164),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_223),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_222),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_162),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_262),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_166),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_196),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_26),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_209),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_188),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_51),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_66),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_60),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_280),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_215),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_367),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_176),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_320),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_341),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_93),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_73),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_349),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_265),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_65),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_162),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_239),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_283),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_313),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_45),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_289),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_211),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_370),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_132),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_315),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_382),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_79),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_299),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_246),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_149),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_266),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_204),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_437),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_288),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_154),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_193),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_106),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_318),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_308),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_346),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_107),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_113),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_196),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_254),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_166),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_188),
.Y(n_548)
);

BUFx10_ASAP7_75t_L g549 ( 
.A(n_98),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_415),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_364),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_438),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_221),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_26),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_38),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_23),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_41),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_156),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_31),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_386),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_122),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_88),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_80),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_355),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_240),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_189),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_83),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_149),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_176),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_38),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_197),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_407),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_255),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_339),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_71),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_164),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_36),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_14),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_302),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_47),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_167),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_106),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_444),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_423),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_252),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_36),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_181),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_115),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_130),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_89),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_231),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_163),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_19),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_293),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_269),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_186),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_393),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_158),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_439),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_225),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_53),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_167),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_440),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_37),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_129),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_297),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_32),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_326),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_42),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_254),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_373),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_67),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_384),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_409),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_435),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_186),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_120),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_216),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_235),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_265),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_387),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_25),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_264),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_422),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_15),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_257),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_377),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_79),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_352),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_112),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_197),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_309),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_374),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_286),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_258),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_10),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_262),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_328),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_216),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_200),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_96),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_101),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_182),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_202),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_426),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_179),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_155),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_147),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_88),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_144),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_114),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_224),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_310),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_9),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_28),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_274),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_165),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_4),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_300),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_175),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_291),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_324),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_331),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_17),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_41),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_138),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_379),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_413),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_354),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_141),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_93),
.Y(n_671)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_332),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_425),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_338),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_406),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_259),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_344),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_51),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_306),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_241),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_27),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_159),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_177),
.Y(n_683)
);

INVx1_ASAP7_75t_SL g684 ( 
.A(n_137),
.Y(n_684)
);

CKINVDCx14_ASAP7_75t_R g685 ( 
.A(n_134),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_428),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_358),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_239),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_252),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_222),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_145),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_210),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_73),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_218),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_194),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_1),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_238),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_63),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_45),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_305),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_230),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_12),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_67),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_46),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_92),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_403),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_363),
.Y(n_707)
);

INVx1_ASAP7_75t_SL g708 ( 
.A(n_19),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_40),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_334),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_13),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_48),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_23),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_8),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_250),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_395),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_366),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_215),
.Y(n_718)
);

CKINVDCx14_ASAP7_75t_R g719 ( 
.A(n_399),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_269),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_357),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_58),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_229),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_378),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_397),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_136),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_290),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_226),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_158),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_194),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_200),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_97),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_97),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_268),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_312),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_52),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_234),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_253),
.Y(n_738)
);

BUFx8_ASAP7_75t_SL g739 ( 
.A(n_146),
.Y(n_739)
);

CKINVDCx6p67_ASAP7_75t_R g740 ( 
.A(n_301),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_417),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_210),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_44),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_174),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_1),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_25),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_145),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_136),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_111),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_303),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_340),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_7),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_75),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_319),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_168),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_237),
.Y(n_756)
);

CKINVDCx20_ASAP7_75t_R g757 ( 
.A(n_322),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_221),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_102),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_362),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_63),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_110),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_411),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_20),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_138),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_155),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_223),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_104),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_65),
.Y(n_769)
);

CKINVDCx20_ASAP7_75t_R g770 ( 
.A(n_163),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_506),
.B(n_0),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_459),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_739),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_446),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_526),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_517),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_517),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_517),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_517),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_484),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_517),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_447),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_449),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_517),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_526),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_548),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_604),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_548),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_604),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_450),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_548),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_548),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_548),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_548),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_660),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_660),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_461),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_744),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_463),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_632),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_660),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_660),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_466),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_660),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_467),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_660),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_709),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_477),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_645),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_709),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_709),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_709),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_709),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_709),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_452),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_481),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_452),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_452),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_482),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_546),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_546),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_546),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_744),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_486),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_559),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_559),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_559),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_602),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_487),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_489),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_602),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_602),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_748),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_616),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_493),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_616),
.Y(n_836)
);

INVxp67_ASAP7_75t_L g837 ( 
.A(n_748),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_616),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_651),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_651),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_651),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_697),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_685),
.B(n_2),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_697),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_697),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_512),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_701),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_520),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_669),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_701),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_506),
.B(n_2),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_733),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_733),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_733),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_743),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_515),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_743),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_679),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_521),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_525),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_527),
.Y(n_862)
);

INVx1_ASAP7_75t_SL g863 ( 
.A(n_445),
.Y(n_863)
);

BUFx8_ASAP7_75t_SL g864 ( 
.A(n_505),
.Y(n_864)
);

INVxp33_ASAP7_75t_L g865 ( 
.A(n_453),
.Y(n_865)
);

BUFx2_ASAP7_75t_L g866 ( 
.A(n_495),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_743),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_495),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_528),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_753),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_520),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_753),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_753),
.Y(n_873)
);

CKINVDCx16_ASAP7_75t_R g874 ( 
.A(n_473),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_475),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_579),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_475),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_495),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_530),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_535),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_501),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_501),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_536),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_501),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_576),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_540),
.Y(n_886)
);

BUFx8_ASAP7_75t_SL g887 ( 
.A(n_534),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_576),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_459),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_541),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_488),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_488),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_488),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_542),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_576),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_560),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_590),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_590),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_590),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_550),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_644),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_551),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_757),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_644),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_564),
.Y(n_905)
);

BUFx3_ASAP7_75t_L g906 ( 
.A(n_475),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_644),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_695),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_695),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_574),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_474),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_583),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_597),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_479),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_606),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_560),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_608),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_621),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_627),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_479),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_629),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_672),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_480),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_634),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_560),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_480),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_483),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_453),
.B(n_3),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_633),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_483),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_507),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_695),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_507),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_509),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_638),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_539),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_633),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_455),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_653),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_455),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_468),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_468),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_485),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_485),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_491),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_511),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_672),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_509),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_511),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_663),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_667),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_633),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_523),
.Y(n_953)
);

INVxp67_ASAP7_75t_SL g954 ( 
.A(n_579),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_656),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_674),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_523),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_613),
.B(n_3),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_491),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_675),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_686),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_543),
.Y(n_962)
);

XNOR2x2_ASAP7_75t_R g963 ( 
.A(n_473),
.B(n_4),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_494),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_687),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_710),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_494),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_498),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_719),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_716),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_717),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_498),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_508),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_724),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_504),
.Y(n_975)
);

CKINVDCx20_ASAP7_75t_R g976 ( 
.A(n_725),
.Y(n_976)
);

CKINVDCx20_ASAP7_75t_R g977 ( 
.A(n_735),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_504),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_513),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_513),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_516),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_516),
.Y(n_982)
);

CKINVDCx14_ASAP7_75t_R g983 ( 
.A(n_613),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_529),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_529),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_741),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_532),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_532),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_754),
.Y(n_989)
);

CKINVDCx16_ASAP7_75t_R g990 ( 
.A(n_508),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_763),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_567),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_451),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_454),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_456),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_L g996 ( 
.A(n_510),
.B(n_5),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_520),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_457),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_533),
.Y(n_999)
);

BUFx10_ASAP7_75t_L g1000 ( 
.A(n_474),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_533),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_544),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_567),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_509),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_552),
.Y(n_1005)
);

CKINVDCx16_ASAP7_75t_R g1006 ( 
.A(n_448),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_544),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_575),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_565),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_458),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_575),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_580),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_580),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_460),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_464),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_465),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_581),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_470),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_520),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_471),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_472),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_581),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_476),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_656),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_582),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_478),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_448),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_582),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_552),
.Y(n_1029)
);

CKINVDCx16_ASAP7_75t_R g1030 ( 
.A(n_448),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_492),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_496),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_497),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_499),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_585),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_740),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_585),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_500),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_589),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_520),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_502),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_589),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_503),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_514),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_572),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_448),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_520),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_572),
.Y(n_1048)
);

CKINVDCx16_ASAP7_75t_R g1049 ( 
.A(n_462),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_518),
.Y(n_1050)
);

BUFx8_ASAP7_75t_SL g1051 ( 
.A(n_568),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_591),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_584),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_519),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_524),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_552),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_537),
.Y(n_1057)
);

BUFx2_ASAP7_75t_SL g1058 ( 
.A(n_522),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_584),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_673),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_656),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_599),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_538),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_545),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_599),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_547),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_673),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_553),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_603),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_740),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_591),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_595),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_595),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_673),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_598),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_659),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_598),
.Y(n_1077)
);

CKINVDCx20_ASAP7_75t_R g1078 ( 
.A(n_740),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_600),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_636),
.Y(n_1080)
);

BUFx10_ASAP7_75t_L g1081 ( 
.A(n_522),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_554),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_555),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_659),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_700),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_510),
.B(n_5),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_600),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_659),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_601),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_601),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_556),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_617),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_617),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_557),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_558),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_700),
.B(n_662),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_618),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_618),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_561),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_623),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_562),
.Y(n_1101)
);

CKINVDCx14_ASAP7_75t_R g1102 ( 
.A(n_462),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_623),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_628),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_662),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_628),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_563),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_630),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_630),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_637),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_637),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_566),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_662),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_569),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_700),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_570),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_650),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_650),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_721),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_462),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_654),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_654),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_571),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_682),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_682),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_573),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_721),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_694),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_603),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_577),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_615),
.B(n_6),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_971),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_993),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_780),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1056),
.Y(n_1135)
);

INVx4_ASAP7_75t_R g1136 ( 
.A(n_863),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1056),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1056),
.Y(n_1138)
);

INVxp33_ASAP7_75t_SL g1139 ( 
.A(n_958),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1056),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_1056),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_976),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_1060),
.Y(n_1143)
);

HB1xp67_ASAP7_75t_L g1144 ( 
.A(n_994),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_800),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_977),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1060),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1060),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_995),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_989),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1060),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_998),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_969),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_848),
.Y(n_1154)
);

INVxp67_ASAP7_75t_SL g1155 ( 
.A(n_1060),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_1010),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_774),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_878),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_809),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_878),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_849),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1014),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_881),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_859),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_881),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_782),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_882),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_882),
.Y(n_1168)
);

CKINVDCx20_ASAP7_75t_R g1169 ( 
.A(n_903),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_983),
.B(n_615),
.Y(n_1170)
);

CKINVDCx20_ASAP7_75t_R g1171 ( 
.A(n_1080),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_864),
.Y(n_1172)
);

INVxp67_ASAP7_75t_SL g1173 ( 
.A(n_948),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_887),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_783),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_790),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_884),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_884),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_885),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_885),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_797),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_888),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_888),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_895),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_895),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_779),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_779),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_799),
.Y(n_1188)
);

HB1xp67_ASAP7_75t_L g1189 ( 
.A(n_1015),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_897),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_897),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_1051),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_898),
.Y(n_1193)
);

INVxp67_ASAP7_75t_SL g1194 ( 
.A(n_948),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_803),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_805),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_898),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_922),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_899),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_876),
.B(n_469),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_776),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_776),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_777),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_808),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_947),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1036),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_816),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_819),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1070),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_954),
.B(n_469),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_1078),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_777),
.Y(n_1212)
);

CKINVDCx16_ASAP7_75t_R g1213 ( 
.A(n_874),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_778),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1043),
.Y(n_1215)
);

CKINVDCx20_ASAP7_75t_R g1216 ( 
.A(n_990),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_778),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1003),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_899),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_824),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_901),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_829),
.B(n_614),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_830),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_901),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_904),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1018),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_835),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_904),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_907),
.Y(n_1229)
);

CKINVDCx16_ASAP7_75t_R g1230 ( 
.A(n_1102),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1020),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_907),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_908),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1016),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_846),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_857),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1021),
.Y(n_1237)
);

INVxp67_ASAP7_75t_SL g1238 ( 
.A(n_948),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_908),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_909),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1023),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_860),
.Y(n_1242)
);

INVxp33_ASAP7_75t_L g1243 ( 
.A(n_775),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_909),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_781),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1026),
.B(n_1031),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_781),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_784),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_784),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_861),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_786),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_786),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_788),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_862),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_869),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1016),
.Y(n_1256)
);

INVxp67_ASAP7_75t_SL g1257 ( 
.A(n_875),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_788),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_791),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_791),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_792),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_792),
.Y(n_1262)
);

CKINVDCx20_ASAP7_75t_R g1263 ( 
.A(n_879),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_875),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_793),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_880),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_793),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_883),
.Y(n_1268)
);

NOR2xp67_ASAP7_75t_L g1269 ( 
.A(n_886),
.B(n_890),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_877),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_894),
.Y(n_1271)
);

INVxp33_ASAP7_75t_SL g1272 ( 
.A(n_900),
.Y(n_1272)
);

INVxp67_ASAP7_75t_L g1273 ( 
.A(n_1044),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_877),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_902),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_795),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_905),
.Y(n_1277)
);

INVxp67_ASAP7_75t_SL g1278 ( 
.A(n_906),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_795),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_796),
.Y(n_1280)
);

INVx3_ASAP7_75t_L g1281 ( 
.A(n_848),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_910),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_796),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_912),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_801),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_801),
.Y(n_1286)
);

INVxp67_ASAP7_75t_SL g1287 ( 
.A(n_906),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_802),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_913),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_802),
.Y(n_1290)
);

CKINVDCx16_ASAP7_75t_R g1291 ( 
.A(n_1006),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_R g1292 ( 
.A(n_1032),
.B(n_578),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_804),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_915),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_934),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1033),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_917),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_918),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_804),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_806),
.Y(n_1300)
);

INVxp67_ASAP7_75t_L g1301 ( 
.A(n_1044),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_806),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1034),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_807),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_807),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_810),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_919),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_810),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_921),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1038),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_811),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_924),
.B(n_721),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_811),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1041),
.B(n_594),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_935),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_812),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_812),
.Y(n_1317)
);

BUFx10_ASAP7_75t_L g1318 ( 
.A(n_773),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_813),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_939),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_950),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_951),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1050),
.B(n_594),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_956),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_813),
.Y(n_1325)
);

CKINVDCx20_ASAP7_75t_R g1326 ( 
.A(n_960),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_814),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_814),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_961),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_965),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_772),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_889),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_934),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_966),
.Y(n_1334)
);

INVxp33_ASAP7_75t_SL g1335 ( 
.A(n_970),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_974),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_914),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_986),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_991),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_1054),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_920),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1055),
.B(n_611),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_923),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_868),
.B(n_1004),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1083),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1057),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1063),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1064),
.B(n_1066),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_926),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_927),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_930),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_936),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1068),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1082),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1091),
.B(n_611),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_962),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_931),
.Y(n_1357)
);

INVxp67_ASAP7_75t_SL g1358 ( 
.A(n_1004),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1094),
.Y(n_1359)
);

CKINVDCx20_ASAP7_75t_R g1360 ( 
.A(n_1009),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1095),
.Y(n_1361)
);

INVxp67_ASAP7_75t_SL g1362 ( 
.A(n_1005),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_933),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_946),
.Y(n_1364)
);

INVxp33_ASAP7_75t_L g1365 ( 
.A(n_973),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1099),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_949),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1101),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_1107),
.Y(n_1369)
);

CKINVDCx20_ASAP7_75t_R g1370 ( 
.A(n_1112),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1114),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1116),
.Y(n_1372)
);

INVx3_ASAP7_75t_L g1373 ( 
.A(n_848),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1123),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1126),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_868),
.B(n_702),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1130),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_848),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1058),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_992),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_953),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_957),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1045),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_1030),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_992),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1048),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1053),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1059),
.Y(n_1388)
);

INVxp33_ASAP7_75t_SL g1389 ( 
.A(n_843),
.Y(n_1389)
);

INVxp33_ASAP7_75t_SL g1390 ( 
.A(n_1131),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1058),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1062),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1049),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1065),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1069),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1083),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1005),
.Y(n_1397)
);

INVxp67_ASAP7_75t_SL g1398 ( 
.A(n_1029),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_911),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1129),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_L g1401 ( 
.A(n_1027),
.B(n_614),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_794),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_866),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_794),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1127),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_1029),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_911),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1127),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1127),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1127),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_911),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1127),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_838),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_838),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_840),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_840),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_785),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1000),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_842),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1000),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_842),
.Y(n_1421)
);

INVxp33_ASAP7_75t_L g1422 ( 
.A(n_785),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_823),
.Y(n_1423)
);

CKINVDCx20_ASAP7_75t_R g1424 ( 
.A(n_823),
.Y(n_1424)
);

CKINVDCx16_ASAP7_75t_R g1425 ( 
.A(n_787),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1000),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_789),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_856),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_856),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_833),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_798),
.Y(n_1431)
);

CKINVDCx14_ASAP7_75t_R g1432 ( 
.A(n_866),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_938),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1081),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1173),
.B(n_1096),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1154),
.Y(n_1436)
);

AOI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1389),
.A2(n_837),
.B1(n_1046),
.B2(n_1027),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1194),
.B(n_1096),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1238),
.B(n_1096),
.Y(n_1439)
);

INVx2_ASAP7_75t_SL g1440 ( 
.A(n_1344),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1154),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1154),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1154),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1158),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1344),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1270),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1186),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1154),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1186),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1257),
.B(n_1096),
.Y(n_1450)
);

BUFx8_ASAP7_75t_L g1451 ( 
.A(n_1149),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1264),
.B(n_1115),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1390),
.B(n_1046),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1187),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1376),
.B(n_1115),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1378),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1270),
.B(n_1067),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1160),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1425),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1163),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1165),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1427),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1333),
.B(n_1067),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1274),
.B(n_1074),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1333),
.B(n_1074),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1187),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1378),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1278),
.B(n_1085),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1378),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1167),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1287),
.B(n_1085),
.Y(n_1471)
);

AND2x2_ASAP7_75t_SL g1472 ( 
.A(n_1314),
.B(n_727),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1376),
.B(n_932),
.Y(n_1473)
);

INVx4_ASAP7_75t_L g1474 ( 
.A(n_1141),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1432),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1402),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1295),
.B(n_815),
.Y(n_1477)
);

AOI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1389),
.A2(n_1139),
.B1(n_1390),
.B2(n_1342),
.Y(n_1478)
);

NOR2xp33_ASAP7_75t_SL g1479 ( 
.A(n_1230),
.B(n_490),
.Y(n_1479)
);

NAND2xp33_ASAP7_75t_L g1480 ( 
.A(n_1312),
.B(n_727),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1141),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1378),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1358),
.B(n_1362),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1153),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1404),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1245),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1397),
.B(n_1119),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1247),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1378),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1281),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1281),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1248),
.A2(n_892),
.B(n_891),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1430),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1281),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1373),
.Y(n_1495)
);

BUFx6f_ASAP7_75t_L g1496 ( 
.A(n_1373),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1373),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1139),
.A2(n_657),
.B1(n_678),
.B2(n_665),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1323),
.A2(n_1120),
.B1(n_852),
.B2(n_996),
.Y(n_1499)
);

NOR2x1_ASAP7_75t_L g1500 ( 
.A(n_1348),
.B(n_928),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1168),
.Y(n_1501)
);

AND2x6_ASAP7_75t_L g1502 ( 
.A(n_1246),
.B(n_727),
.Y(n_1502)
);

BUFx6f_ASAP7_75t_L g1503 ( 
.A(n_1412),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1135),
.Y(n_1504)
);

INVxp33_ASAP7_75t_SL g1505 ( 
.A(n_1399),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1398),
.B(n_891),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1177),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1355),
.A2(n_1200),
.B1(n_1210),
.B2(n_1292),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1249),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1412),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1137),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1138),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1405),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1178),
.B(n_932),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1406),
.B(n_892),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1352),
.Y(n_1516)
);

INVx5_ASAP7_75t_L g1517 ( 
.A(n_1149),
.Y(n_1517)
);

BUFx6f_ASAP7_75t_L g1518 ( 
.A(n_1140),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1179),
.B(n_815),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1234),
.A2(n_1120),
.B1(n_1086),
.B2(n_771),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1251),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1252),
.Y(n_1522)
);

BUFx6f_ASAP7_75t_L g1523 ( 
.A(n_1147),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1148),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1180),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1151),
.Y(n_1526)
);

INVx1_ASAP7_75t_SL g1527 ( 
.A(n_1356),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1182),
.B(n_817),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1408),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1143),
.B(n_893),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1183),
.B(n_817),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1409),
.Y(n_1532)
);

INVxp67_ASAP7_75t_L g1533 ( 
.A(n_1170),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1410),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1201),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1379),
.B(n_490),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1253),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1403),
.A2(n_1256),
.B1(n_1301),
.B2(n_1273),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1272),
.B(n_490),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1380),
.A2(n_703),
.B1(n_728),
.B2(n_688),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1155),
.B(n_893),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1222),
.B(n_896),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1184),
.Y(n_1543)
);

INVxp33_ASAP7_75t_SL g1544 ( 
.A(n_1399),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1201),
.A2(n_916),
.B(n_896),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1185),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1258),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1259),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1190),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1191),
.B(n_818),
.Y(n_1550)
);

AND2x2_ASAP7_75t_SL g1551 ( 
.A(n_1237),
.B(n_624),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1193),
.Y(n_1552)
);

AND2x6_ASAP7_75t_L g1553 ( 
.A(n_1197),
.B(n_624),
.Y(n_1553)
);

CKINVDCx20_ASAP7_75t_R g1554 ( 
.A(n_1360),
.Y(n_1554)
);

AOI22x1_ASAP7_75t_SL g1555 ( 
.A1(n_1417),
.A2(n_770),
.B1(n_684),
.B2(n_708),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1260),
.Y(n_1556)
);

AND2x4_ASAP7_75t_L g1557 ( 
.A(n_1199),
.B(n_818),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1261),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1219),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1262),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1221),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1265),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1202),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1224),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1225),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1267),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1276),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1202),
.A2(n_925),
.B(n_916),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1401),
.B(n_925),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1279),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1228),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1280),
.A2(n_937),
.B(n_929),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1283),
.B(n_929),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1285),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1345),
.A2(n_1215),
.B1(n_1391),
.B2(n_1379),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1286),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1229),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1232),
.B(n_1233),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1288),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1239),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1240),
.B(n_820),
.Y(n_1581)
);

OAI22x1_ASAP7_75t_SL g1582 ( 
.A1(n_1423),
.A2(n_684),
.B1(n_708),
.B2(n_592),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1290),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1293),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1244),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1331),
.B(n_820),
.Y(n_1586)
);

OAI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1391),
.A2(n_692),
.B1(n_928),
.B2(n_587),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1299),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1300),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1302),
.Y(n_1590)
);

AND2x2_ASAP7_75t_SL g1591 ( 
.A(n_1237),
.B(n_661),
.Y(n_1591)
);

INVx4_ASAP7_75t_L g1592 ( 
.A(n_1304),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1332),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1305),
.A2(n_952),
.B(n_937),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1407),
.B(n_490),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1306),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1337),
.B(n_821),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1308),
.Y(n_1598)
);

INVxp67_ASAP7_75t_L g1599 ( 
.A(n_1133),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1311),
.Y(n_1600)
);

AND2x6_ASAP7_75t_L g1601 ( 
.A(n_1341),
.B(n_661),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1396),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1144),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1313),
.Y(n_1604)
);

NOR2x1_ASAP7_75t_L g1605 ( 
.A(n_1269),
.B(n_668),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1343),
.B(n_821),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1203),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1316),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1203),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1317),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1319),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1325),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1327),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1433),
.B(n_822),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1328),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1212),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1396),
.Y(n_1617)
);

BUFx6f_ASAP7_75t_L g1618 ( 
.A(n_1212),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1152),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1214),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1349),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1214),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1350),
.B(n_822),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1351),
.B(n_952),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1217),
.Y(n_1625)
);

BUFx8_ASAP7_75t_SL g1626 ( 
.A(n_1172),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1357),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1272),
.A2(n_588),
.B1(n_593),
.B2(n_586),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1217),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1433),
.B(n_825),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1363),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1364),
.A2(n_1024),
.B(n_955),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1367),
.B(n_825),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1381),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1413),
.Y(n_1635)
);

BUFx6f_ASAP7_75t_L g1636 ( 
.A(n_1382),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1413),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1383),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1386),
.B(n_826),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1414),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1431),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1387),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1414),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1388),
.B(n_1392),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1394),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1395),
.Y(n_1646)
);

BUFx8_ASAP7_75t_L g1647 ( 
.A(n_1136),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1335),
.A2(n_596),
.B1(n_607),
.B2(n_605),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1400),
.A2(n_1024),
.B(n_955),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1415),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1415),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1385),
.A2(n_720),
.B1(n_592),
.B2(n_963),
.Y(n_1652)
);

BUFx12f_ASAP7_75t_L g1653 ( 
.A(n_1318),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1416),
.Y(n_1654)
);

OAI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1416),
.A2(n_1076),
.B(n_1061),
.Y(n_1655)
);

INVx4_ASAP7_75t_L g1656 ( 
.A(n_1419),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1419),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1335),
.B(n_865),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1421),
.B(n_826),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1421),
.B(n_827),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1428),
.A2(n_1076),
.B(n_1061),
.Y(n_1661)
);

BUFx6f_ASAP7_75t_L g1662 ( 
.A(n_1428),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1153),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1429),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1429),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1156),
.Y(n_1666)
);

INVxp33_ASAP7_75t_SL g1667 ( 
.A(n_1407),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_SL g1668 ( 
.A(n_1411),
.B(n_1081),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1365),
.A2(n_619),
.B1(n_620),
.B2(n_609),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1162),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1422),
.B(n_827),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1189),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1226),
.A2(n_1088),
.B(n_1084),
.Y(n_1673)
);

INVx3_ASAP7_75t_L g1674 ( 
.A(n_1157),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1231),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1243),
.B(n_828),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1241),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1296),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1411),
.B(n_1084),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1418),
.A2(n_1105),
.B(n_1088),
.Y(n_1680)
);

CKINVDCx5p33_ASAP7_75t_R g1681 ( 
.A(n_1132),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1418),
.A2(n_1113),
.B(n_1105),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1303),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1310),
.A2(n_625),
.B1(n_626),
.B2(n_622),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1157),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1420),
.B(n_828),
.Y(n_1686)
);

AND2x2_ASAP7_75t_SL g1687 ( 
.A(n_1213),
.B(n_668),
.Y(n_1687)
);

AND2x6_ASAP7_75t_L g1688 ( 
.A(n_1166),
.B(n_677),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1166),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1420),
.B(n_1113),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1175),
.Y(n_1691)
);

OAI22x1_ASAP7_75t_L g1692 ( 
.A1(n_1393),
.A2(n_963),
.B1(n_720),
.B2(n_1132),
.Y(n_1692)
);

BUFx12f_ASAP7_75t_L g1693 ( 
.A(n_1318),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1426),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1426),
.B(n_1119),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1434),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1175),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1176),
.A2(n_635),
.B1(n_640),
.B2(n_631),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1434),
.B(n_848),
.Y(n_1699)
);

INVx4_ASAP7_75t_L g1700 ( 
.A(n_1176),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1181),
.B(n_831),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1181),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1188),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1188),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1195),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1195),
.A2(n_832),
.B(n_831),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1196),
.B(n_832),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1196),
.B(n_834),
.Y(n_1708)
);

OAI22x1_ASAP7_75t_SL g1709 ( 
.A1(n_1424),
.A2(n_642),
.B1(n_643),
.B2(n_641),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1204),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1204),
.Y(n_1711)
);

BUFx6f_ASAP7_75t_L g1712 ( 
.A(n_1207),
.Y(n_1712)
);

BUFx6f_ASAP7_75t_L g1713 ( 
.A(n_1207),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1208),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1216),
.A2(n_647),
.B1(n_648),
.B2(n_646),
.Y(n_1715)
);

INVx6_ASAP7_75t_L g1716 ( 
.A(n_1318),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1142),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1208),
.B(n_871),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1220),
.A2(n_652),
.B1(n_655),
.B2(n_649),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1220),
.A2(n_664),
.B1(n_666),
.B2(n_658),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1447),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1446),
.Y(n_1722)
);

AOI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1472),
.A2(n_1346),
.B1(n_1347),
.B2(n_1340),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1676),
.B(n_1340),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1639),
.Y(n_1725)
);

INVx8_ASAP7_75t_L g1726 ( 
.A(n_1653),
.Y(n_1726)
);

AND2x4_ASAP7_75t_SL g1727 ( 
.A(n_1685),
.B(n_1134),
.Y(n_1727)
);

OAI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1508),
.A2(n_1347),
.B1(n_1353),
.B2(n_1346),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1457),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1676),
.B(n_1353),
.Y(n_1730)
);

INVx8_ASAP7_75t_L g1731 ( 
.A(n_1653),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1472),
.A2(n_1359),
.B1(n_1361),
.B2(n_1354),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1440),
.B(n_1236),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1658),
.B(n_1354),
.Y(n_1734)
);

AO22x2_ASAP7_75t_L g1735 ( 
.A1(n_1555),
.A2(n_702),
.B1(n_718),
.B2(n_704),
.Y(n_1735)
);

OA22x2_ASAP7_75t_L g1736 ( 
.A1(n_1478),
.A2(n_1366),
.B1(n_1368),
.B2(n_1361),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1655),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1551),
.A2(n_1369),
.B1(n_1371),
.B2(n_1368),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1551),
.A2(n_1371),
.B1(n_1372),
.B2(n_1369),
.Y(n_1739)
);

AO22x2_ASAP7_75t_L g1740 ( 
.A1(n_1555),
.A2(n_704),
.B1(n_729),
.B2(n_718),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1539),
.A2(n_1499),
.B1(n_1445),
.B2(n_1440),
.Y(n_1741)
);

AND2x2_ASAP7_75t_SL g1742 ( 
.A(n_1591),
.B(n_1291),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1655),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_SL g1744 ( 
.A1(n_1498),
.A2(n_1198),
.B1(n_1205),
.B2(n_1171),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1445),
.A2(n_1375),
.B1(n_1377),
.B2(n_1372),
.Y(n_1745)
);

AO22x2_ASAP7_75t_L g1746 ( 
.A1(n_1587),
.A2(n_731),
.B1(n_732),
.B2(n_729),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1447),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1591),
.A2(n_1377),
.B1(n_1375),
.B2(n_1254),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1449),
.Y(n_1749)
);

INVx8_ASAP7_75t_L g1750 ( 
.A(n_1693),
.Y(n_1750)
);

INVx4_ASAP7_75t_L g1751 ( 
.A(n_1481),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1716),
.B(n_972),
.Y(n_1752)
);

OAI22xp33_ASAP7_75t_SL g1753 ( 
.A1(n_1479),
.A2(n_1254),
.B1(n_1255),
.B2(n_1236),
.Y(n_1753)
);

AO22x2_ASAP7_75t_L g1754 ( 
.A1(n_1538),
.A2(n_732),
.B1(n_734),
.B2(n_731),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1540),
.A2(n_1652),
.B1(n_1554),
.B2(n_1145),
.Y(n_1755)
);

OAI22xp33_ASAP7_75t_L g1756 ( 
.A1(n_1437),
.A2(n_1450),
.B1(n_1533),
.B2(n_1520),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1449),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1688),
.A2(n_1268),
.B1(n_1271),
.B2(n_1255),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1473),
.B(n_1268),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_SL g1760 ( 
.A1(n_1536),
.A2(n_1275),
.B1(n_1277),
.B2(n_1271),
.Y(n_1760)
);

AO22x2_ASAP7_75t_L g1761 ( 
.A1(n_1705),
.A2(n_1714),
.B1(n_1595),
.B2(n_1617),
.Y(n_1761)
);

AO22x2_ASAP7_75t_L g1762 ( 
.A1(n_1705),
.A2(n_749),
.B1(n_766),
.B2(n_746),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1639),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1454),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1438),
.A2(n_1277),
.B1(n_1282),
.B2(n_1275),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1438),
.B(n_1282),
.Y(n_1766)
);

AO22x2_ASAP7_75t_L g1767 ( 
.A1(n_1714),
.A2(n_766),
.B1(n_706),
.B2(n_707),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1626),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_R g1769 ( 
.A(n_1681),
.B(n_1142),
.Y(n_1769)
);

OAI22xp33_ASAP7_75t_SL g1770 ( 
.A1(n_1483),
.A2(n_1289),
.B1(n_1294),
.B2(n_1284),
.Y(n_1770)
);

OAI22xp33_ASAP7_75t_SL g1771 ( 
.A1(n_1452),
.A2(n_1289),
.B1(n_1294),
.B2(n_1284),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1466),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1466),
.Y(n_1773)
);

AO22x2_ASAP7_75t_L g1774 ( 
.A1(n_1617),
.A2(n_706),
.B1(n_707),
.B2(n_677),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1457),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1481),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1586),
.Y(n_1777)
);

OA22x2_ASAP7_75t_L g1778 ( 
.A1(n_1575),
.A2(n_1307),
.B1(n_1309),
.B2(n_1297),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1688),
.A2(n_1307),
.B1(n_1309),
.B2(n_1297),
.Y(n_1779)
);

INVx4_ASAP7_75t_L g1780 ( 
.A(n_1481),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1473),
.B(n_1315),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1659),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1446),
.B(n_938),
.Y(n_1783)
);

XNOR2xp5_ASAP7_75t_L g1784 ( 
.A(n_1554),
.B(n_1159),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1618),
.Y(n_1785)
);

AOI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1688),
.A2(n_1322),
.B1(n_1324),
.B2(n_1315),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1438),
.B(n_1322),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1688),
.A2(n_1330),
.B1(n_1336),
.B2(n_1324),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1459),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1661),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1527),
.B(n_1462),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1671),
.B(n_1330),
.Y(n_1792)
);

OAI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1679),
.A2(n_1338),
.B1(n_1336),
.B2(n_1384),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1618),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1688),
.A2(n_1338),
.B1(n_1223),
.B2(n_1235),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1661),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1671),
.B(n_1081),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1618),
.Y(n_1798)
);

AO22x2_ASAP7_75t_L g1799 ( 
.A1(n_1669),
.A2(n_1720),
.B1(n_1719),
.B2(n_1703),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1453),
.B(n_1227),
.Y(n_1800)
);

AOI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1688),
.A2(n_1242),
.B1(n_1263),
.B2(n_1250),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1545),
.Y(n_1802)
);

AO22x2_ASAP7_75t_L g1803 ( 
.A1(n_1689),
.A2(n_751),
.B1(n_760),
.B2(n_750),
.Y(n_1803)
);

OAI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1690),
.A2(n_1695),
.B1(n_1517),
.B2(n_1464),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1545),
.Y(n_1805)
);

OA22x2_ASAP7_75t_L g1806 ( 
.A1(n_1715),
.A2(n_1393),
.B1(n_671),
.B2(n_676),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1502),
.A2(n_1266),
.B1(n_1320),
.B2(n_1298),
.Y(n_1807)
);

OAI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1517),
.A2(n_751),
.B1(n_760),
.B2(n_750),
.Y(n_1808)
);

OAI22xp33_ASAP7_75t_SL g1809 ( 
.A1(n_1468),
.A2(n_1150),
.B1(n_1146),
.B2(n_680),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1618),
.Y(n_1810)
);

OR2x6_ASAP7_75t_L g1811 ( 
.A(n_1716),
.B(n_940),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1502),
.A2(n_1321),
.B1(n_1329),
.B2(n_1326),
.Y(n_1812)
);

OR2x6_ASAP7_75t_L g1813 ( 
.A(n_1716),
.B(n_940),
.Y(n_1813)
);

XOR2xp5_ASAP7_75t_L g1814 ( 
.A(n_1516),
.B(n_1161),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1502),
.A2(n_1334),
.B1(n_1339),
.B2(n_1370),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1462),
.B(n_1146),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1455),
.B(n_1374),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1502),
.A2(n_1218),
.B1(n_1150),
.B2(n_1169),
.Y(n_1818)
);

AO22x2_ASAP7_75t_L g1819 ( 
.A1(n_1689),
.A2(n_942),
.B1(n_943),
.B2(n_941),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1708),
.B(n_462),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1618),
.Y(n_1821)
);

OR2x6_ASAP7_75t_L g1822 ( 
.A(n_1716),
.B(n_941),
.Y(n_1822)
);

NAND2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1694),
.B(n_670),
.Y(n_1823)
);

OAI22xp33_ASAP7_75t_SL g1824 ( 
.A1(n_1718),
.A2(n_683),
.B1(n_689),
.B2(n_681),
.Y(n_1824)
);

OAI22xp33_ASAP7_75t_R g1825 ( 
.A1(n_1582),
.A2(n_1602),
.B1(n_942),
.B2(n_944),
.Y(n_1825)
);

BUFx6f_ASAP7_75t_L g1826 ( 
.A(n_1457),
.Y(n_1826)
);

NAND3x1_ASAP7_75t_L g1827 ( 
.A(n_1674),
.B(n_944),
.C(n_943),
.Y(n_1827)
);

OAI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1684),
.A2(n_691),
.B1(n_693),
.B2(n_690),
.Y(n_1828)
);

AO22x2_ASAP7_75t_L g1829 ( 
.A1(n_1703),
.A2(n_1702),
.B1(n_1670),
.B2(n_1675),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1650),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_R g1831 ( 
.A1(n_1641),
.A2(n_959),
.B1(n_964),
.B2(n_945),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1439),
.B(n_871),
.Y(n_1832)
);

OA22x2_ASAP7_75t_L g1833 ( 
.A1(n_1698),
.A2(n_698),
.B1(n_699),
.B2(n_696),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1708),
.B(n_531),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1701),
.B(n_531),
.Y(n_1835)
);

AO22x2_ASAP7_75t_L g1836 ( 
.A1(n_1666),
.A2(n_959),
.B1(n_964),
.B2(n_945),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1568),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1502),
.A2(n_1164),
.B1(n_711),
.B2(n_712),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1500),
.B(n_1206),
.Y(n_1839)
);

OA22x2_ASAP7_75t_L g1840 ( 
.A1(n_1628),
.A2(n_713),
.B1(n_714),
.B2(n_705),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1568),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1650),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1701),
.B(n_1707),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1502),
.A2(n_722),
.B1(n_726),
.B2(n_715),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1632),
.Y(n_1845)
);

OA22x2_ASAP7_75t_L g1846 ( 
.A1(n_1648),
.A2(n_736),
.B1(n_737),
.B2(n_730),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1621),
.A2(n_742),
.B1(n_745),
.B2(n_738),
.Y(n_1847)
);

INVxp67_ASAP7_75t_SL g1848 ( 
.A(n_1650),
.Y(n_1848)
);

OAI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1627),
.A2(n_752),
.B1(n_755),
.B2(n_747),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1650),
.Y(n_1850)
);

OAI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1645),
.A2(n_758),
.B1(n_759),
.B2(n_756),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1701),
.A2(n_762),
.B1(n_764),
.B2(n_761),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1707),
.A2(n_767),
.B1(n_768),
.B2(n_765),
.Y(n_1853)
);

OR2x2_ASAP7_75t_L g1854 ( 
.A(n_1493),
.B(n_967),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1463),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1707),
.B(n_1686),
.Y(n_1856)
);

AOI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1439),
.A2(n_769),
.B1(n_836),
.B2(n_834),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1514),
.B(n_531),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1439),
.B(n_1477),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1477),
.B(n_871),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1514),
.B(n_531),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1659),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1471),
.A2(n_839),
.B1(n_841),
.B2(n_836),
.Y(n_1863)
);

OAI22xp5_ASAP7_75t_L g1864 ( 
.A1(n_1435),
.A2(n_841),
.B1(n_844),
.B2(n_839),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1586),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1471),
.B(n_1209),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1471),
.A2(n_845),
.B1(n_847),
.B2(n_844),
.Y(n_1867)
);

OAI22xp33_ASAP7_75t_SL g1868 ( 
.A1(n_1644),
.A2(n_968),
.B1(n_975),
.B2(n_967),
.Y(n_1868)
);

INVx2_ASAP7_75t_L g1869 ( 
.A(n_1650),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1692),
.A2(n_1211),
.B1(n_1192),
.B2(n_1174),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1706),
.A2(n_847),
.B1(n_850),
.B2(n_845),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1517),
.B(n_549),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1477),
.B(n_1487),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1706),
.A2(n_851),
.B1(n_853),
.B2(n_850),
.Y(n_1874)
);

OAI22xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1666),
.A2(n_975),
.B1(n_978),
.B2(n_968),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1706),
.A2(n_853),
.B1(n_854),
.B2(n_851),
.Y(n_1876)
);

AO22x2_ASAP7_75t_L g1877 ( 
.A1(n_1670),
.A2(n_979),
.B1(n_980),
.B2(n_978),
.Y(n_1877)
);

OAI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1517),
.A2(n_855),
.B1(n_858),
.B2(n_854),
.Y(n_1878)
);

AO22x2_ASAP7_75t_L g1879 ( 
.A1(n_1675),
.A2(n_980),
.B1(n_981),
.B2(n_979),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1463),
.B(n_981),
.Y(n_1880)
);

OAI22xp33_ASAP7_75t_SL g1881 ( 
.A1(n_1699),
.A2(n_984),
.B1(n_985),
.B2(n_982),
.Y(n_1881)
);

OR2x6_ASAP7_75t_L g1882 ( 
.A(n_1685),
.B(n_982),
.Y(n_1882)
);

INVx3_ASAP7_75t_L g1883 ( 
.A(n_1659),
.Y(n_1883)
);

INVx2_ASAP7_75t_L g1884 ( 
.A(n_1654),
.Y(n_1884)
);

CKINVDCx20_ASAP7_75t_R g1885 ( 
.A(n_1647),
.Y(n_1885)
);

OAI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1517),
.A2(n_858),
.B1(n_867),
.B2(n_855),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1463),
.B(n_549),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1686),
.B(n_549),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1686),
.A2(n_870),
.B1(n_872),
.B2(n_867),
.Y(n_1889)
);

OAI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1444),
.A2(n_872),
.B1(n_873),
.B2(n_870),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1654),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1654),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1654),
.Y(n_1893)
);

AO22x2_ASAP7_75t_L g1894 ( 
.A1(n_1672),
.A2(n_988),
.B1(n_999),
.B2(n_987),
.Y(n_1894)
);

OAI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1444),
.A2(n_873),
.B1(n_999),
.B2(n_988),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1654),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1662),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1687),
.A2(n_1002),
.B1(n_1007),
.B2(n_1001),
.Y(n_1898)
);

AO22x2_ASAP7_75t_L g1899 ( 
.A1(n_1677),
.A2(n_1002),
.B1(n_1007),
.B2(n_1001),
.Y(n_1899)
);

AND2x2_ASAP7_75t_SL g1900 ( 
.A(n_1687),
.B(n_1493),
.Y(n_1900)
);

OR2x6_ASAP7_75t_L g1901 ( 
.A(n_1685),
.B(n_1128),
.Y(n_1901)
);

BUFx10_ASAP7_75t_L g1902 ( 
.A(n_1685),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1677),
.B(n_549),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1578),
.A2(n_1011),
.B1(n_1012),
.B2(n_1008),
.Y(n_1904)
);

AO22x2_ASAP7_75t_L g1905 ( 
.A1(n_1683),
.A2(n_1678),
.B1(n_1710),
.B2(n_1674),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1632),
.Y(n_1906)
);

AOI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1578),
.A2(n_1011),
.B1(n_1012),
.B2(n_1008),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1692),
.A2(n_1017),
.B1(n_1022),
.B2(n_1013),
.Y(n_1908)
);

CKINVDCx6p67_ASAP7_75t_R g1909 ( 
.A(n_1693),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1632),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1465),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1578),
.A2(n_1128),
.B1(n_1017),
.B2(n_1022),
.Y(n_1912)
);

AOI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1480),
.A2(n_1025),
.B1(n_1028),
.B2(n_1013),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1662),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1597),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_SL g1916 ( 
.A1(n_1681),
.A2(n_1028),
.B1(n_1035),
.B2(n_1025),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1597),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1501),
.A2(n_1037),
.B1(n_1039),
.B2(n_1035),
.Y(n_1918)
);

OAI22xp33_ASAP7_75t_SL g1919 ( 
.A1(n_1683),
.A2(n_1039),
.B1(n_1042),
.B2(n_1037),
.Y(n_1919)
);

INVx5_ASAP7_75t_L g1920 ( 
.A(n_1601),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1662),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1649),
.Y(n_1922)
);

OAI22xp33_ASAP7_75t_SL g1923 ( 
.A1(n_1674),
.A2(n_1052),
.B1(n_1071),
.B2(n_1042),
.Y(n_1923)
);

INVx8_ASAP7_75t_L g1924 ( 
.A(n_1685),
.Y(n_1924)
);

XNOR2xp5_ASAP7_75t_L g1925 ( 
.A(n_1484),
.B(n_271),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1480),
.A2(n_1071),
.B1(n_1072),
.B2(n_1052),
.Y(n_1926)
);

OA22x2_ASAP7_75t_L g1927 ( 
.A1(n_1668),
.A2(n_1696),
.B1(n_1603),
.B2(n_1619),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1662),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1597),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1710),
.B(n_1465),
.Y(n_1930)
);

OAI22xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1710),
.A2(n_1073),
.B1(n_1075),
.B2(n_1072),
.Y(n_1931)
);

OAI22xp33_ASAP7_75t_L g1932 ( 
.A1(n_1501),
.A2(n_1075),
.B1(n_1077),
.B2(n_1073),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1606),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1465),
.A2(n_1125),
.B1(n_1079),
.B2(n_1087),
.Y(n_1934)
);

OAI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1592),
.A2(n_1079),
.B1(n_1087),
.B2(n_1077),
.Y(n_1935)
);

OAI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1507),
.A2(n_1561),
.B1(n_1564),
.B2(n_1525),
.Y(n_1936)
);

OR2x6_ASAP7_75t_L g1937 ( 
.A(n_1691),
.B(n_1089),
.Y(n_1937)
);

OAI22xp33_ASAP7_75t_SL g1938 ( 
.A1(n_1593),
.A2(n_1090),
.B1(n_1092),
.B2(n_1089),
.Y(n_1938)
);

AOI22xp5_ASAP7_75t_L g1939 ( 
.A1(n_1593),
.A2(n_1125),
.B1(n_1092),
.B2(n_1093),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1599),
.B(n_610),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1649),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1662),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1475),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1631),
.A2(n_1124),
.B1(n_1093),
.B2(n_1097),
.Y(n_1944)
);

AO22x2_ASAP7_75t_L g1945 ( 
.A1(n_1697),
.A2(n_1097),
.B1(n_1098),
.B2(n_1090),
.Y(n_1945)
);

AO22x2_ASAP7_75t_L g1946 ( 
.A1(n_1697),
.A2(n_1100),
.B1(n_1103),
.B2(n_1098),
.Y(n_1946)
);

OAI22xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1631),
.A2(n_1103),
.B1(n_1104),
.B2(n_1100),
.Y(n_1947)
);

AO22x2_ASAP7_75t_L g1948 ( 
.A1(n_1700),
.A2(n_1106),
.B1(n_1108),
.B2(n_1104),
.Y(n_1948)
);

AO22x2_ASAP7_75t_L g1949 ( 
.A1(n_1700),
.A2(n_1108),
.B1(n_1109),
.B2(n_1106),
.Y(n_1949)
);

OR2x6_ASAP7_75t_L g1950 ( 
.A(n_1691),
.B(n_1109),
.Y(n_1950)
);

AOI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1458),
.A2(n_1124),
.B1(n_1111),
.B2(n_1117),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1460),
.A2(n_1111),
.B1(n_1117),
.B2(n_1110),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1505),
.B(n_1544),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1700),
.B(n_610),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1649),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1691),
.B(n_610),
.Y(n_1956)
);

OAI22xp33_ASAP7_75t_SL g1957 ( 
.A1(n_1506),
.A2(n_1118),
.B1(n_1121),
.B2(n_1110),
.Y(n_1957)
);

AO22x2_ASAP7_75t_L g1958 ( 
.A1(n_1507),
.A2(n_1121),
.B1(n_1122),
.B2(n_1118),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1635),
.Y(n_1959)
);

AOI22x1_ASAP7_75t_SL g1960 ( 
.A1(n_1717),
.A2(n_1484),
.B1(n_1663),
.B2(n_1709),
.Y(n_1960)
);

OA22x2_ASAP7_75t_L g1961 ( 
.A1(n_1663),
.A2(n_1122),
.B1(n_639),
.B2(n_723),
.Y(n_1961)
);

OAI22xp33_ASAP7_75t_L g1962 ( 
.A1(n_1525),
.A2(n_1564),
.B1(n_1565),
.B2(n_1561),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1616),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1616),
.Y(n_1964)
);

OAI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1565),
.A2(n_1047),
.B1(n_997),
.B2(n_1019),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1592),
.A2(n_997),
.B1(n_1019),
.B2(n_871),
.Y(n_1966)
);

OAI22xp33_ASAP7_75t_SL g1967 ( 
.A1(n_1515),
.A2(n_639),
.B1(n_723),
.B2(n_612),
.Y(n_1967)
);

XNOR2xp5_ASAP7_75t_L g1968 ( 
.A(n_1717),
.B(n_272),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1691),
.B(n_612),
.Y(n_1969)
);

OA22x2_ASAP7_75t_L g1970 ( 
.A1(n_1571),
.A2(n_639),
.B1(n_723),
.B2(n_612),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1635),
.Y(n_1971)
);

OAI22xp33_ASAP7_75t_L g1972 ( 
.A1(n_1571),
.A2(n_1580),
.B1(n_1585),
.B2(n_1577),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1505),
.B(n_612),
.Y(n_1973)
);

AO22x2_ASAP7_75t_L g1974 ( 
.A1(n_1577),
.A2(n_723),
.B1(n_639),
.B2(n_8),
.Y(n_1974)
);

AO22x2_ASAP7_75t_L g1975 ( 
.A1(n_1580),
.A2(n_9),
.B1(n_6),
.B2(n_7),
.Y(n_1975)
);

OAI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1585),
.A2(n_1047),
.B1(n_997),
.B2(n_1019),
.Y(n_1976)
);

AO22x2_ASAP7_75t_L g1977 ( 
.A1(n_1461),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1977)
);

XNOR2xp5_ASAP7_75t_L g1978 ( 
.A(n_1544),
.B(n_275),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1635),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1470),
.A2(n_997),
.B1(n_1019),
.B2(n_871),
.Y(n_1980)
);

AND2x4_ASAP7_75t_L g1981 ( 
.A(n_1543),
.B(n_1546),
.Y(n_1981)
);

AOI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1549),
.A2(n_1019),
.B1(n_1040),
.B2(n_997),
.Y(n_1982)
);

AOI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1552),
.A2(n_1047),
.B1(n_1040),
.B2(n_278),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1691),
.B(n_1040),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1704),
.B(n_1040),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1667),
.B(n_1559),
.Y(n_1986)
);

OAI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1542),
.A2(n_1047),
.B1(n_1040),
.B2(n_14),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1637),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1592),
.B(n_1047),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1637),
.Y(n_1990)
);

OAI22xp33_ASAP7_75t_SL g1991 ( 
.A1(n_1667),
.A2(n_15),
.B1(n_11),
.B2(n_13),
.Y(n_1991)
);

INVx2_ASAP7_75t_SL g1992 ( 
.A(n_1605),
.Y(n_1992)
);

OAI22xp33_ASAP7_75t_SL g1993 ( 
.A1(n_1590),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1713),
.B(n_18),
.Y(n_1994)
);

AOI22xp5_ASAP7_75t_L g1995 ( 
.A1(n_1601),
.A2(n_1636),
.B1(n_1638),
.B2(n_1634),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1606),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1606),
.Y(n_1997)
);

INVx5_ASAP7_75t_L g1998 ( 
.A(n_1601),
.Y(n_1998)
);

OAI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1704),
.A2(n_1712),
.B1(n_1713),
.B2(n_1711),
.Y(n_1999)
);

AND2x2_ASAP7_75t_SL g2000 ( 
.A(n_1704),
.B(n_20),
.Y(n_2000)
);

OAI22xp33_ASAP7_75t_SL g2001 ( 
.A1(n_1590),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_2001)
);

AOI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1601),
.A2(n_1636),
.B1(n_1638),
.B2(n_1634),
.Y(n_2002)
);

OAI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1713),
.A2(n_1711),
.B1(n_1712),
.B2(n_1704),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1637),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1963),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1963),
.Y(n_2006)
);

OR2x6_ASAP7_75t_L g2007 ( 
.A(n_1924),
.B(n_1704),
.Y(n_2007)
);

OAI22xp5_ASAP7_75t_L g2008 ( 
.A1(n_1859),
.A2(n_1712),
.B1(n_1713),
.B2(n_1711),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1734),
.B(n_1711),
.Y(n_2009)
);

AOI22xp33_ASAP7_75t_L g2010 ( 
.A1(n_1782),
.A2(n_1553),
.B1(n_1601),
.B2(n_1656),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1964),
.Y(n_2011)
);

NOR2xp33_ASAP7_75t_L g2012 ( 
.A(n_1792),
.B(n_1724),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1789),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1826),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1782),
.A2(n_1553),
.B1(n_1601),
.B2(n_1656),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1882),
.Y(n_2016)
);

AND2x6_ASAP7_75t_L g2017 ( 
.A(n_1845),
.B(n_1711),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1964),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1845),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1999),
.B(n_1712),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_1769),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1873),
.B(n_1608),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1906),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1906),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1910),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1910),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1922),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1902),
.Y(n_2028)
);

INVx2_ASAP7_75t_L g2029 ( 
.A(n_1922),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1941),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1902),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_2003),
.B(n_1712),
.Y(n_2032)
);

NOR2x1p5_ASAP7_75t_L g2033 ( 
.A(n_1909),
.B(n_1713),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1959),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1741),
.B(n_1634),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1862),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1862),
.Y(n_2037)
);

XOR2x2_ASAP7_75t_SL g2038 ( 
.A(n_1898),
.B(n_1451),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1930),
.B(n_1612),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1883),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1924),
.B(n_1673),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1722),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1883),
.Y(n_2043)
);

INVx4_ASAP7_75t_L g2044 ( 
.A(n_1751),
.Y(n_2044)
);

BUFx3_ASAP7_75t_L g2045 ( 
.A(n_1722),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1797),
.B(n_1612),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1941),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1826),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1971),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1979),
.Y(n_2050)
);

INVx4_ASAP7_75t_SL g2051 ( 
.A(n_1955),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1988),
.Y(n_2052)
);

NOR2xp33_ASAP7_75t_L g2053 ( 
.A(n_1730),
.B(n_1647),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1936),
.B(n_1613),
.Y(n_2054)
);

NAND2xp33_ASAP7_75t_L g2055 ( 
.A(n_1920),
.B(n_1553),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1990),
.Y(n_2056)
);

INVx4_ASAP7_75t_SL g2057 ( 
.A(n_1955),
.Y(n_2057)
);

INVx8_ASAP7_75t_L g2058 ( 
.A(n_1882),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2004),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1777),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_1800),
.B(n_1647),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1865),
.Y(n_2062)
);

AND2x4_ASAP7_75t_L g2063 ( 
.A(n_1729),
.B(n_1623),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1843),
.B(n_1634),
.Y(n_2064)
);

AOI22xp5_ASAP7_75t_L g2065 ( 
.A1(n_1759),
.A2(n_1636),
.B1(n_1638),
.B2(n_1634),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1962),
.B(n_1613),
.Y(n_2066)
);

NAND2xp33_ASAP7_75t_L g2067 ( 
.A(n_1920),
.B(n_1553),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1802),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1802),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1805),
.Y(n_2070)
);

INVx4_ASAP7_75t_L g2071 ( 
.A(n_1751),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1805),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1915),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1837),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1972),
.B(n_1725),
.Y(n_2075)
);

INVx4_ASAP7_75t_L g2076 ( 
.A(n_1776),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1917),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1826),
.B(n_1623),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1804),
.B(n_1636),
.Y(n_2079)
);

INVx4_ASAP7_75t_L g2080 ( 
.A(n_1776),
.Y(n_2080)
);

NOR3xp33_ASAP7_75t_L g2081 ( 
.A(n_1728),
.B(n_1856),
.C(n_1793),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1763),
.B(n_1680),
.Y(n_2082)
);

AOI22xp33_ASAP7_75t_L g2083 ( 
.A1(n_2000),
.A2(n_1553),
.B1(n_1656),
.B2(n_1680),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1929),
.B(n_1615),
.Y(n_2084)
);

INVx5_ASAP7_75t_L g2085 ( 
.A(n_1920),
.Y(n_2085)
);

INVxp33_ASAP7_75t_SL g2086 ( 
.A(n_1784),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1933),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_1781),
.A2(n_1638),
.B1(n_1642),
.B2(n_1636),
.Y(n_2088)
);

BUFx6f_ASAP7_75t_L g2089 ( 
.A(n_1998),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_1837),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1785),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_1996),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1820),
.B(n_1680),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1997),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1841),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1834),
.B(n_1682),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_1903),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1998),
.B(n_1638),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1841),
.Y(n_2099)
);

INVx3_ASAP7_75t_L g2100 ( 
.A(n_1794),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_1798),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1737),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1956),
.B(n_1969),
.Y(n_2103)
);

INVx6_ASAP7_75t_L g2104 ( 
.A(n_1780),
.Y(n_2104)
);

NAND2xp33_ASAP7_75t_L g2105 ( 
.A(n_1998),
.B(n_1995),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1880),
.B(n_1615),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1880),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1721),
.Y(n_2108)
);

OAI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1723),
.A2(n_1646),
.B1(n_1642),
.B2(n_1682),
.Y(n_2109)
);

HB1xp67_ASAP7_75t_L g2110 ( 
.A(n_1901),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1858),
.B(n_1682),
.Y(n_2111)
);

BUFx3_ASAP7_75t_L g2112 ( 
.A(n_1722),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1985),
.B(n_1642),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_1791),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1747),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_1854),
.B(n_1816),
.Y(n_2116)
);

BUFx10_ASAP7_75t_L g2117 ( 
.A(n_1953),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1766),
.B(n_1642),
.Y(n_2118)
);

AND2x2_ASAP7_75t_SL g2119 ( 
.A(n_1742),
.B(n_1474),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1737),
.Y(n_2120)
);

NAND2xp33_ASAP7_75t_L g2121 ( 
.A(n_2002),
.B(n_1553),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_1787),
.B(n_1642),
.Y(n_2122)
);

BUFx2_ASAP7_75t_L g2123 ( 
.A(n_1817),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1743),
.Y(n_2124)
);

AND2x6_ASAP7_75t_L g2125 ( 
.A(n_1743),
.B(n_1535),
.Y(n_2125)
);

INVx5_ASAP7_75t_L g2126 ( 
.A(n_1901),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1790),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1790),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1749),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_1872),
.B(n_1646),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1796),
.Y(n_2131)
);

NAND3xp33_ASAP7_75t_L g2132 ( 
.A(n_1973),
.B(n_1451),
.C(n_1646),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1796),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_1733),
.B(n_1646),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1757),
.Y(n_2135)
);

BUFx3_ASAP7_75t_L g2136 ( 
.A(n_1727),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_1810),
.Y(n_2137)
);

AOI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1799),
.A2(n_1504),
.B1(n_1486),
.B2(n_1488),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1764),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1772),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1773),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1821),
.Y(n_2142)
);

INVx1_ASAP7_75t_SL g2143 ( 
.A(n_1943),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1981),
.B(n_1783),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1981),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1783),
.B(n_1535),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1756),
.A2(n_1504),
.B1(n_1509),
.B2(n_1486),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_L g2148 ( 
.A(n_1780),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1830),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_1814),
.Y(n_2150)
);

AND2x4_ASAP7_75t_L g2151 ( 
.A(n_1775),
.B(n_1623),
.Y(n_2151)
);

INVx4_ASAP7_75t_L g2152 ( 
.A(n_1937),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1745),
.B(n_1535),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1842),
.Y(n_2154)
);

INVx4_ASAP7_75t_L g2155 ( 
.A(n_1937),
.Y(n_2155)
);

NOR3xp33_ASAP7_75t_L g2156 ( 
.A(n_1765),
.B(n_1624),
.C(n_1519),
.Y(n_2156)
);

INVx2_ASAP7_75t_L g2157 ( 
.A(n_1850),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1894),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_1950),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1869),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_1884),
.Y(n_2161)
);

BUFx6f_ASAP7_75t_L g2162 ( 
.A(n_1855),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_1892),
.Y(n_2163)
);

BUFx6f_ASAP7_75t_L g2164 ( 
.A(n_1911),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1893),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1861),
.B(n_1563),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_1896),
.Y(n_2167)
);

BUFx8_ASAP7_75t_SL g2168 ( 
.A(n_1768),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1986),
.B(n_1451),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1894),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_SL g2171 ( 
.A(n_1758),
.B(n_1563),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_1819),
.B(n_1614),
.Y(n_2172)
);

BUFx3_ASAP7_75t_L g2173 ( 
.A(n_1726),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_SL g2174 ( 
.A(n_1779),
.B(n_1563),
.Y(n_2174)
);

BUFx10_ASAP7_75t_L g2175 ( 
.A(n_1866),
.Y(n_2175)
);

NAND2xp33_ASAP7_75t_L g2176 ( 
.A(n_1827),
.B(n_1607),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_1897),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1786),
.B(n_1607),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1788),
.B(n_1607),
.Y(n_2179)
);

AND2x4_ASAP7_75t_L g2180 ( 
.A(n_1994),
.B(n_1633),
.Y(n_2180)
);

HB1xp67_ASAP7_75t_L g2181 ( 
.A(n_1950),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_1732),
.B(n_1738),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1899),
.Y(n_2183)
);

AND2x2_ASAP7_75t_SL g2184 ( 
.A(n_1900),
.B(n_1474),
.Y(n_2184)
);

INVx2_ASAP7_75t_SL g2185 ( 
.A(n_1905),
.Y(n_2185)
);

BUFx2_ASAP7_75t_L g2186 ( 
.A(n_1752),
.Y(n_2186)
);

NOR2xp33_ASAP7_75t_L g2187 ( 
.A(n_1739),
.B(n_1504),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1914),
.Y(n_2188)
);

INVx8_ASAP7_75t_L g2189 ( 
.A(n_1811),
.Y(n_2189)
);

INVx5_ASAP7_75t_L g2190 ( 
.A(n_1811),
.Y(n_2190)
);

INVx2_ASAP7_75t_SL g2191 ( 
.A(n_1905),
.Y(n_2191)
);

OR2x6_ASAP7_75t_L g2192 ( 
.A(n_1813),
.B(n_1673),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1748),
.B(n_1609),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1921),
.Y(n_2194)
);

INVx1_ASAP7_75t_SL g2195 ( 
.A(n_1916),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_SL g2196 ( 
.A(n_1760),
.B(n_1609),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1928),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1942),
.Y(n_2198)
);

INVx3_ASAP7_75t_L g2199 ( 
.A(n_1832),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_SL g2200 ( 
.A(n_1824),
.B(n_1609),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1819),
.B(n_1614),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1899),
.Y(n_2202)
);

NOR2xp33_ASAP7_75t_L g2203 ( 
.A(n_1839),
.B(n_1474),
.Y(n_2203)
);

INVx5_ASAP7_75t_L g2204 ( 
.A(n_1813),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1860),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1958),
.Y(n_2206)
);

INVx5_ASAP7_75t_L g2207 ( 
.A(n_1822),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_L g2208 ( 
.A(n_1888),
.B(n_1521),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1958),
.Y(n_2209)
);

BUFx10_ASAP7_75t_L g2210 ( 
.A(n_1940),
.Y(n_2210)
);

BUFx6f_ASAP7_75t_L g2211 ( 
.A(n_1822),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1989),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1863),
.Y(n_2213)
);

AND2x6_ASAP7_75t_L g2214 ( 
.A(n_1871),
.B(n_1620),
.Y(n_2214)
);

INVxp33_ASAP7_75t_SL g2215 ( 
.A(n_1744),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1848),
.B(n_1521),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1867),
.Y(n_2217)
);

NAND2xp33_ASAP7_75t_R g2218 ( 
.A(n_1954),
.B(n_1633),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1829),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1891),
.B(n_1522),
.Y(n_2220)
);

NAND3xp33_ASAP7_75t_L g2221 ( 
.A(n_1852),
.B(n_1519),
.C(n_1633),
.Y(n_2221)
);

AND2x2_ASAP7_75t_L g2222 ( 
.A(n_1835),
.B(n_1630),
.Y(n_2222)
);

BUFx3_ASAP7_75t_L g2223 ( 
.A(n_1726),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1992),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1829),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1874),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1876),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1803),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1803),
.Y(n_2229)
);

INVx2_ASAP7_75t_SL g2230 ( 
.A(n_1836),
.Y(n_2230)
);

INVx2_ASAP7_75t_SL g2231 ( 
.A(n_1836),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1877),
.Y(n_2232)
);

INVx1_ASAP7_75t_SL g2233 ( 
.A(n_1752),
.Y(n_2233)
);

INVx4_ASAP7_75t_L g2234 ( 
.A(n_1945),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_1795),
.B(n_1522),
.Y(n_2235)
);

NAND2xp33_ASAP7_75t_R g2236 ( 
.A(n_1960),
.B(n_1528),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1877),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_1761),
.A2(n_1548),
.B1(n_1556),
.B2(n_1537),
.Y(n_2238)
);

AND2x6_ASAP7_75t_L g2239 ( 
.A(n_1887),
.B(n_1620),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1935),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_1879),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1864),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_1984),
.Y(n_2243)
);

NOR2xp33_ASAP7_75t_L g2244 ( 
.A(n_1838),
.B(n_1537),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1879),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_SL g2246 ( 
.A(n_1923),
.B(n_1503),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1881),
.B(n_1548),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_1904),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1774),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1907),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1912),
.Y(n_2251)
);

BUFx3_ASAP7_75t_L g2252 ( 
.A(n_1731),
.Y(n_2252)
);

BUFx10_ASAP7_75t_L g2253 ( 
.A(n_1831),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_1945),
.B(n_1630),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_1946),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_1840),
.A2(n_1556),
.B1(n_1562),
.B2(n_1560),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_1931),
.B(n_1503),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_1889),
.B(n_1560),
.Y(n_2258)
);

INVx5_ASAP7_75t_L g2259 ( 
.A(n_1731),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1774),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1938),
.Y(n_2261)
);

OR2x2_ASAP7_75t_L g2262 ( 
.A(n_1818),
.B(n_1528),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1947),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1934),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1828),
.B(n_1503),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_SL g2266 ( 
.A(n_1770),
.B(n_1503),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_1750),
.Y(n_2267)
);

INVx3_ASAP7_75t_L g2268 ( 
.A(n_1946),
.Y(n_2268)
);

INVx1_ASAP7_75t_SL g2269 ( 
.A(n_1823),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1913),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1957),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1939),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_1771),
.B(n_1503),
.Y(n_2273)
);

INVx2_ASAP7_75t_SL g2274 ( 
.A(n_1948),
.Y(n_2274)
);

BUFx2_ASAP7_75t_L g2275 ( 
.A(n_1948),
.Y(n_2275)
);

NAND2xp33_ASAP7_75t_L g2276 ( 
.A(n_1761),
.B(n_1510),
.Y(n_2276)
);

INVx2_ASAP7_75t_SL g2277 ( 
.A(n_1949),
.Y(n_2277)
);

INVx8_ASAP7_75t_L g2278 ( 
.A(n_1750),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_1944),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_L g2280 ( 
.A(n_1807),
.B(n_1562),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_1949),
.B(n_1528),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1919),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1926),
.Y(n_2283)
);

INVx5_ASAP7_75t_L g2284 ( 
.A(n_1878),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1754),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1875),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_1908),
.Y(n_2287)
);

INVx3_ASAP7_75t_L g2288 ( 
.A(n_1927),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_SL g2289 ( 
.A(n_1753),
.B(n_1844),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_SL g2290 ( 
.A(n_1857),
.B(n_1510),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2005),
.Y(n_2291)
);

INVx1_ASAP7_75t_SL g2292 ( 
.A(n_2143),
.Y(n_2292)
);

BUFx6f_ASAP7_75t_L g2293 ( 
.A(n_2014),
.Y(n_2293)
);

AO22x2_ASAP7_75t_L g2294 ( 
.A1(n_2229),
.A2(n_1975),
.B1(n_1977),
.B2(n_1974),
.Y(n_2294)
);

CKINVDCx20_ASAP7_75t_R g2295 ( 
.A(n_2168),
.Y(n_2295)
);

NAND2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2126),
.B(n_1664),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2005),
.Y(n_2297)
);

CKINVDCx20_ASAP7_75t_R g2298 ( 
.A(n_2168),
.Y(n_2298)
);

INVx1_ASAP7_75t_SL g2299 ( 
.A(n_2013),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_2014),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2104),
.Y(n_2301)
);

AND2x4_ASAP7_75t_L g2302 ( 
.A(n_2042),
.B(n_1812),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2006),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2006),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2068),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2011),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2012),
.B(n_1815),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2018),
.Y(n_2308)
);

INVx3_ASAP7_75t_L g2309 ( 
.A(n_2104),
.Y(n_2309)
);

NAND2x1p5_ASAP7_75t_L g2310 ( 
.A(n_2126),
.B(n_1664),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2139),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_2103),
.B(n_1801),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2185),
.Y(n_2313)
);

INVx2_ASAP7_75t_L g2314 ( 
.A(n_2139),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_L g2315 ( 
.A(n_2116),
.B(n_1809),
.Y(n_2315)
);

AND2x4_ASAP7_75t_L g2316 ( 
.A(n_2042),
.B(n_2045),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_2222),
.B(n_2116),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_2195),
.B(n_2097),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_2068),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2069),
.Y(n_2320)
);

CKINVDCx5p33_ASAP7_75t_R g2321 ( 
.A(n_2021),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2182),
.A2(n_1736),
.B1(n_1778),
.B2(n_1846),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2069),
.Y(n_2323)
);

INVxp67_ASAP7_75t_SL g2324 ( 
.A(n_2019),
.Y(n_2324)
);

AND2x6_ASAP7_75t_L g2325 ( 
.A(n_2228),
.B(n_1983),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_2136),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2185),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2045),
.B(n_1531),
.Y(n_2328)
);

INVxp67_ASAP7_75t_L g2329 ( 
.A(n_2114),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_2191),
.Y(n_2330)
);

OR2x2_ASAP7_75t_SL g2331 ( 
.A(n_2132),
.B(n_1755),
.Y(n_2331)
);

INVx2_ASAP7_75t_SL g2332 ( 
.A(n_2123),
.Y(n_2332)
);

AO22x2_ASAP7_75t_L g2333 ( 
.A1(n_2229),
.A2(n_1975),
.B1(n_1977),
.B2(n_1974),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2191),
.Y(n_2334)
);

BUFx2_ASAP7_75t_L g2335 ( 
.A(n_2186),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2070),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2222),
.B(n_1978),
.Y(n_2337)
);

INVx3_ASAP7_75t_L g2338 ( 
.A(n_2104),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2060),
.Y(n_2339)
);

AND2x4_ASAP7_75t_L g2340 ( 
.A(n_2112),
.B(n_1531),
.Y(n_2340)
);

OR2x6_ASAP7_75t_L g2341 ( 
.A(n_2058),
.B(n_1870),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2046),
.B(n_2009),
.Y(n_2342)
);

INVxp67_ASAP7_75t_L g2343 ( 
.A(n_2144),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2070),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_2136),
.Y(n_2345)
);

BUFx6f_ASAP7_75t_L g2346 ( 
.A(n_2014),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2062),
.Y(n_2347)
);

NOR2xp33_ASAP7_75t_L g2348 ( 
.A(n_2287),
.B(n_1853),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2073),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2072),
.Y(n_2350)
);

INVx2_ASAP7_75t_L g2351 ( 
.A(n_2072),
.Y(n_2351)
);

NAND3x1_ASAP7_75t_L g2352 ( 
.A(n_2169),
.B(n_2061),
.C(n_2053),
.Y(n_2352)
);

BUFx6f_ASAP7_75t_L g2353 ( 
.A(n_2014),
.Y(n_2353)
);

AND2x2_ASAP7_75t_L g2354 ( 
.A(n_2254),
.B(n_1754),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2074),
.Y(n_2355)
);

NAND3x1_ASAP7_75t_L g2356 ( 
.A(n_2081),
.B(n_1960),
.C(n_1825),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2117),
.B(n_1833),
.Y(n_2357)
);

AND3x4_ASAP7_75t_L g2358 ( 
.A(n_2285),
.B(n_1825),
.C(n_1831),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_2126),
.B(n_2184),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2112),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2022),
.B(n_1767),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_2104),
.Y(n_2362)
);

BUFx6f_ASAP7_75t_L g2363 ( 
.A(n_2014),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2077),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2074),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2087),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_2152),
.B(n_1531),
.Y(n_2367)
);

BUFx6f_ASAP7_75t_L g2368 ( 
.A(n_2048),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2092),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2090),
.Y(n_2370)
);

BUFx3_ASAP7_75t_L g2371 ( 
.A(n_2267),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2254),
.B(n_1762),
.Y(n_2372)
);

INVx4_ASAP7_75t_L g2373 ( 
.A(n_2126),
.Y(n_2373)
);

BUFx3_ASAP7_75t_L g2374 ( 
.A(n_2267),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2094),
.Y(n_2375)
);

AND2x6_ASAP7_75t_L g2376 ( 
.A(n_2228),
.B(n_1622),
.Y(n_2376)
);

BUFx2_ASAP7_75t_L g2377 ( 
.A(n_2016),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2141),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2141),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2117),
.B(n_1847),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2048),
.Y(n_2381)
);

CKINVDCx5p33_ASAP7_75t_R g2382 ( 
.A(n_2021),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2142),
.Y(n_2383)
);

INVx4_ASAP7_75t_L g2384 ( 
.A(n_2126),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2019),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2023),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2075),
.B(n_1767),
.Y(n_2387)
);

INVx4_ASAP7_75t_L g2388 ( 
.A(n_2048),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_2142),
.Y(n_2389)
);

AOI22xp5_ASAP7_75t_L g2390 ( 
.A1(n_2280),
.A2(n_2218),
.B1(n_2184),
.B2(n_2187),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2117),
.B(n_1849),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2090),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2234),
.B(n_1851),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2023),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2203),
.B(n_1746),
.Y(n_2395)
);

INVx1_ASAP7_75t_SL g2396 ( 
.A(n_2233),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_SL g2397 ( 
.A(n_2119),
.B(n_1886),
.Y(n_2397)
);

INVxp67_ASAP7_75t_L g2398 ( 
.A(n_2219),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2095),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2024),
.Y(n_2400)
);

AND2x6_ASAP7_75t_L g2401 ( 
.A(n_2228),
.B(n_1622),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2288),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2024),
.Y(n_2403)
);

INVx4_ASAP7_75t_L g2404 ( 
.A(n_2048),
.Y(n_2404)
);

INVx3_ASAP7_75t_L g2405 ( 
.A(n_2044),
.Y(n_2405)
);

INVx2_ASAP7_75t_SL g2406 ( 
.A(n_2288),
.Y(n_2406)
);

INVxp67_ASAP7_75t_L g2407 ( 
.A(n_2225),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2044),
.Y(n_2408)
);

HB1xp67_ASAP7_75t_L g2409 ( 
.A(n_2230),
.Y(n_2409)
);

BUFx3_ASAP7_75t_L g2410 ( 
.A(n_2267),
.Y(n_2410)
);

NOR2xp33_ASAP7_75t_L g2411 ( 
.A(n_2234),
.B(n_1991),
.Y(n_2411)
);

AND2x2_ASAP7_75t_SL g2412 ( 
.A(n_2119),
.B(n_1625),
.Y(n_2412)
);

INVx1_ASAP7_75t_SL g2413 ( 
.A(n_2150),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_L g2414 ( 
.A(n_2234),
.B(n_1806),
.Y(n_2414)
);

OAI22xp5_ASAP7_75t_SL g2415 ( 
.A1(n_2215),
.A2(n_1925),
.B1(n_1968),
.B2(n_1885),
.Y(n_2415)
);

NAND2xp5_ASAP7_75t_L g2416 ( 
.A(n_2166),
.B(n_1746),
.Y(n_2416)
);

AO22x2_ASAP7_75t_L g2417 ( 
.A1(n_2249),
.A2(n_1762),
.B1(n_1740),
.B2(n_1735),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2025),
.Y(n_2418)
);

AO22x2_ASAP7_75t_L g2419 ( 
.A1(n_2249),
.A2(n_1740),
.B1(n_1735),
.B2(n_1993),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2025),
.Y(n_2420)
);

AOI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2235),
.A2(n_1808),
.B1(n_1574),
.B2(n_1576),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2026),
.Y(n_2422)
);

AND2x4_ASAP7_75t_L g2423 ( 
.A(n_2152),
.B(n_1550),
.Y(n_2423)
);

AND2x4_ASAP7_75t_L g2424 ( 
.A(n_2152),
.B(n_1550),
.Y(n_2424)
);

NAND3xp33_ASAP7_75t_SL g2425 ( 
.A(n_2156),
.B(n_2269),
.C(n_2289),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2262),
.B(n_1967),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2026),
.Y(n_2427)
);

INVx4_ASAP7_75t_L g2428 ( 
.A(n_2007),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2095),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2099),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2089),
.Y(n_2431)
);

AO22x2_ASAP7_75t_L g2432 ( 
.A1(n_2260),
.A2(n_2001),
.B1(n_1961),
.B2(n_1970),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2027),
.Y(n_2433)
);

OR2x6_ASAP7_75t_SL g2434 ( 
.A(n_2008),
.B(n_1566),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_2099),
.Y(n_2435)
);

OAI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2020),
.A2(n_2032),
.B1(n_2035),
.B2(n_2054),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2089),
.Y(n_2437)
);

INVxp33_ASAP7_75t_L g2438 ( 
.A(n_2110),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_2172),
.B(n_1550),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2149),
.Y(n_2440)
);

NAND2x1p5_ASAP7_75t_L g2441 ( 
.A(n_2190),
.B(n_1494),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2155),
.B(n_1557),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2172),
.B(n_2201),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2089),
.Y(n_2444)
);

NOR2xp33_ASAP7_75t_L g2445 ( 
.A(n_2262),
.B(n_1868),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2255),
.B(n_2275),
.Y(n_2446)
);

NOR2xp33_ASAP7_75t_L g2447 ( 
.A(n_2230),
.B(n_1918),
.Y(n_2447)
);

INVx2_ASAP7_75t_SL g2448 ( 
.A(n_2181),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2201),
.B(n_1557),
.Y(n_2449)
);

AOI22xp33_ASAP7_75t_L g2450 ( 
.A1(n_2232),
.A2(n_1987),
.B1(n_1581),
.B2(n_1557),
.Y(n_2450)
);

BUFx3_ASAP7_75t_L g2451 ( 
.A(n_2267),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_2044),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2027),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2039),
.B(n_1581),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2093),
.B(n_1581),
.Y(n_2455)
);

INVxp67_ASAP7_75t_SL g2456 ( 
.A(n_2029),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2029),
.Y(n_2457)
);

INVx4_ASAP7_75t_L g2458 ( 
.A(n_2007),
.Y(n_2458)
);

INVx2_ASAP7_75t_L g2459 ( 
.A(n_2102),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2030),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2231),
.B(n_2086),
.Y(n_2461)
);

AND2x4_ASAP7_75t_L g2462 ( 
.A(n_2155),
.B(n_1951),
.Y(n_2462)
);

NAND2x1p5_ASAP7_75t_L g2463 ( 
.A(n_2190),
.B(n_1494),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_2089),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2086),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2093),
.B(n_1932),
.Y(n_2466)
);

BUFx2_ASAP7_75t_L g2467 ( 
.A(n_2285),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2030),
.Y(n_2468)
);

INVx4_ASAP7_75t_L g2469 ( 
.A(n_2007),
.Y(n_2469)
);

BUFx2_ASAP7_75t_L g2470 ( 
.A(n_2211),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2047),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2102),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2278),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2120),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2096),
.B(n_1566),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2281),
.B(n_1952),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_2089),
.Y(n_2477)
);

NOR2xp33_ASAP7_75t_L g2478 ( 
.A(n_2231),
.B(n_2274),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2047),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2084),
.Y(n_2480)
);

AND2x4_ASAP7_75t_L g2481 ( 
.A(n_2155),
.B(n_1574),
.Y(n_2481)
);

NOR2xp33_ASAP7_75t_L g2482 ( 
.A(n_2274),
.B(n_1895),
.Y(n_2482)
);

AOI22xp5_ASAP7_75t_SL g2483 ( 
.A1(n_2215),
.A2(n_2038),
.B1(n_2253),
.B2(n_2107),
.Y(n_2483)
);

AOI22xp33_ASAP7_75t_SL g2484 ( 
.A1(n_2253),
.A2(n_28),
.B1(n_21),
.B2(n_27),
.Y(n_2484)
);

NOR2xp33_ASAP7_75t_L g2485 ( 
.A(n_2277),
.B(n_1576),
.Y(n_2485)
);

CKINVDCx11_ASAP7_75t_R g2486 ( 
.A(n_2278),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2149),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2154),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2281),
.B(n_1660),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2096),
.B(n_1579),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2108),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2115),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2154),
.Y(n_2493)
);

AND2x4_ASAP7_75t_L g2494 ( 
.A(n_2159),
.B(n_1579),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2129),
.Y(n_2495)
);

AND2x4_ASAP7_75t_L g2496 ( 
.A(n_2159),
.B(n_1583),
.Y(n_2496)
);

AOI22xp33_ASAP7_75t_L g2497 ( 
.A1(n_2232),
.A2(n_1643),
.B1(n_1651),
.B2(n_1640),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2159),
.B(n_1583),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2135),
.Y(n_2499)
);

INVx4_ASAP7_75t_L g2500 ( 
.A(n_2007),
.Y(n_2500)
);

AO22x2_ASAP7_75t_L g2501 ( 
.A1(n_2260),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2120),
.Y(n_2502)
);

AND2x4_ASAP7_75t_L g2503 ( 
.A(n_2145),
.B(n_1588),
.Y(n_2503)
);

INVx1_ASAP7_75t_SL g2504 ( 
.A(n_2173),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2140),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2106),
.B(n_2286),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2071),
.Y(n_2507)
);

AND2x4_ASAP7_75t_L g2508 ( 
.A(n_2145),
.B(n_1588),
.Y(n_2508)
);

INVx3_ASAP7_75t_L g2509 ( 
.A(n_2071),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2124),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2124),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2127),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2127),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2128),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2128),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2071),
.Y(n_2516)
);

AND2x6_ASAP7_75t_L g2517 ( 
.A(n_2268),
.B(n_1625),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2211),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2131),
.Y(n_2519)
);

BUFx6f_ASAP7_75t_L g2520 ( 
.A(n_2148),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2131),
.Y(n_2521)
);

AND2x6_ASAP7_75t_L g2522 ( 
.A(n_2268),
.B(n_2111),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2133),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2133),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2036),
.Y(n_2525)
);

OAI22xp33_ASAP7_75t_L g2526 ( 
.A1(n_2390),
.A2(n_2237),
.B1(n_2245),
.B2(n_2241),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_SL g2527 ( 
.A(n_2307),
.B(n_2145),
.Y(n_2527)
);

OAI21xp5_ASAP7_75t_L g2528 ( 
.A1(n_2342),
.A2(n_2032),
.B(n_2020),
.Y(n_2528)
);

NOR2xp33_ASAP7_75t_L g2529 ( 
.A(n_2348),
.B(n_2253),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2467),
.Y(n_2530)
);

BUFx3_ASAP7_75t_L g2531 ( 
.A(n_2326),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2342),
.B(n_2237),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_SL g2533 ( 
.A(n_2318),
.B(n_2145),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2480),
.B(n_2241),
.Y(n_2534)
);

INVx8_ASAP7_75t_L g2535 ( 
.A(n_2517),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2317),
.B(n_2245),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_2312),
.B(n_2248),
.Y(n_2537)
);

OR2x6_ASAP7_75t_L g2538 ( 
.A(n_2373),
.B(n_2058),
.Y(n_2538)
);

INVx4_ASAP7_75t_L g2539 ( 
.A(n_2373),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2312),
.B(n_2250),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_2343),
.B(n_2251),
.Y(n_2541)
);

NOR2xp33_ASAP7_75t_L g2542 ( 
.A(n_2348),
.B(n_2210),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2343),
.B(n_2264),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2306),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2291),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_SL g2546 ( 
.A(n_2318),
.B(n_2190),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2489),
.B(n_2272),
.Y(n_2547)
);

AOI22xp33_ASAP7_75t_L g2548 ( 
.A1(n_2501),
.A2(n_2271),
.B1(n_2209),
.B2(n_2206),
.Y(n_2548)
);

NAND2x1_ASAP7_75t_L g2549 ( 
.A(n_2405),
.B(n_2148),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2387),
.B(n_2279),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2308),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2510),
.Y(n_2552)
);

AND2x4_ASAP7_75t_L g2553 ( 
.A(n_2473),
.B(n_2063),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_2332),
.B(n_2190),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2506),
.B(n_2111),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2324),
.B(n_2282),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2291),
.Y(n_2557)
);

AOI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2501),
.A2(n_2289),
.B1(n_2170),
.B2(n_2183),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2511),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2512),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2324),
.B(n_2261),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_SL g2562 ( 
.A(n_2337),
.B(n_2190),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2329),
.B(n_2204),
.Y(n_2563)
);

INVxp33_ASAP7_75t_L g2564 ( 
.A(n_2315),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2456),
.B(n_2263),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2514),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2456),
.B(n_2134),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2361),
.B(n_2066),
.Y(n_2568)
);

O2A1O1Ixp33_ASAP7_75t_L g2569 ( 
.A1(n_2395),
.A2(n_2196),
.B(n_2153),
.C(n_2200),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_L g2570 ( 
.A(n_2413),
.B(n_2210),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2445),
.B(n_2208),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2515),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2519),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2445),
.B(n_2224),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_2447),
.B(n_2443),
.Y(n_2575)
);

INVx4_ASAP7_75t_L g2576 ( 
.A(n_2384),
.Y(n_2576)
);

OAI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2412),
.A2(n_2207),
.B1(n_2204),
.B2(n_2065),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2524),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2447),
.B(n_2439),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_2329),
.B(n_2210),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_2446),
.B(n_2277),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2449),
.B(n_2224),
.Y(n_2582)
);

NOR2xp33_ASAP7_75t_L g2583 ( 
.A(n_2446),
.B(n_2175),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2339),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2347),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2292),
.B(n_2204),
.Y(n_2586)
);

INVx3_ASAP7_75t_L g2587 ( 
.A(n_2520),
.Y(n_2587)
);

BUFx5_ASAP7_75t_L g2588 ( 
.A(n_2522),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_L g2589 ( 
.A(n_2299),
.B(n_2224),
.Y(n_2589)
);

AOI22xp33_ASAP7_75t_L g2590 ( 
.A1(n_2501),
.A2(n_2158),
.B1(n_2202),
.B2(n_2268),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2476),
.B(n_2240),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_2412),
.B(n_2204),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2349),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2426),
.A2(n_2180),
.B1(n_2244),
.B2(n_2063),
.Y(n_2594)
);

INVx2_ASAP7_75t_SL g2595 ( 
.A(n_2326),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2364),
.Y(n_2596)
);

OAI21xp33_ASAP7_75t_L g2597 ( 
.A1(n_2426),
.A2(n_2256),
.B(n_2217),
.Y(n_2597)
);

AOI22xp33_ASAP7_75t_L g2598 ( 
.A1(n_2436),
.A2(n_2242),
.B1(n_2035),
.B2(n_2153),
.Y(n_2598)
);

A2O1A1Ixp33_ASAP7_75t_L g2599 ( 
.A1(n_2425),
.A2(n_2196),
.B(n_2221),
.C(n_2193),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_2448),
.B(n_2204),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2482),
.B(n_2213),
.Y(n_2601)
);

INVx3_ASAP7_75t_L g2602 ( 
.A(n_2520),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2482),
.B(n_2180),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_SL g2604 ( 
.A(n_2461),
.B(n_2207),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2461),
.B(n_2411),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_L g2606 ( 
.A1(n_2359),
.A2(n_2207),
.B1(n_2088),
.B2(n_2083),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2297),
.Y(n_2607)
);

AND2x2_ASAP7_75t_L g2608 ( 
.A(n_2372),
.B(n_2063),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2297),
.Y(n_2609)
);

NOR2xp33_ASAP7_75t_L g2610 ( 
.A(n_2411),
.B(n_2146),
.Y(n_2610)
);

NAND2x1p5_ASAP7_75t_L g2611 ( 
.A(n_2384),
.B(n_2207),
.Y(n_2611)
);

NOR2xp67_ASAP7_75t_L g2612 ( 
.A(n_2321),
.B(n_2259),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2454),
.B(n_2205),
.Y(n_2613)
);

OAI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2359),
.A2(n_2207),
.B1(n_2434),
.B2(n_2416),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_R g2615 ( 
.A(n_2382),
.B(n_2278),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_SL g2616 ( 
.A(n_2295),
.B(n_2259),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2366),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_2345),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2354),
.B(n_2151),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_L g2620 ( 
.A(n_2465),
.B(n_2211),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_SL g2621 ( 
.A(n_2302),
.B(n_2038),
.Y(n_2621)
);

OAI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2322),
.A2(n_2284),
.B1(n_2193),
.B2(n_2130),
.Y(n_2622)
);

INVx2_ASAP7_75t_SL g2623 ( 
.A(n_2345),
.Y(n_2623)
);

NOR2xp33_ASAP7_75t_L g2624 ( 
.A(n_2327),
.B(n_2211),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2520),
.Y(n_2625)
);

AOI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2380),
.A2(n_2078),
.B1(n_2151),
.B2(n_2239),
.Y(n_2626)
);

AOI22xp5_ASAP7_75t_L g2627 ( 
.A1(n_2380),
.A2(n_2078),
.B1(n_2151),
.B2(n_2239),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2369),
.B(n_2058),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2375),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_SL g2630 ( 
.A(n_2302),
.B(n_2078),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2316),
.B(n_2162),
.Y(n_2631)
);

NOR2xp67_ASAP7_75t_L g2632 ( 
.A(n_2425),
.B(n_2259),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2305),
.Y(n_2633)
);

BUFx6f_ASAP7_75t_L g2634 ( 
.A(n_2520),
.Y(n_2634)
);

NOR2xp33_ASAP7_75t_L g2635 ( 
.A(n_2327),
.B(n_2162),
.Y(n_2635)
);

AND3x1_ASAP7_75t_L g2636 ( 
.A(n_2414),
.B(n_2236),
.C(n_2238),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2305),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_2316),
.B(n_2162),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_SL g2639 ( 
.A(n_2328),
.B(n_2162),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_L g2640 ( 
.A(n_2478),
.B(n_2058),
.Y(n_2640)
);

AND2x2_ASAP7_75t_L g2641 ( 
.A(n_2438),
.B(n_2164),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2303),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2319),
.Y(n_2643)
);

NAND2xp5_ASAP7_75t_L g2644 ( 
.A(n_2478),
.B(n_2239),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2328),
.B(n_2164),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2409),
.B(n_2239),
.Y(n_2646)
);

NOR2xp67_ASAP7_75t_L g2647 ( 
.A(n_2402),
.B(n_2259),
.Y(n_2647)
);

AND2x6_ASAP7_75t_SL g2648 ( 
.A(n_2341),
.B(n_2247),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2409),
.B(n_2398),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2398),
.B(n_2239),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2377),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2438),
.B(n_2164),
.Y(n_2652)
);

AND3x1_ASAP7_75t_L g2653 ( 
.A(n_2414),
.B(n_2138),
.C(n_2031),
.Y(n_2653)
);

CKINVDCx20_ASAP7_75t_R g2654 ( 
.A(n_2295),
.Y(n_2654)
);

CKINVDCx5p33_ASAP7_75t_R g2655 ( 
.A(n_2298),
.Y(n_2655)
);

INVx2_ASAP7_75t_SL g2656 ( 
.A(n_2335),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2319),
.Y(n_2657)
);

NAND2x1_ASAP7_75t_L g2658 ( 
.A(n_2405),
.B(n_2148),
.Y(n_2658)
);

AND2x6_ASAP7_75t_L g2659 ( 
.A(n_2408),
.B(n_2082),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2304),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_2313),
.B(n_2164),
.Y(n_2661)
);

NAND3xp33_ASAP7_75t_L g2662 ( 
.A(n_2391),
.B(n_2200),
.C(n_2273),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2407),
.B(n_2239),
.Y(n_2663)
);

OR2x6_ASAP7_75t_L g2664 ( 
.A(n_2428),
.B(n_2189),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2431),
.Y(n_2665)
);

INVx2_ASAP7_75t_L g2666 ( 
.A(n_2320),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_L g2667 ( 
.A1(n_2484),
.A2(n_2270),
.B1(n_2283),
.B2(n_2214),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2407),
.B(n_2270),
.Y(n_2668)
);

INVx2_ASAP7_75t_L g2669 ( 
.A(n_2320),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_L g2670 ( 
.A(n_2396),
.B(n_2189),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_SL g2671 ( 
.A1(n_2393),
.A2(n_2223),
.B1(n_2252),
.B2(n_2173),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2340),
.B(n_2367),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2340),
.B(n_2028),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2485),
.B(n_2491),
.Y(n_2674)
);

NOR2xp33_ASAP7_75t_L g2675 ( 
.A(n_2393),
.B(n_2189),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2323),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2360),
.B(n_2273),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2485),
.B(n_2492),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2323),
.Y(n_2679)
);

NAND2xp5_ASAP7_75t_L g2680 ( 
.A(n_2495),
.B(n_2283),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2336),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2367),
.B(n_2028),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2462),
.B(n_2033),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_2484),
.A2(n_2214),
.B1(n_2266),
.B2(n_2227),
.Y(n_2684)
);

NOR2xp33_ASAP7_75t_L g2685 ( 
.A(n_2391),
.B(n_2189),
.Y(n_2685)
);

INVx2_ASAP7_75t_SL g2686 ( 
.A(n_2504),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2336),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2344),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2499),
.B(n_2082),
.Y(n_2689)
);

NOR2xp33_ASAP7_75t_L g2690 ( 
.A(n_2357),
.B(n_2031),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2505),
.B(n_2212),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2344),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2350),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2350),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_SL g2695 ( 
.A(n_2423),
.B(n_2259),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_SL g2696 ( 
.A1(n_2483),
.A2(n_2284),
.B1(n_2017),
.B2(n_2121),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_SL g2697 ( 
.A(n_2423),
.B(n_2284),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2351),
.Y(n_2698)
);

OR2x6_ASAP7_75t_L g2699 ( 
.A(n_2428),
.B(n_2278),
.Y(n_2699)
);

OR2x2_ASAP7_75t_L g2700 ( 
.A(n_2406),
.B(n_2266),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_2294),
.A2(n_2214),
.B1(n_2227),
.B2(n_2226),
.Y(n_2701)
);

NOR2xp33_ASAP7_75t_SL g2702 ( 
.A(n_2298),
.B(n_2223),
.Y(n_2702)
);

AOI22xp5_ASAP7_75t_L g2703 ( 
.A1(n_2357),
.A2(n_2265),
.B1(n_2118),
.B2(n_2122),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2330),
.B(n_2037),
.Y(n_2704)
);

NOR2xp33_ASAP7_75t_L g2705 ( 
.A(n_2334),
.B(n_2040),
.Y(n_2705)
);

AND2x6_ASAP7_75t_SL g2706 ( 
.A(n_2341),
.B(n_2192),
.Y(n_2706)
);

NOR3xp33_ASAP7_75t_L g2707 ( 
.A(n_2397),
.B(n_2265),
.C(n_2122),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_SL g2708 ( 
.A(n_2424),
.B(n_2284),
.Y(n_2708)
);

BUFx3_ASAP7_75t_L g2709 ( 
.A(n_2371),
.Y(n_2709)
);

INVx3_ASAP7_75t_L g2710 ( 
.A(n_2431),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2466),
.B(n_2226),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2351),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2293),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2537),
.B(n_2540),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_L g2715 ( 
.A(n_2601),
.B(n_2522),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2584),
.Y(n_2716)
);

OR2x6_ASAP7_75t_L g2717 ( 
.A(n_2535),
.B(n_2458),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_L g2718 ( 
.A(n_2575),
.B(n_2522),
.Y(n_2718)
);

INVx2_ASAP7_75t_SL g2719 ( 
.A(n_2531),
.Y(n_2719)
);

CKINVDCx5p33_ASAP7_75t_R g2720 ( 
.A(n_2655),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2585),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2571),
.B(n_2421),
.Y(n_2722)
);

INVx5_ASAP7_75t_L g2723 ( 
.A(n_2659),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2654),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2593),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2596),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2535),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2579),
.B(n_2522),
.Y(n_2728)
);

NOR2x2_ASAP7_75t_L g2729 ( 
.A(n_2664),
.B(n_2341),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2608),
.B(n_2419),
.Y(n_2730)
);

AOI22xp5_ASAP7_75t_L g2731 ( 
.A1(n_2529),
.A2(n_2352),
.B1(n_2356),
.B2(n_2462),
.Y(n_2731)
);

AND2x4_ASAP7_75t_L g2732 ( 
.A(n_2553),
.B(n_2473),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2545),
.Y(n_2733)
);

INVx6_ASAP7_75t_L g2734 ( 
.A(n_2699),
.Y(n_2734)
);

INVxp67_ASAP7_75t_L g2735 ( 
.A(n_2651),
.Y(n_2735)
);

INVx1_ASAP7_75t_SL g2736 ( 
.A(n_2651),
.Y(n_2736)
);

INVxp67_ASAP7_75t_SL g2737 ( 
.A(n_2567),
.Y(n_2737)
);

NAND2xp5_ASAP7_75t_L g2738 ( 
.A(n_2568),
.B(n_2522),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2617),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2550),
.B(n_2385),
.Y(n_2740)
);

INVxp67_ASAP7_75t_SL g2741 ( 
.A(n_2556),
.Y(n_2741)
);

INVx2_ASAP7_75t_L g2742 ( 
.A(n_2557),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2607),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2629),
.Y(n_2744)
);

CKINVDCx8_ASAP7_75t_R g2745 ( 
.A(n_2648),
.Y(n_2745)
);

INVx2_ASAP7_75t_SL g2746 ( 
.A(n_2595),
.Y(n_2746)
);

NAND2x1p5_ASAP7_75t_L g2747 ( 
.A(n_2697),
.B(n_2458),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2605),
.B(n_2147),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2605),
.B(n_2397),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2544),
.Y(n_2750)
);

CKINVDCx5p33_ASAP7_75t_R g2751 ( 
.A(n_2615),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2551),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2552),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2559),
.Y(n_2754)
);

INVx3_ASAP7_75t_L g2755 ( 
.A(n_2535),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2560),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2610),
.B(n_2386),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2609),
.Y(n_2758)
);

NOR2xp33_ASAP7_75t_L g2759 ( 
.A(n_2564),
.B(n_2415),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2566),
.Y(n_2760)
);

HB1xp67_ASAP7_75t_L g2761 ( 
.A(n_2677),
.Y(n_2761)
);

INVx2_ASAP7_75t_SL g2762 ( 
.A(n_2618),
.Y(n_2762)
);

BUFx6f_ASAP7_75t_L g2763 ( 
.A(n_2709),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2572),
.Y(n_2764)
);

INVx3_ASAP7_75t_L g2765 ( 
.A(n_2634),
.Y(n_2765)
);

AOI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2529),
.A2(n_2358),
.B1(n_2442),
.B2(n_2424),
.Y(n_2766)
);

NAND2xp5_ASAP7_75t_L g2767 ( 
.A(n_2610),
.B(n_2394),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2573),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2666),
.Y(n_2769)
);

INVx2_ASAP7_75t_SL g2770 ( 
.A(n_2623),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2578),
.Y(n_2771)
);

BUFx3_ASAP7_75t_L g2772 ( 
.A(n_2656),
.Y(n_2772)
);

HB1xp67_ASAP7_75t_L g2773 ( 
.A(n_2649),
.Y(n_2773)
);

AND2x6_ASAP7_75t_L g2774 ( 
.A(n_2626),
.B(n_2408),
.Y(n_2774)
);

OR2x2_ASAP7_75t_SL g2775 ( 
.A(n_2591),
.B(n_2331),
.Y(n_2775)
);

BUFx6f_ASAP7_75t_L g2776 ( 
.A(n_2713),
.Y(n_2776)
);

INVx5_ASAP7_75t_L g2777 ( 
.A(n_2659),
.Y(n_2777)
);

BUFx6f_ASAP7_75t_L g2778 ( 
.A(n_2713),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2669),
.Y(n_2779)
);

BUFx3_ASAP7_75t_L g2780 ( 
.A(n_2686),
.Y(n_2780)
);

INVx2_ASAP7_75t_SL g2781 ( 
.A(n_2641),
.Y(n_2781)
);

INVx3_ASAP7_75t_L g2782 ( 
.A(n_2634),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2553),
.B(n_2371),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2667),
.A2(n_2358),
.B1(n_2294),
.B2(n_2333),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_SL g2785 ( 
.A(n_2542),
.B(n_2109),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2642),
.Y(n_2786)
);

INVx4_ASAP7_75t_L g2787 ( 
.A(n_2634),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2660),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2542),
.B(n_2603),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2679),
.Y(n_2790)
);

AND3x1_ASAP7_75t_SL g2791 ( 
.A(n_2530),
.B(n_2417),
.C(n_2333),
.Y(n_2791)
);

INVx1_ASAP7_75t_SL g2792 ( 
.A(n_2652),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2633),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_SL g2794 ( 
.A(n_2594),
.B(n_2574),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2681),
.Y(n_2795)
);

CKINVDCx5p33_ASAP7_75t_R g2796 ( 
.A(n_2570),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_2664),
.B(n_2374),
.Y(n_2797)
);

INVx3_ASAP7_75t_L g2798 ( 
.A(n_2634),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2637),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_SL g2800 ( 
.A(n_2653),
.B(n_2597),
.Y(n_2800)
);

BUFx12f_ASAP7_75t_L g2801 ( 
.A(n_2538),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2683),
.B(n_2419),
.Y(n_2802)
);

INVx2_ASAP7_75t_SL g2803 ( 
.A(n_2589),
.Y(n_2803)
);

INVx2_ASAP7_75t_SL g2804 ( 
.A(n_2620),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2636),
.A2(n_2442),
.B1(n_2494),
.B2(n_2481),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2687),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2532),
.B(n_2400),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2688),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2643),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2711),
.B(n_2403),
.Y(n_2810)
);

INVx2_ASAP7_75t_SL g2811 ( 
.A(n_2670),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2561),
.B(n_2418),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2692),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2657),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2676),
.Y(n_2815)
);

BUFx12f_ASAP7_75t_L g2816 ( 
.A(n_2538),
.Y(n_2816)
);

AND2x4_ASAP7_75t_L g2817 ( 
.A(n_2664),
.B(n_2374),
.Y(n_2817)
);

INVx1_ASAP7_75t_SL g2818 ( 
.A(n_2702),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2693),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_L g2820 ( 
.A1(n_2667),
.A2(n_2294),
.B1(n_2333),
.B2(n_2417),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2712),
.Y(n_2821)
);

CKINVDCx5p33_ASAP7_75t_R g2822 ( 
.A(n_2580),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2565),
.B(n_2420),
.Y(n_2823)
);

INVx3_ASAP7_75t_L g2824 ( 
.A(n_2539),
.Y(n_2824)
);

INVx4_ASAP7_75t_L g2825 ( 
.A(n_2538),
.Y(n_2825)
);

BUFx3_ASAP7_75t_L g2826 ( 
.A(n_2624),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2694),
.Y(n_2827)
);

INVx2_ASAP7_75t_SL g2828 ( 
.A(n_2671),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2698),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2700),
.Y(n_2830)
);

AND2x6_ASAP7_75t_L g2831 ( 
.A(n_2627),
.B(n_2452),
.Y(n_2831)
);

INVx4_ASAP7_75t_L g2832 ( 
.A(n_2713),
.Y(n_2832)
);

NAND2xp5_ASAP7_75t_L g2833 ( 
.A(n_2613),
.B(n_2422),
.Y(n_2833)
);

HB1xp67_ASAP7_75t_L g2834 ( 
.A(n_2635),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2624),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2526),
.B(n_2427),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2526),
.B(n_2598),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_2580),
.Y(n_2838)
);

BUFx2_ASAP7_75t_L g2839 ( 
.A(n_2665),
.Y(n_2839)
);

OR2x6_ASAP7_75t_L g2840 ( 
.A(n_2699),
.B(n_2469),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2598),
.B(n_2433),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2619),
.B(n_2419),
.Y(n_2842)
);

OR2x6_ASAP7_75t_L g2843 ( 
.A(n_2699),
.B(n_2708),
.Y(n_2843)
);

BUFx3_ASAP7_75t_L g2844 ( 
.A(n_2665),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2547),
.B(n_2525),
.Y(n_2845)
);

INVx1_ASAP7_75t_SL g2846 ( 
.A(n_2583),
.Y(n_2846)
);

AND2x4_ASAP7_75t_L g2847 ( 
.A(n_2672),
.B(n_2410),
.Y(n_2847)
);

OR2x4_ASAP7_75t_L g2848 ( 
.A(n_2583),
.B(n_2368),
.Y(n_2848)
);

CKINVDCx5p33_ASAP7_75t_R g2849 ( 
.A(n_2706),
.Y(n_2849)
);

AND2x6_ASAP7_75t_L g2850 ( 
.A(n_2703),
.B(n_2452),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2536),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2680),
.Y(n_2852)
);

AOI22xp33_ASAP7_75t_L g2853 ( 
.A1(n_2621),
.A2(n_2417),
.B1(n_2432),
.B2(n_2325),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2668),
.Y(n_2854)
);

INVx3_ASAP7_75t_L g2855 ( 
.A(n_2539),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2534),
.Y(n_2856)
);

INVx2_ASAP7_75t_L g2857 ( 
.A(n_2691),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2555),
.B(n_2453),
.Y(n_2858)
);

AND2x4_ASAP7_75t_L g2859 ( 
.A(n_2630),
.B(n_2410),
.Y(n_2859)
);

INVx2_ASAP7_75t_SL g2860 ( 
.A(n_2710),
.Y(n_2860)
);

AO22x1_ASAP7_75t_L g2861 ( 
.A1(n_2675),
.A2(n_2481),
.B1(n_2496),
.B2(n_2494),
.Y(n_2861)
);

AND2x2_ASAP7_75t_L g2862 ( 
.A(n_2581),
.B(n_2432),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_SL g2863 ( 
.A(n_2696),
.B(n_2528),
.Y(n_2863)
);

INVx5_ASAP7_75t_L g2864 ( 
.A(n_2659),
.Y(n_2864)
);

NOR2xp33_ASAP7_75t_L g2865 ( 
.A(n_2533),
.B(n_2470),
.Y(n_2865)
);

HB1xp67_ASAP7_75t_L g2866 ( 
.A(n_2635),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_2710),
.Y(n_2867)
);

INVx3_ASAP7_75t_SL g2868 ( 
.A(n_2586),
.Y(n_2868)
);

NAND2xp5_ASAP7_75t_L g2869 ( 
.A(n_2701),
.B(n_2457),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2541),
.Y(n_2870)
);

INVx1_ASAP7_75t_SL g2871 ( 
.A(n_2640),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_2576),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2543),
.Y(n_2873)
);

HB1xp67_ASAP7_75t_L g2874 ( 
.A(n_2707),
.Y(n_2874)
);

AND2x4_ASAP7_75t_L g2875 ( 
.A(n_2612),
.B(n_2451),
.Y(n_2875)
);

INVx3_ASAP7_75t_L g2876 ( 
.A(n_2576),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2674),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2704),
.Y(n_2878)
);

AOI22xp5_ASAP7_75t_L g2879 ( 
.A1(n_2562),
.A2(n_2498),
.B1(n_2508),
.B2(n_2503),
.Y(n_2879)
);

BUFx3_ASAP7_75t_L g2880 ( 
.A(n_2587),
.Y(n_2880)
);

AND2x6_ASAP7_75t_SL g2881 ( 
.A(n_2685),
.B(n_2498),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2704),
.Y(n_2882)
);

INVx1_ASAP7_75t_SL g2883 ( 
.A(n_2628),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2701),
.B(n_2460),
.Y(n_2884)
);

OAI21xp5_ASAP7_75t_L g2885 ( 
.A1(n_2599),
.A2(n_2662),
.B(n_2569),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2587),
.Y(n_2886)
);

INVx3_ASAP7_75t_L g2887 ( 
.A(n_2611),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2684),
.B(n_2468),
.Y(n_2888)
);

CKINVDCx5p33_ASAP7_75t_R g2889 ( 
.A(n_2690),
.Y(n_2889)
);

HB1xp67_ASAP7_75t_L g2890 ( 
.A(n_2707),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2705),
.Y(n_2891)
);

OR2x4_ASAP7_75t_L g2892 ( 
.A(n_2581),
.B(n_2368),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_2546),
.B(n_2582),
.Y(n_2893)
);

INVx2_ASAP7_75t_SL g2894 ( 
.A(n_2602),
.Y(n_2894)
);

CKINVDCx5p33_ASAP7_75t_R g2895 ( 
.A(n_2713),
.Y(n_2895)
);

INVx5_ASAP7_75t_L g2896 ( 
.A(n_2659),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2611),
.Y(n_2897)
);

INVx4_ASAP7_75t_L g2898 ( 
.A(n_2602),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2705),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2714),
.B(n_2678),
.Y(n_2900)
);

OR2x2_ASAP7_75t_L g2901 ( 
.A(n_2761),
.B(n_2527),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2885),
.A2(n_2105),
.B(n_2606),
.Y(n_2902)
);

AND2x4_ASAP7_75t_L g2903 ( 
.A(n_2825),
.B(n_2563),
.Y(n_2903)
);

AO21x2_ASAP7_75t_L g2904 ( 
.A1(n_2785),
.A2(n_2632),
.B(n_2079),
.Y(n_2904)
);

AOI21xp5_ASAP7_75t_L g2905 ( 
.A1(n_2748),
.A2(n_2105),
.B(n_2577),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2733),
.Y(n_2906)
);

AOI22x1_ASAP7_75t_L g2907 ( 
.A1(n_2889),
.A2(n_2432),
.B1(n_2310),
.B2(n_2296),
.Y(n_2907)
);

NOR2xp67_ASAP7_75t_L g2908 ( 
.A(n_2803),
.B(n_2252),
.Y(n_2908)
);

NAND2xp5_ASAP7_75t_L g2909 ( 
.A(n_2714),
.B(n_2548),
.Y(n_2909)
);

BUFx6f_ASAP7_75t_L g2910 ( 
.A(n_2763),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2761),
.Y(n_2911)
);

NAND2x1p5_ASAP7_75t_L g2912 ( 
.A(n_2723),
.B(n_2604),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2792),
.B(n_2548),
.Y(n_2913)
);

INVx4_ASAP7_75t_L g2914 ( 
.A(n_2763),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2870),
.B(n_2684),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_L g2916 ( 
.A(n_2873),
.B(n_2558),
.Y(n_2916)
);

NOR2xp33_ASAP7_75t_L g2917 ( 
.A(n_2846),
.B(n_2518),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2748),
.A2(n_2785),
.B(n_2722),
.Y(n_2918)
);

OR2x6_ASAP7_75t_L g2919 ( 
.A(n_2843),
.B(n_2569),
.Y(n_2919)
);

INVx6_ASAP7_75t_L g2920 ( 
.A(n_2763),
.Y(n_2920)
);

A2O1A1Ixp33_ASAP7_75t_L g2921 ( 
.A1(n_2731),
.A2(n_2696),
.B(n_2661),
.C(n_2622),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2742),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2722),
.A2(n_2079),
.B(n_2067),
.Y(n_2923)
);

NOR2xp67_ASAP7_75t_L g2924 ( 
.A(n_2796),
.B(n_2682),
.Y(n_2924)
);

NAND3xp33_ASAP7_75t_SL g2925 ( 
.A(n_2745),
.B(n_2616),
.C(n_2600),
.Y(n_2925)
);

AOI22xp33_ASAP7_75t_L g2926 ( 
.A1(n_2749),
.A2(n_2614),
.B1(n_2592),
.B2(n_2503),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2743),
.Y(n_2927)
);

AOI21xp5_ASAP7_75t_L g2928 ( 
.A1(n_2737),
.A2(n_2067),
.B(n_2055),
.Y(n_2928)
);

AOI21xp5_ASAP7_75t_L g2929 ( 
.A1(n_2737),
.A2(n_2055),
.B(n_2121),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2758),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2789),
.B(n_2590),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2741),
.A2(n_2658),
.B(n_2549),
.Y(n_2932)
);

BUFx8_ASAP7_75t_L g2933 ( 
.A(n_2804),
.Y(n_2933)
);

NOR2xp33_ASAP7_75t_L g2934 ( 
.A(n_2789),
.B(n_2673),
.Y(n_2934)
);

NAND2xp5_ASAP7_75t_L g2935 ( 
.A(n_2877),
.B(n_2854),
.Y(n_2935)
);

AND2x2_ASAP7_75t_L g2936 ( 
.A(n_2781),
.B(n_2661),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2811),
.B(n_2588),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2769),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_L g2939 ( 
.A(n_2772),
.Y(n_2939)
);

O2A1O1Ixp33_ASAP7_75t_SL g2940 ( 
.A1(n_2800),
.A2(n_2749),
.B(n_2767),
.C(n_2757),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_L g2941 ( 
.A(n_2871),
.B(n_2590),
.Y(n_2941)
);

A2O1A1Ixp33_ASAP7_75t_L g2942 ( 
.A1(n_2800),
.A2(n_2759),
.B(n_2845),
.C(n_2766),
.Y(n_2942)
);

INVx2_ASAP7_75t_L g2943 ( 
.A(n_2779),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_SL g2944 ( 
.A(n_2822),
.B(n_2588),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2790),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_2838),
.B(n_2588),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_R g2947 ( 
.A(n_2724),
.B(n_2486),
.Y(n_2947)
);

AND2x4_ASAP7_75t_L g2948 ( 
.A(n_2825),
.B(n_2554),
.Y(n_2948)
);

AOI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2794),
.A2(n_2325),
.B1(n_2276),
.B2(n_2650),
.Y(n_2949)
);

O2A1O1Ixp33_ASAP7_75t_L g2950 ( 
.A1(n_2845),
.A2(n_2276),
.B(n_2645),
.C(n_2639),
.Y(n_2950)
);

AOI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2794),
.A2(n_2325),
.B1(n_2663),
.B2(n_2644),
.Y(n_2951)
);

NAND3xp33_ASAP7_75t_L g2952 ( 
.A(n_2893),
.B(n_2837),
.C(n_2863),
.Y(n_2952)
);

O2A1O1Ixp33_ASAP7_75t_L g2953 ( 
.A1(n_2863),
.A2(n_2837),
.B(n_2767),
.C(n_2757),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2802),
.B(n_2631),
.Y(n_2954)
);

BUFx12f_ASAP7_75t_L g2955 ( 
.A(n_2720),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_2741),
.A2(n_2174),
.B(n_2171),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2773),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2833),
.A2(n_2174),
.B(n_2171),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_SL g2959 ( 
.A(n_2805),
.B(n_2883),
.Y(n_2959)
);

AOI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2833),
.A2(n_2179),
.B(n_2178),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2795),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_SL g2962 ( 
.A(n_2828),
.B(n_2588),
.Y(n_2962)
);

AOI21xp33_ASAP7_75t_L g2963 ( 
.A1(n_2893),
.A2(n_2646),
.B(n_2118),
.Y(n_2963)
);

AND2x2_ASAP7_75t_L g2964 ( 
.A(n_2730),
.B(n_2638),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2857),
.B(n_2689),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2738),
.A2(n_2199),
.B(n_2113),
.Y(n_2966)
);

BUFx6f_ASAP7_75t_L g2967 ( 
.A(n_2780),
.Y(n_2967)
);

AOI22xp5_ASAP7_75t_L g2968 ( 
.A1(n_2759),
.A2(n_2325),
.B1(n_2176),
.B2(n_2508),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2852),
.B(n_2471),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2773),
.Y(n_2970)
);

AOI21xp5_ASAP7_75t_L g2971 ( 
.A1(n_2723),
.A2(n_2179),
.B(n_2178),
.Y(n_2971)
);

CKINVDCx5p33_ASAP7_75t_R g2972 ( 
.A(n_2751),
.Y(n_2972)
);

AOI33xp33_ASAP7_75t_L g2973 ( 
.A1(n_2784),
.A2(n_2450),
.A3(n_1890),
.B1(n_2052),
.B2(n_2056),
.B3(n_2050),
.Y(n_2973)
);

OAI21xp5_ASAP7_75t_L g2974 ( 
.A1(n_2740),
.A2(n_2064),
.B(n_2290),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2830),
.B(n_2851),
.Y(n_2975)
);

AOI22xp5_ASAP7_75t_L g2976 ( 
.A1(n_2862),
.A2(n_2325),
.B1(n_2176),
.B2(n_2376),
.Y(n_2976)
);

AOI21xp5_ASAP7_75t_L g2977 ( 
.A1(n_2723),
.A2(n_2148),
.B(n_2290),
.Y(n_2977)
);

AOI21xp5_ASAP7_75t_L g2978 ( 
.A1(n_2723),
.A2(n_2148),
.B(n_2064),
.Y(n_2978)
);

OAI321xp33_ASAP7_75t_L g2979 ( 
.A1(n_2784),
.A2(n_2450),
.A3(n_2695),
.B1(n_2310),
.B2(n_2296),
.C(n_2258),
.Y(n_2979)
);

NAND2xp33_ASAP7_75t_L g2980 ( 
.A(n_2849),
.B(n_2588),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2716),
.Y(n_2981)
);

INVx1_ASAP7_75t_L g2982 ( 
.A(n_2721),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2806),
.Y(n_2983)
);

AOI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2777),
.A2(n_2509),
.B(n_2507),
.Y(n_2984)
);

AOI21xp5_ASAP7_75t_L g2985 ( 
.A1(n_2777),
.A2(n_2509),
.B(n_2507),
.Y(n_2985)
);

NAND2xp5_ASAP7_75t_L g2986 ( 
.A(n_2856),
.B(n_2899),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2808),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2776),
.Y(n_2988)
);

BUFx4f_ASAP7_75t_SL g2989 ( 
.A(n_2801),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2775),
.B(n_2451),
.Y(n_2990)
);

A2O1A1Ixp33_ASAP7_75t_SL g2991 ( 
.A1(n_2865),
.A2(n_2625),
.B(n_2314),
.C(n_2378),
.Y(n_2991)
);

AOI21xp5_ASAP7_75t_L g2992 ( 
.A1(n_2777),
.A2(n_2516),
.B(n_2080),
.Y(n_2992)
);

A2O1A1Ixp33_ASAP7_75t_SL g2993 ( 
.A1(n_2865),
.A2(n_2625),
.B(n_2379),
.C(n_2311),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2725),
.Y(n_2994)
);

CKINVDCx10_ASAP7_75t_R g2995 ( 
.A(n_2717),
.Y(n_2995)
);

OAI22x1_ASAP7_75t_L g2996 ( 
.A1(n_2874),
.A2(n_2500),
.B1(n_2469),
.B2(n_2479),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2834),
.B(n_2383),
.Y(n_2997)
);

BUFx2_ASAP7_75t_L g2998 ( 
.A(n_2826),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2878),
.B(n_2355),
.Y(n_2999)
);

NOR2xp33_ASAP7_75t_L g3000 ( 
.A(n_2818),
.B(n_2486),
.Y(n_3000)
);

INVx2_ASAP7_75t_SL g3001 ( 
.A(n_2719),
.Y(n_3001)
);

NOR2xp33_ASAP7_75t_L g3002 ( 
.A(n_2835),
.B(n_2049),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_L g3003 ( 
.A(n_2882),
.B(n_2355),
.Y(n_3003)
);

OAI22x1_ASAP7_75t_L g3004 ( 
.A1(n_2874),
.A2(n_2500),
.B1(n_2370),
.B2(n_2392),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2891),
.B(n_2365),
.Y(n_3005)
);

BUFx8_ASAP7_75t_SL g3006 ( 
.A(n_2816),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2736),
.B(n_2740),
.Y(n_3007)
);

BUFx2_ASAP7_75t_L g3008 ( 
.A(n_2895),
.Y(n_3008)
);

OAI22xp5_ASAP7_75t_L g3009 ( 
.A1(n_2892),
.A2(n_2647),
.B1(n_2284),
.B2(n_2497),
.Y(n_3009)
);

AOI22xp33_ASAP7_75t_L g3010 ( 
.A1(n_2890),
.A2(n_2850),
.B1(n_2774),
.B2(n_2831),
.Y(n_3010)
);

AOI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2861),
.A2(n_2257),
.B(n_2246),
.Y(n_3011)
);

OA22x2_ASAP7_75t_L g3012 ( 
.A1(n_2879),
.A2(n_2404),
.B1(n_2388),
.B2(n_2389),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2813),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2834),
.B(n_2365),
.Y(n_3014)
);

AOI22xp5_ASAP7_75t_L g3015 ( 
.A1(n_2853),
.A2(n_2376),
.B1(n_2401),
.B2(n_2214),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2866),
.B(n_2370),
.Y(n_3016)
);

OAI22xp5_ASAP7_75t_L g3017 ( 
.A1(n_2892),
.A2(n_2497),
.B1(n_2043),
.B2(n_2463),
.Y(n_3017)
);

BUFx2_ASAP7_75t_L g3018 ( 
.A(n_2848),
.Y(n_3018)
);

INVx4_ASAP7_75t_L g3019 ( 
.A(n_2783),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2726),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2848),
.B(n_2881),
.Y(n_3021)
);

BUFx6f_ASAP7_75t_L g3022 ( 
.A(n_2776),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2827),
.Y(n_3023)
);

AOI21xp5_ASAP7_75t_L g3024 ( 
.A1(n_2777),
.A2(n_2516),
.B(n_2080),
.Y(n_3024)
);

OAI21xp5_ASAP7_75t_L g3025 ( 
.A1(n_2738),
.A2(n_2455),
.B(n_2220),
.Y(n_3025)
);

OR2x6_ASAP7_75t_L g3026 ( 
.A(n_2843),
.B(n_2441),
.Y(n_3026)
);

AND2x2_ASAP7_75t_L g3027 ( 
.A(n_2866),
.B(n_2842),
.Y(n_3027)
);

O2A1O1Ixp33_ASAP7_75t_L g3028 ( 
.A1(n_2868),
.A2(n_2890),
.B(n_2735),
.C(n_2715),
.Y(n_3028)
);

INVx2_ASAP7_75t_L g3029 ( 
.A(n_2786),
.Y(n_3029)
);

NOR3xp33_ASAP7_75t_L g3030 ( 
.A(n_2715),
.B(n_2404),
.C(n_2388),
.Y(n_3030)
);

NOR2x1_ASAP7_75t_L g3031 ( 
.A(n_2824),
.B(n_2392),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2735),
.B(n_2810),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2810),
.B(n_2399),
.Y(n_3033)
);

AOI21xp5_ASAP7_75t_L g3034 ( 
.A1(n_2864),
.A2(n_2080),
.B(n_2076),
.Y(n_3034)
);

OAI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2853),
.A2(n_2463),
.B1(n_2441),
.B2(n_2015),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_2868),
.B(n_2368),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2807),
.B(n_2399),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2739),
.Y(n_3038)
);

INVxp67_ASAP7_75t_R g3039 ( 
.A(n_2729),
.Y(n_3039)
);

NOR2xp67_ASAP7_75t_L g3040 ( 
.A(n_2746),
.B(n_2301),
.Y(n_3040)
);

BUFx6f_ASAP7_75t_L g3041 ( 
.A(n_2776),
.Y(n_3041)
);

NAND3xp33_ASAP7_75t_L g3042 ( 
.A(n_2718),
.B(n_2059),
.C(n_2243),
.Y(n_3042)
);

AOI22x1_ASAP7_75t_L g3043 ( 
.A1(n_2747),
.A2(n_2368),
.B1(n_2381),
.B2(n_2440),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2788),
.B(n_2487),
.Y(n_3044)
);

AOI21xp5_ASAP7_75t_L g3045 ( 
.A1(n_2864),
.A2(n_2076),
.B(n_2475),
.Y(n_3045)
);

AND2x4_ASAP7_75t_L g3046 ( 
.A(n_2797),
.B(n_2817),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2864),
.A2(n_2076),
.B(n_2490),
.Y(n_3047)
);

AOI21xp5_ASAP7_75t_L g3048 ( 
.A1(n_2864),
.A2(n_2216),
.B(n_2085),
.Y(n_3048)
);

CKINVDCx5p33_ASAP7_75t_R g3049 ( 
.A(n_2762),
.Y(n_3049)
);

OAI22xp5_ASAP7_75t_L g3050 ( 
.A1(n_2820),
.A2(n_2010),
.B1(n_2192),
.B2(n_2243),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_SL g3051 ( 
.A(n_2847),
.B(n_2381),
.Y(n_3051)
);

INVx6_ASAP7_75t_L g3052 ( 
.A(n_2783),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2807),
.B(n_2429),
.Y(n_3053)
);

OAI22xp5_ASAP7_75t_L g3054 ( 
.A1(n_2820),
.A2(n_2192),
.B1(n_2243),
.B2(n_2488),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2829),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2744),
.Y(n_3056)
);

O2A1O1Ixp33_ASAP7_75t_L g3057 ( 
.A1(n_2836),
.A2(n_2192),
.B(n_2098),
.C(n_2493),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2858),
.B(n_2429),
.Y(n_3058)
);

HB1xp67_ASAP7_75t_L g3059 ( 
.A(n_2839),
.Y(n_3059)
);

NOR2xp67_ASAP7_75t_SL g3060 ( 
.A(n_2896),
.B(n_2301),
.Y(n_3060)
);

AND2x4_ASAP7_75t_SL g3061 ( 
.A(n_2732),
.B(n_2381),
.Y(n_3061)
);

OA21x2_ASAP7_75t_L g3062 ( 
.A1(n_2841),
.A2(n_2435),
.B(n_2430),
.Y(n_3062)
);

O2A1O1Ixp33_ASAP7_75t_L g3063 ( 
.A1(n_2836),
.A2(n_2098),
.B(n_1589),
.C(n_1598),
.Y(n_3063)
);

O2A1O1Ixp33_ASAP7_75t_L g3064 ( 
.A1(n_2718),
.A2(n_1589),
.B(n_1598),
.C(n_1596),
.Y(n_3064)
);

OAI22xp5_ASAP7_75t_L g3065 ( 
.A1(n_2728),
.A2(n_2243),
.B1(n_2338),
.B2(n_2309),
.Y(n_3065)
);

INVxp67_ASAP7_75t_L g3066 ( 
.A(n_2770),
.Y(n_3066)
);

AOI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2896),
.A2(n_2085),
.B(n_2309),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2858),
.B(n_2430),
.Y(n_3068)
);

NAND2x1p5_ASAP7_75t_L g3069 ( 
.A(n_2896),
.B(n_2293),
.Y(n_3069)
);

NOR2x1_ASAP7_75t_L g3070 ( 
.A(n_2824),
.B(n_2435),
.Y(n_3070)
);

CKINVDCx5p33_ASAP7_75t_R g3071 ( 
.A(n_2844),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2812),
.B(n_2459),
.Y(n_3072)
);

OAI21xp33_ASAP7_75t_L g3073 ( 
.A1(n_2888),
.A2(n_2472),
.B(n_2459),
.Y(n_3073)
);

AOI22xp5_ASAP7_75t_L g3074 ( 
.A1(n_2728),
.A2(n_2376),
.B1(n_2401),
.B2(n_2214),
.Y(n_3074)
);

AOI21xp5_ASAP7_75t_L g3075 ( 
.A1(n_2896),
.A2(n_2085),
.B(n_2338),
.Y(n_3075)
);

O2A1O1Ixp33_ASAP7_75t_SL g3076 ( 
.A1(n_2812),
.A2(n_2474),
.B(n_2502),
.C(n_2472),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2750),
.Y(n_3077)
);

AOI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2823),
.A2(n_2085),
.B(n_2362),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2823),
.B(n_2474),
.Y(n_3079)
);

A2O1A1Ixp33_ASAP7_75t_L g3080 ( 
.A1(n_2888),
.A2(n_2199),
.B(n_2362),
.C(n_2243),
.Y(n_3080)
);

NAND3xp33_ASAP7_75t_L g3081 ( 
.A(n_2869),
.B(n_2513),
.C(n_2502),
.Y(n_3081)
);

INVx2_ASAP7_75t_L g3082 ( 
.A(n_2752),
.Y(n_3082)
);

AOI21xp5_ASAP7_75t_L g3083 ( 
.A1(n_2843),
.A2(n_2085),
.B(n_2041),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2847),
.B(n_2381),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2859),
.B(n_2513),
.Y(n_3085)
);

OAI22xp5_ASAP7_75t_L g3086 ( 
.A1(n_2747),
.A2(n_2199),
.B1(n_2300),
.B2(n_2293),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2840),
.A2(n_2041),
.B(n_2293),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_SL g3088 ( 
.A(n_2859),
.B(n_2797),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2850),
.A2(n_2659),
.B(n_2214),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2840),
.A2(n_2717),
.B(n_2869),
.Y(n_3090)
);

A2O1A1Ixp33_ASAP7_75t_L g3091 ( 
.A1(n_2884),
.A2(n_2034),
.B(n_2523),
.C(n_2521),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2753),
.Y(n_3092)
);

NAND3xp33_ASAP7_75t_L g3093 ( 
.A(n_2884),
.B(n_2523),
.C(n_2521),
.Y(n_3093)
);

OAI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2734),
.A2(n_2840),
.B1(n_2756),
.B2(n_2760),
.Y(n_3094)
);

OAI22xp5_ASAP7_75t_L g3095 ( 
.A1(n_2734),
.A2(n_2764),
.B1(n_2768),
.B2(n_2754),
.Y(n_3095)
);

OAI21x1_ASAP7_75t_L g3096 ( 
.A1(n_3078),
.A2(n_2755),
.B(n_2727),
.Y(n_3096)
);

OAI21x1_ASAP7_75t_SL g3097 ( 
.A1(n_2953),
.A2(n_2771),
.B(n_2793),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2918),
.B(n_3007),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2957),
.Y(n_3099)
);

INVxp67_ASAP7_75t_SL g3100 ( 
.A(n_2970),
.Y(n_3100)
);

OAI21x1_ASAP7_75t_L g3101 ( 
.A1(n_3083),
.A2(n_2755),
.B(n_2727),
.Y(n_3101)
);

O2A1O1Ixp5_ASAP7_75t_SL g3102 ( 
.A1(n_2959),
.A2(n_2809),
.B(n_2814),
.C(n_2799),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2911),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2981),
.Y(n_3104)
);

OAI22xp5_ASAP7_75t_L g3105 ( 
.A1(n_2942),
.A2(n_2734),
.B1(n_2819),
.B2(n_2815),
.Y(n_3105)
);

AOI21xp5_ASAP7_75t_L g3106 ( 
.A1(n_2905),
.A2(n_2928),
.B(n_2929),
.Y(n_3106)
);

BUFx2_ASAP7_75t_L g3107 ( 
.A(n_2933),
.Y(n_3107)
);

AO21x2_ASAP7_75t_L g3108 ( 
.A1(n_2956),
.A2(n_2821),
.B(n_1976),
.Y(n_3108)
);

INVx4_ASAP7_75t_L g3109 ( 
.A(n_2910),
.Y(n_3109)
);

AO31x2_ASAP7_75t_L g3110 ( 
.A1(n_3004),
.A2(n_2832),
.A3(n_2787),
.B(n_2898),
.Y(n_3110)
);

OAI21x1_ASAP7_75t_L g3111 ( 
.A1(n_2971),
.A2(n_2897),
.B(n_2887),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2923),
.A2(n_2897),
.B(n_2887),
.Y(n_3112)
);

OAI21xp5_ASAP7_75t_L g3113 ( 
.A1(n_2952),
.A2(n_2850),
.B(n_2831),
.Y(n_3113)
);

OAI22xp5_ASAP7_75t_L g3114 ( 
.A1(n_2952),
.A2(n_2791),
.B1(n_2732),
.B2(n_2860),
.Y(n_3114)
);

AOI21xp5_ASAP7_75t_L g3115 ( 
.A1(n_2977),
.A2(n_2872),
.B(n_2855),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_3032),
.B(n_2900),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_SL g3117 ( 
.A1(n_3028),
.A2(n_2894),
.B(n_2867),
.Y(n_3117)
);

A2O1A1Ixp33_ASAP7_75t_L g3118 ( 
.A1(n_2921),
.A2(n_2875),
.B(n_2872),
.C(n_2855),
.Y(n_3118)
);

OAI21x1_ASAP7_75t_L g3119 ( 
.A1(n_2966),
.A2(n_2782),
.B(n_2765),
.Y(n_3119)
);

INVx1_ASAP7_75t_L g3120 ( 
.A(n_2982),
.Y(n_3120)
);

AO21x1_ASAP7_75t_L g3121 ( 
.A1(n_3095),
.A2(n_2898),
.B(n_2832),
.Y(n_3121)
);

AO31x2_ASAP7_75t_L g3122 ( 
.A1(n_3080),
.A2(n_2787),
.A3(n_1966),
.B(n_2160),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_3029),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2958),
.A2(n_2876),
.B(n_2850),
.Y(n_3124)
);

OAI21x1_ASAP7_75t_L g3125 ( 
.A1(n_3011),
.A2(n_2782),
.B(n_2765),
.Y(n_3125)
);

AND2x2_ASAP7_75t_SL g3126 ( 
.A(n_2980),
.B(n_2778),
.Y(n_3126)
);

AOI21xp5_ASAP7_75t_L g3127 ( 
.A1(n_2960),
.A2(n_2850),
.B(n_2041),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_3057),
.A2(n_2041),
.B(n_2300),
.Y(n_3128)
);

O2A1O1Ixp5_ASAP7_75t_SL g3129 ( 
.A1(n_2937),
.A2(n_2798),
.B(n_2091),
.C(n_2101),
.Y(n_3129)
);

OA21x2_ASAP7_75t_L g3130 ( 
.A1(n_3090),
.A2(n_2160),
.B(n_2157),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_3027),
.B(n_2798),
.Y(n_3131)
);

OAI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_2931),
.A2(n_2791),
.B1(n_2886),
.B2(n_2880),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2935),
.B(n_2774),
.Y(n_3133)
);

OAI21x1_ASAP7_75t_SL g3134 ( 
.A1(n_2950),
.A2(n_2165),
.B(n_2157),
.Y(n_3134)
);

OAI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_3064),
.A2(n_2831),
.B(n_2774),
.Y(n_3135)
);

BUFx10_ASAP7_75t_L g3136 ( 
.A(n_2972),
.Y(n_3136)
);

BUFx6f_ASAP7_75t_L g3137 ( 
.A(n_2939),
.Y(n_3137)
);

NAND2x1_ASAP7_75t_L g3138 ( 
.A(n_2919),
.B(n_2774),
.Y(n_3138)
);

OAI21xp5_ASAP7_75t_L g3139 ( 
.A1(n_3042),
.A2(n_2831),
.B(n_2774),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2994),
.Y(n_3140)
);

OAI21x1_ASAP7_75t_L g3141 ( 
.A1(n_3087),
.A2(n_2100),
.B(n_2091),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_3077),
.Y(n_3142)
);

INVx2_ASAP7_75t_SL g3143 ( 
.A(n_2920),
.Y(n_3143)
);

OAI21xp33_ASAP7_75t_SL g3144 ( 
.A1(n_3012),
.A2(n_2177),
.B(n_2165),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2975),
.B(n_2831),
.Y(n_3145)
);

OA21x2_ASAP7_75t_L g3146 ( 
.A1(n_3042),
.A2(n_2188),
.B(n_2177),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_3020),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_SL g3148 ( 
.A(n_3060),
.B(n_3021),
.Y(n_3148)
);

BUFx2_ASAP7_75t_L g3149 ( 
.A(n_2933),
.Y(n_3149)
);

AND2x4_ASAP7_75t_L g3150 ( 
.A(n_3018),
.B(n_2300),
.Y(n_3150)
);

OAI21x1_ASAP7_75t_L g3151 ( 
.A1(n_3048),
.A2(n_2101),
.B(n_2100),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_2978),
.A2(n_2346),
.B(n_2300),
.Y(n_3152)
);

OAI21x1_ASAP7_75t_L g3153 ( 
.A1(n_2932),
.A2(n_3047),
.B(n_3045),
.Y(n_3153)
);

OAI21xp5_ASAP7_75t_L g3154 ( 
.A1(n_2940),
.A2(n_2017),
.B(n_2517),
.Y(n_3154)
);

NOR2xp67_ASAP7_75t_L g3155 ( 
.A(n_3066),
.B(n_2034),
.Y(n_3155)
);

NOR4xp25_ASAP7_75t_L g3156 ( 
.A(n_2979),
.B(n_34),
.C(n_29),
.D(n_33),
.Y(n_3156)
);

OAI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2974),
.A2(n_3063),
.B(n_3025),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_3038),
.Y(n_3158)
);

OAI22xp5_ASAP7_75t_L g3159 ( 
.A1(n_3015),
.A2(n_2353),
.B1(n_2363),
.B2(n_2346),
.Y(n_3159)
);

AOI21xp5_ASAP7_75t_L g3160 ( 
.A1(n_3034),
.A2(n_2353),
.B(n_2346),
.Y(n_3160)
);

OAI21x1_ASAP7_75t_L g3161 ( 
.A1(n_3067),
.A2(n_2137),
.B(n_2101),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3056),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2992),
.A2(n_3024),
.B(n_3089),
.Y(n_3163)
);

AOI21xp5_ASAP7_75t_L g3164 ( 
.A1(n_2979),
.A2(n_2353),
.B(n_2346),
.Y(n_3164)
);

NAND3xp33_ASAP7_75t_L g3165 ( 
.A(n_2934),
.B(n_1600),
.C(n_1596),
.Y(n_3165)
);

OAI21x1_ASAP7_75t_L g3166 ( 
.A1(n_3075),
.A2(n_2161),
.B(n_2137),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3092),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_3039),
.B(n_2353),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2990),
.A2(n_2517),
.B1(n_2376),
.B2(n_2401),
.Y(n_3169)
);

AO31x2_ASAP7_75t_L g3170 ( 
.A1(n_2996),
.A2(n_2188),
.A3(n_2197),
.B(n_2194),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_3082),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3055),
.Y(n_3172)
);

AOI221xp5_ASAP7_75t_SL g3173 ( 
.A1(n_3054),
.A2(n_2363),
.B1(n_1965),
.B2(n_35),
.C(n_33),
.Y(n_3173)
);

AO21x2_ASAP7_75t_L g3174 ( 
.A1(n_2991),
.A2(n_2197),
.B(n_2194),
.Y(n_3174)
);

OAI21x1_ASAP7_75t_L g3175 ( 
.A1(n_3065),
.A2(n_2161),
.B(n_2137),
.Y(n_3175)
);

BUFx8_ASAP7_75t_SL g3176 ( 
.A(n_2955),
.Y(n_3176)
);

AO21x1_ASAP7_75t_L g3177 ( 
.A1(n_2986),
.A2(n_2916),
.B(n_2941),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2997),
.B(n_34),
.Y(n_3178)
);

INVx3_ASAP7_75t_L g3179 ( 
.A(n_3046),
.Y(n_3179)
);

AO31x2_ASAP7_75t_L g3180 ( 
.A1(n_3091),
.A2(n_2198),
.A3(n_1629),
.B(n_1643),
.Y(n_3180)
);

OAI21x1_ASAP7_75t_L g3181 ( 
.A1(n_3043),
.A2(n_2163),
.B(n_2161),
.Y(n_3181)
);

AOI21xp5_ASAP7_75t_SL g3182 ( 
.A1(n_2925),
.A2(n_3050),
.B(n_3009),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2909),
.B(n_2017),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_2998),
.Y(n_3184)
);

OAI21x1_ASAP7_75t_L g3185 ( 
.A1(n_2984),
.A2(n_2985),
.B(n_2912),
.Y(n_3185)
);

AND2x4_ASAP7_75t_L g3186 ( 
.A(n_2901),
.B(n_2363),
.Y(n_3186)
);

OAI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2949),
.A2(n_2017),
.B(n_2517),
.Y(n_3187)
);

OAI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_3015),
.A2(n_2363),
.B1(n_2198),
.B2(n_2034),
.Y(n_3188)
);

BUFx6f_ASAP7_75t_L g3189 ( 
.A(n_2939),
.Y(n_3189)
);

OAI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2949),
.A2(n_2017),
.B(n_2517),
.Y(n_3190)
);

OAI21xp5_ASAP7_75t_L g3191 ( 
.A1(n_2951),
.A2(n_2017),
.B(n_2376),
.Y(n_3191)
);

NOR2xp67_ASAP7_75t_SL g3192 ( 
.A(n_2967),
.B(n_2431),
.Y(n_3192)
);

OAI21x1_ASAP7_75t_L g3193 ( 
.A1(n_2907),
.A2(n_3062),
.B(n_3086),
.Y(n_3193)
);

OAI21x1_ASAP7_75t_L g3194 ( 
.A1(n_3062),
.A2(n_2167),
.B(n_2163),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2915),
.B(n_1640),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_3014),
.B(n_1651),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_2954),
.B(n_35),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_3016),
.B(n_1657),
.Y(n_3198)
);

BUFx6f_ASAP7_75t_L g3199 ( 
.A(n_2939),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_2913),
.B(n_37),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_L g3201 ( 
.A1(n_3069),
.A2(n_2167),
.B(n_1629),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2965),
.B(n_39),
.Y(n_3202)
);

AO31x2_ASAP7_75t_L g3203 ( 
.A1(n_3017),
.A2(n_1665),
.A3(n_1657),
.B(n_1604),
.Y(n_3203)
);

AOI221x1_ASAP7_75t_L g3204 ( 
.A1(n_3030),
.A2(n_1485),
.B1(n_1476),
.B2(n_43),
.C(n_40),
.Y(n_3204)
);

OAI21x1_ASAP7_75t_L g3205 ( 
.A1(n_3069),
.A2(n_1604),
.B(n_1600),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_SL g3206 ( 
.A(n_2924),
.B(n_2431),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_3059),
.B(n_42),
.Y(n_3207)
);

OAI21x1_ASAP7_75t_L g3208 ( 
.A1(n_3074),
.A2(n_1610),
.B(n_1485),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2936),
.B(n_43),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2906),
.B(n_44),
.Y(n_3210)
);

INVxp67_ASAP7_75t_SL g3211 ( 
.A(n_3081),
.Y(n_3211)
);

AOI21xp5_ASAP7_75t_L g3212 ( 
.A1(n_3076),
.A2(n_2477),
.B(n_2444),
.Y(n_3212)
);

OAI21x1_ASAP7_75t_L g3213 ( 
.A1(n_3074),
.A2(n_1610),
.B(n_1476),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2919),
.B(n_1665),
.Y(n_3214)
);

NOR4xp25_ASAP7_75t_L g3215 ( 
.A(n_2973),
.B(n_3010),
.C(n_2963),
.D(n_2962),
.Y(n_3215)
);

INVx1_ASAP7_75t_L g3216 ( 
.A(n_2922),
.Y(n_3216)
);

OAI22xp5_ASAP7_75t_L g3217 ( 
.A1(n_2968),
.A2(n_2444),
.B1(n_2464),
.B2(n_2437),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2927),
.B(n_46),
.Y(n_3218)
);

AND3x2_ASAP7_75t_L g3219 ( 
.A(n_3008),
.B(n_47),
.C(n_48),
.Y(n_3219)
);

OAI21xp33_ASAP7_75t_L g3220 ( 
.A1(n_2968),
.A2(n_1569),
.B(n_1573),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2919),
.B(n_49),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_3073),
.A2(n_3093),
.B(n_3081),
.Y(n_3222)
);

CKINVDCx12_ASAP7_75t_R g3223 ( 
.A(n_3085),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2930),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3073),
.B(n_3093),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_L g3226 ( 
.A1(n_2944),
.A2(n_2401),
.B1(n_2125),
.B2(n_1558),
.Y(n_3226)
);

OAI21x1_ASAP7_75t_L g3227 ( 
.A1(n_3072),
.A2(n_1532),
.B(n_1513),
.Y(n_3227)
);

OAI21x1_ASAP7_75t_L g3228 ( 
.A1(n_3079),
.A2(n_1532),
.B(n_1513),
.Y(n_3228)
);

O2A1O1Ixp5_ASAP7_75t_L g3229 ( 
.A1(n_2946),
.A2(n_1541),
.B(n_1530),
.C(n_1532),
.Y(n_3229)
);

NAND3xp33_ASAP7_75t_SL g3230 ( 
.A(n_3002),
.B(n_1982),
.C(n_1980),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2938),
.Y(n_3231)
);

AOI21x1_ASAP7_75t_L g3232 ( 
.A1(n_3036),
.A2(n_1572),
.B(n_1492),
.Y(n_3232)
);

AO31x2_ASAP7_75t_L g3233 ( 
.A1(n_3094),
.A2(n_2057),
.A3(n_2051),
.B(n_2125),
.Y(n_3233)
);

OAI21x1_ASAP7_75t_L g3234 ( 
.A1(n_3037),
.A2(n_1534),
.B(n_1513),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_2904),
.B(n_49),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2943),
.Y(n_3236)
);

AOI221x1_ASAP7_75t_L g3237 ( 
.A1(n_2917),
.A2(n_53),
.B1(n_50),
.B2(n_52),
.C(n_54),
.Y(n_3237)
);

BUFx2_ASAP7_75t_L g3238 ( 
.A(n_3046),
.Y(n_3238)
);

BUFx2_ASAP7_75t_SL g3239 ( 
.A(n_2908),
.Y(n_3239)
);

OAI21x1_ASAP7_75t_L g3240 ( 
.A1(n_3053),
.A2(n_1534),
.B(n_1492),
.Y(n_3240)
);

AO31x2_ASAP7_75t_L g3241 ( 
.A1(n_3035),
.A2(n_3033),
.A3(n_3068),
.B(n_3058),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_2993),
.A2(n_2477),
.B(n_2444),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_2910),
.Y(n_3243)
);

OAI21x1_ASAP7_75t_L g3244 ( 
.A1(n_3031),
.A2(n_1534),
.B(n_1492),
.Y(n_3244)
);

AOI21x1_ASAP7_75t_L g3245 ( 
.A1(n_3070),
.A2(n_1594),
.B(n_1572),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_2904),
.B(n_50),
.Y(n_3246)
);

OAI21x1_ASAP7_75t_L g3247 ( 
.A1(n_2951),
.A2(n_2969),
.B(n_2926),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_2945),
.B(n_55),
.Y(n_3248)
);

INVx2_ASAP7_75t_SL g3249 ( 
.A(n_2910),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2961),
.Y(n_3250)
);

AOI211x1_ASAP7_75t_L g3251 ( 
.A1(n_3088),
.A2(n_3051),
.B(n_3084),
.C(n_2964),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2983),
.B(n_55),
.Y(n_3252)
);

NAND3xp33_ASAP7_75t_SL g3253 ( 
.A(n_3049),
.B(n_56),
.C(n_57),
.Y(n_3253)
);

AO21x1_ASAP7_75t_L g3254 ( 
.A1(n_2999),
.A2(n_56),
.B(n_57),
.Y(n_3254)
);

CKINVDCx5p33_ASAP7_75t_R g3255 ( 
.A(n_2947),
.Y(n_3255)
);

OAI21x1_ASAP7_75t_L g3256 ( 
.A1(n_3003),
.A2(n_1594),
.B(n_1572),
.Y(n_3256)
);

AOI21xp5_ASAP7_75t_L g3257 ( 
.A1(n_3026),
.A2(n_2477),
.B(n_2464),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2987),
.B(n_58),
.Y(n_3258)
);

INVx2_ASAP7_75t_SL g3259 ( 
.A(n_2967),
.Y(n_3259)
);

AOI221xp5_ASAP7_75t_L g3260 ( 
.A1(n_3001),
.A2(n_1558),
.B1(n_1570),
.B2(n_1567),
.C(n_1547),
.Y(n_3260)
);

OAI21xp5_ASAP7_75t_L g3261 ( 
.A1(n_2976),
.A2(n_2401),
.B(n_2125),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_L g3262 ( 
.A(n_3013),
.B(n_59),
.Y(n_3262)
);

INVx4_ASAP7_75t_L g3263 ( 
.A(n_2988),
.Y(n_3263)
);

AO21x1_ASAP7_75t_L g3264 ( 
.A1(n_3005),
.A2(n_59),
.B(n_60),
.Y(n_3264)
);

OAI21x1_ASAP7_75t_L g3265 ( 
.A1(n_3023),
.A2(n_1594),
.B(n_1456),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_SL g3266 ( 
.A(n_2914),
.B(n_3006),
.Y(n_3266)
);

AOI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3000),
.A2(n_2948),
.B1(n_2903),
.B2(n_2976),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_3026),
.A2(n_2464),
.B(n_2437),
.Y(n_3268)
);

OAI21xp5_ASAP7_75t_L g3269 ( 
.A1(n_2948),
.A2(n_2125),
.B(n_1494),
.Y(n_3269)
);

NAND2x1p5_ASAP7_75t_L g3270 ( 
.A(n_2903),
.B(n_2437),
.Y(n_3270)
);

BUFx6f_ASAP7_75t_L g3271 ( 
.A(n_2967),
.Y(n_3271)
);

OAI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3044),
.A2(n_3040),
.B(n_2914),
.Y(n_3272)
);

INVx2_ASAP7_75t_L g3273 ( 
.A(n_2988),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_SL g3274 ( 
.A(n_3019),
.B(n_3071),
.Y(n_3274)
);

OAI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_3019),
.A2(n_2125),
.B(n_1456),
.Y(n_3275)
);

AO31x2_ASAP7_75t_L g3276 ( 
.A1(n_2995),
.A2(n_2057),
.A3(n_2051),
.B(n_2125),
.Y(n_3276)
);

OAI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2989),
.A2(n_2477),
.B1(n_2464),
.B2(n_66),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_3061),
.A2(n_2057),
.B(n_2051),
.Y(n_3278)
);

AND2x2_ASAP7_75t_SL g3279 ( 
.A(n_2988),
.B(n_3022),
.Y(n_3279)
);

OAI21x1_ASAP7_75t_L g3280 ( 
.A1(n_3022),
.A2(n_1456),
.B(n_1436),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_3022),
.A2(n_2057),
.B(n_2051),
.Y(n_3281)
);

OAI21x1_ASAP7_75t_L g3282 ( 
.A1(n_3041),
.A2(n_1469),
.B(n_1436),
.Y(n_3282)
);

OAI21x1_ASAP7_75t_L g3283 ( 
.A1(n_3041),
.A2(n_1469),
.B(n_1436),
.Y(n_3283)
);

INVx1_ASAP7_75t_L g3284 ( 
.A(n_3041),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3052),
.B(n_61),
.Y(n_3285)
);

OAI21x1_ASAP7_75t_L g3286 ( 
.A1(n_3052),
.A2(n_1469),
.B(n_1481),
.Y(n_3286)
);

BUFx3_ASAP7_75t_L g3287 ( 
.A(n_2933),
.Y(n_3287)
);

OAI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2918),
.A2(n_61),
.B(n_64),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_2934),
.B(n_64),
.Y(n_3289)
);

INVx3_ASAP7_75t_L g3290 ( 
.A(n_3046),
.Y(n_3290)
);

NAND2x1p5_ASAP7_75t_L g3291 ( 
.A(n_3060),
.B(n_1547),
.Y(n_3291)
);

AOI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_2902),
.A2(n_1558),
.B(n_1547),
.Y(n_3292)
);

OAI21x1_ASAP7_75t_L g3293 ( 
.A1(n_3078),
.A2(n_1558),
.B(n_1547),
.Y(n_3293)
);

INVx2_ASAP7_75t_SL g3294 ( 
.A(n_2920),
.Y(n_3294)
);

AO31x2_ASAP7_75t_L g3295 ( 
.A1(n_3083),
.A2(n_70),
.A3(n_68),
.B(n_69),
.Y(n_3295)
);

NAND2xp5_ASAP7_75t_L g3296 ( 
.A(n_2953),
.B(n_68),
.Y(n_3296)
);

INVx2_ASAP7_75t_SL g3297 ( 
.A(n_2920),
.Y(n_3297)
);

OAI21x1_ASAP7_75t_L g3298 ( 
.A1(n_3078),
.A2(n_1558),
.B(n_1547),
.Y(n_3298)
);

O2A1O1Ixp5_ASAP7_75t_L g3299 ( 
.A1(n_2918),
.A2(n_71),
.B(n_69),
.C(n_70),
.Y(n_3299)
);

A2O1A1Ixp33_ASAP7_75t_L g3300 ( 
.A1(n_3288),
.A2(n_75),
.B(n_72),
.C(n_74),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3104),
.Y(n_3301)
);

AOI21xp5_ASAP7_75t_L g3302 ( 
.A1(n_3222),
.A2(n_1570),
.B(n_1567),
.Y(n_3302)
);

OR2x2_ASAP7_75t_L g3303 ( 
.A(n_3100),
.B(n_72),
.Y(n_3303)
);

OAI21xp5_ASAP7_75t_L g3304 ( 
.A1(n_3288),
.A2(n_74),
.B(n_76),
.Y(n_3304)
);

O2A1O1Ixp33_ASAP7_75t_L g3305 ( 
.A1(n_3296),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_3305)
);

AO32x2_ASAP7_75t_L g3306 ( 
.A1(n_3132),
.A2(n_77),
.A3(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3120),
.Y(n_3307)
);

A2O1A1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_3296),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3098),
.B(n_82),
.Y(n_3309)
);

OAI21x1_ASAP7_75t_L g3310 ( 
.A1(n_3153),
.A2(n_281),
.B(n_276),
.Y(n_3310)
);

INVx2_ASAP7_75t_SL g3311 ( 
.A(n_3137),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_3116),
.B(n_84),
.Y(n_3312)
);

OAI21x1_ASAP7_75t_L g3313 ( 
.A1(n_3193),
.A2(n_287),
.B(n_285),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_3106),
.A2(n_1570),
.B(n_1567),
.Y(n_3314)
);

AOI21x1_ASAP7_75t_L g3315 ( 
.A1(n_3235),
.A2(n_84),
.B(n_85),
.Y(n_3315)
);

OAI21xp5_ASAP7_75t_SL g3316 ( 
.A1(n_3219),
.A2(n_85),
.B(n_86),
.Y(n_3316)
);

OAI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_3105),
.A2(n_86),
.B(n_87),
.Y(n_3317)
);

AOI221xp5_ASAP7_75t_SL g3318 ( 
.A1(n_3105),
.A2(n_3221),
.B1(n_3289),
.B2(n_3277),
.C(n_3114),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3157),
.A2(n_3127),
.B(n_3113),
.Y(n_3319)
);

OAI22xp5_ASAP7_75t_L g3320 ( 
.A1(n_3118),
.A2(n_1570),
.B1(n_1584),
.B2(n_1567),
.Y(n_3320)
);

AOI221x1_ASAP7_75t_L g3321 ( 
.A1(n_3221),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.C(n_91),
.Y(n_3321)
);

OA21x2_ASAP7_75t_L g3322 ( 
.A1(n_3177),
.A2(n_90),
.B(n_91),
.Y(n_3322)
);

AOI21x1_ASAP7_75t_L g3323 ( 
.A1(n_3235),
.A2(n_92),
.B(n_94),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3140),
.Y(n_3324)
);

BUFx6f_ASAP7_75t_L g3325 ( 
.A(n_3137),
.Y(n_3325)
);

A2O1A1Ixp33_ASAP7_75t_L g3326 ( 
.A1(n_3113),
.A2(n_96),
.B(n_94),
.C(n_95),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3157),
.A2(n_1570),
.B(n_1567),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_3147),
.Y(n_3328)
);

NAND3xp33_ASAP7_75t_L g3329 ( 
.A(n_3237),
.B(n_1611),
.C(n_1584),
.Y(n_3329)
);

AND2x4_ASAP7_75t_L g3330 ( 
.A(n_3179),
.B(n_95),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_3139),
.A2(n_1611),
.B(n_1584),
.Y(n_3331)
);

OAI21x1_ASAP7_75t_L g3332 ( 
.A1(n_3292),
.A2(n_294),
.B(n_292),
.Y(n_3332)
);

AO32x2_ASAP7_75t_L g3333 ( 
.A1(n_3132),
.A2(n_98),
.A3(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_3139),
.A2(n_1611),
.B(n_1584),
.Y(n_3334)
);

O2A1O1Ixp33_ASAP7_75t_L g3335 ( 
.A1(n_3253),
.A2(n_102),
.B(n_99),
.C(n_100),
.Y(n_3335)
);

INVx2_ASAP7_75t_L g3336 ( 
.A(n_3142),
.Y(n_3336)
);

AOI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_3156),
.A2(n_1611),
.B(n_1584),
.Y(n_3337)
);

AND2x2_ASAP7_75t_L g3338 ( 
.A(n_3238),
.B(n_103),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3172),
.B(n_103),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_L g3340 ( 
.A(n_3137),
.Y(n_3340)
);

BUFx6f_ASAP7_75t_L g3341 ( 
.A(n_3189),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_3171),
.Y(n_3342)
);

OAI21x1_ASAP7_75t_L g3343 ( 
.A1(n_3293),
.A2(n_3298),
.B(n_3185),
.Y(n_3343)
);

OAI21xp5_ASAP7_75t_L g3344 ( 
.A1(n_3299),
.A2(n_104),
.B(n_105),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_3145),
.B(n_105),
.Y(n_3345)
);

AO31x2_ASAP7_75t_L g3346 ( 
.A1(n_3128),
.A2(n_109),
.A3(n_107),
.B(n_108),
.Y(n_3346)
);

A2O1A1Ixp33_ASAP7_75t_L g3347 ( 
.A1(n_3154),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_3347)
);

OAI21x1_ASAP7_75t_L g3348 ( 
.A1(n_3163),
.A2(n_296),
.B(n_295),
.Y(n_3348)
);

NOR2xp67_ASAP7_75t_L g3349 ( 
.A(n_3103),
.B(n_111),
.Y(n_3349)
);

A2O1A1Ixp33_ASAP7_75t_L g3350 ( 
.A1(n_3154),
.A2(n_115),
.B(n_112),
.C(n_114),
.Y(n_3350)
);

BUFx2_ASAP7_75t_L g3351 ( 
.A(n_3184),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_SL g3352 ( 
.A(n_3148),
.B(n_1611),
.Y(n_3352)
);

OR2x2_ASAP7_75t_L g3353 ( 
.A(n_3099),
.B(n_116),
.Y(n_3353)
);

AOI21xp5_ASAP7_75t_L g3354 ( 
.A1(n_3156),
.A2(n_1512),
.B(n_1511),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3158),
.Y(n_3355)
);

AO31x2_ASAP7_75t_L g3356 ( 
.A1(n_3204),
.A2(n_118),
.A3(n_116),
.B(n_117),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3133),
.B(n_117),
.Y(n_3357)
);

O2A1O1Ixp33_ASAP7_75t_L g3358 ( 
.A1(n_3277),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_3358)
);

NAND2xp5_ASAP7_75t_L g3359 ( 
.A(n_3123),
.B(n_119),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_SL g3360 ( 
.A(n_3176),
.B(n_1510),
.Y(n_3360)
);

BUFx6f_ASAP7_75t_L g3361 ( 
.A(n_3189),
.Y(n_3361)
);

CKINVDCx20_ASAP7_75t_R g3362 ( 
.A(n_3255),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3162),
.Y(n_3363)
);

OAI21x1_ASAP7_75t_L g3364 ( 
.A1(n_3227),
.A2(n_311),
.B(n_304),
.Y(n_3364)
);

OAI21x1_ASAP7_75t_L g3365 ( 
.A1(n_3228),
.A2(n_316),
.B(n_314),
.Y(n_3365)
);

OAI21x1_ASAP7_75t_L g3366 ( 
.A1(n_3234),
.A2(n_321),
.B(n_317),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3216),
.B(n_121),
.Y(n_3367)
);

AO32x2_ASAP7_75t_L g3368 ( 
.A1(n_3114),
.A2(n_122),
.A3(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_3368)
);

OAI21x1_ASAP7_75t_L g3369 ( 
.A1(n_3129),
.A2(n_325),
.B(n_323),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3167),
.Y(n_3370)
);

NAND3x1_ASAP7_75t_L g3371 ( 
.A(n_3267),
.B(n_123),
.C(n_124),
.Y(n_3371)
);

OAI21x1_ASAP7_75t_L g3372 ( 
.A1(n_3194),
.A2(n_3124),
.B(n_3212),
.Y(n_3372)
);

OAI21x1_ASAP7_75t_L g3373 ( 
.A1(n_3102),
.A2(n_329),
.B(n_327),
.Y(n_3373)
);

AND2x2_ASAP7_75t_L g3374 ( 
.A(n_3290),
.B(n_125),
.Y(n_3374)
);

AO31x2_ASAP7_75t_L g3375 ( 
.A1(n_3121),
.A2(n_126),
.A3(n_127),
.B(n_128),
.Y(n_3375)
);

BUFx6f_ASAP7_75t_SL g3376 ( 
.A(n_3287),
.Y(n_3376)
);

INVxp67_ASAP7_75t_L g3377 ( 
.A(n_3189),
.Y(n_3377)
);

NOR2xp67_ASAP7_75t_L g3378 ( 
.A(n_3259),
.B(n_126),
.Y(n_3378)
);

OAI21x1_ASAP7_75t_L g3379 ( 
.A1(n_3208),
.A2(n_335),
.B(n_333),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3224),
.Y(n_3380)
);

HB1xp67_ASAP7_75t_L g3381 ( 
.A(n_3214),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_3199),
.Y(n_3382)
);

NOR3xp33_ASAP7_75t_L g3383 ( 
.A(n_3214),
.B(n_127),
.C(n_128),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3250),
.Y(n_3384)
);

A2O1A1Ixp33_ASAP7_75t_L g3385 ( 
.A1(n_3138),
.A2(n_129),
.B(n_130),
.C(n_131),
.Y(n_3385)
);

AO31x2_ASAP7_75t_L g3386 ( 
.A1(n_3217),
.A2(n_131),
.A3(n_132),
.B(n_133),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3231),
.Y(n_3387)
);

INVx6_ASAP7_75t_L g3388 ( 
.A(n_3136),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_3290),
.Y(n_3389)
);

OAI22xp33_ASAP7_75t_L g3390 ( 
.A1(n_3148),
.A2(n_1526),
.B1(n_1524),
.B2(n_1523),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3236),
.Y(n_3391)
);

AOI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_3135),
.A2(n_1512),
.B(n_1511),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3246),
.Y(n_3393)
);

NAND2xp33_ASAP7_75t_R g3394 ( 
.A(n_3107),
.B(n_133),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3246),
.Y(n_3395)
);

AOI221xp5_ASAP7_75t_SL g3396 ( 
.A1(n_3200),
.A2(n_134),
.B1(n_135),
.B2(n_137),
.C(n_139),
.Y(n_3396)
);

OA21x2_ASAP7_75t_L g3397 ( 
.A1(n_3125),
.A2(n_3096),
.B(n_3272),
.Y(n_3397)
);

OAI21xp5_ASAP7_75t_L g3398 ( 
.A1(n_3215),
.A2(n_135),
.B(n_139),
.Y(n_3398)
);

AO21x2_ASAP7_75t_L g3399 ( 
.A1(n_3117),
.A2(n_140),
.B(n_141),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3131),
.B(n_140),
.Y(n_3400)
);

INVx2_ASAP7_75t_SL g3401 ( 
.A(n_3199),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_3225),
.A2(n_1512),
.B(n_1511),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3149),
.B(n_142),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3241),
.B(n_143),
.Y(n_3404)
);

AO21x2_ASAP7_75t_L g3405 ( 
.A1(n_3165),
.A2(n_143),
.B(n_144),
.Y(n_3405)
);

OAI21x1_ASAP7_75t_L g3406 ( 
.A1(n_3213),
.A2(n_337),
.B(n_336),
.Y(n_3406)
);

BUFx2_ASAP7_75t_R g3407 ( 
.A(n_3274),
.Y(n_3407)
);

INVx2_ASAP7_75t_L g3408 ( 
.A(n_3284),
.Y(n_3408)
);

AO21x1_ASAP7_75t_L g3409 ( 
.A1(n_3207),
.A2(n_146),
.B(n_147),
.Y(n_3409)
);

OAI21xp5_ASAP7_75t_L g3410 ( 
.A1(n_3215),
.A2(n_148),
.B(n_150),
.Y(n_3410)
);

O2A1O1Ixp5_ASAP7_75t_L g3411 ( 
.A1(n_3254),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3273),
.Y(n_3412)
);

AO31x2_ASAP7_75t_L g3413 ( 
.A1(n_3217),
.A2(n_151),
.A3(n_152),
.B(n_153),
.Y(n_3413)
);

CKINVDCx11_ASAP7_75t_R g3414 ( 
.A(n_3136),
.Y(n_3414)
);

INVx4_ASAP7_75t_L g3415 ( 
.A(n_3199),
.Y(n_3415)
);

AOI221xp5_ASAP7_75t_L g3416 ( 
.A1(n_3264),
.A2(n_153),
.B1(n_154),
.B2(n_156),
.C(n_157),
.Y(n_3416)
);

AO31x2_ASAP7_75t_L g3417 ( 
.A1(n_3159),
.A2(n_157),
.A3(n_159),
.B(n_160),
.Y(n_3417)
);

NAND2xp5_ASAP7_75t_L g3418 ( 
.A(n_3241),
.B(n_160),
.Y(n_3418)
);

AOI21xp5_ASAP7_75t_L g3419 ( 
.A1(n_3225),
.A2(n_3182),
.B(n_3211),
.Y(n_3419)
);

NAND3xp33_ASAP7_75t_L g3420 ( 
.A(n_3173),
.B(n_1512),
.C(n_1511),
.Y(n_3420)
);

BUFx3_ASAP7_75t_L g3421 ( 
.A(n_3271),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3241),
.B(n_161),
.Y(n_3422)
);

AOI21xp5_ASAP7_75t_L g3423 ( 
.A1(n_3165),
.A2(n_1512),
.B(n_1511),
.Y(n_3423)
);

OA22x2_ASAP7_75t_L g3424 ( 
.A1(n_3272),
.A2(n_161),
.B1(n_168),
.B2(n_169),
.Y(n_3424)
);

CKINVDCx8_ASAP7_75t_R g3425 ( 
.A(n_3239),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_3247),
.B(n_169),
.Y(n_3426)
);

AND2x4_ASAP7_75t_L g3427 ( 
.A(n_3101),
.B(n_170),
.Y(n_3427)
);

AOI21xp5_ASAP7_75t_L g3428 ( 
.A1(n_3187),
.A2(n_1523),
.B(n_1518),
.Y(n_3428)
);

INVx5_ASAP7_75t_L g3429 ( 
.A(n_3271),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_SL g3430 ( 
.A(n_3126),
.B(n_1518),
.Y(n_3430)
);

BUFx10_ASAP7_75t_L g3431 ( 
.A(n_3271),
.Y(n_3431)
);

OAI22xp5_ASAP7_75t_L g3432 ( 
.A1(n_3169),
.A2(n_1526),
.B1(n_1524),
.B2(n_1523),
.Y(n_3432)
);

AOI21xp5_ASAP7_75t_L g3433 ( 
.A1(n_3187),
.A2(n_1523),
.B(n_1518),
.Y(n_3433)
);

BUFx3_ASAP7_75t_L g3434 ( 
.A(n_3143),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3295),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_3119),
.Y(n_3436)
);

AOI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_3190),
.A2(n_1523),
.B(n_1518),
.Y(n_3437)
);

OAI21x1_ASAP7_75t_L g3438 ( 
.A1(n_3151),
.A2(n_345),
.B(n_342),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3097),
.Y(n_3439)
);

AO21x1_ASAP7_75t_L g3440 ( 
.A1(n_3206),
.A2(n_170),
.B(n_171),
.Y(n_3440)
);

NAND2x1p5_ASAP7_75t_L g3441 ( 
.A(n_3192),
.B(n_1518),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_3294),
.Y(n_3442)
);

OAI21x1_ASAP7_75t_L g3443 ( 
.A1(n_3141),
.A2(n_348),
.B(n_347),
.Y(n_3443)
);

OAI22x1_ASAP7_75t_L g3444 ( 
.A1(n_3197),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3186),
.Y(n_3445)
);

AO31x2_ASAP7_75t_L g3446 ( 
.A1(n_3159),
.A2(n_172),
.A3(n_173),
.B(n_174),
.Y(n_3446)
);

AO31x2_ASAP7_75t_L g3447 ( 
.A1(n_3188),
.A2(n_177),
.A3(n_178),
.B(n_180),
.Y(n_3447)
);

INVx3_ASAP7_75t_L g3448 ( 
.A(n_3109),
.Y(n_3448)
);

INVxp67_ASAP7_75t_L g3449 ( 
.A(n_3297),
.Y(n_3449)
);

AOI21xp5_ASAP7_75t_L g3450 ( 
.A1(n_3190),
.A2(n_1526),
.B(n_1524),
.Y(n_3450)
);

CKINVDCx11_ASAP7_75t_R g3451 ( 
.A(n_3109),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3195),
.B(n_178),
.Y(n_3452)
);

AOI21xp5_ASAP7_75t_L g3453 ( 
.A1(n_3275),
.A2(n_1526),
.B(n_1524),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3195),
.B(n_180),
.Y(n_3454)
);

INVx1_ASAP7_75t_SL g3455 ( 
.A(n_3279),
.Y(n_3455)
);

AOI22xp5_ASAP7_75t_L g3456 ( 
.A1(n_3266),
.A2(n_1526),
.B1(n_1524),
.B2(n_1529),
.Y(n_3456)
);

OAI21x1_ASAP7_75t_L g3457 ( 
.A1(n_3134),
.A2(n_3112),
.B(n_3175),
.Y(n_3457)
);

AOI21x1_ASAP7_75t_L g3458 ( 
.A1(n_3115),
.A2(n_183),
.B(n_184),
.Y(n_3458)
);

AOI21xp5_ASAP7_75t_L g3459 ( 
.A1(n_3191),
.A2(n_1510),
.B(n_1529),
.Y(n_3459)
);

AND2x2_ASAP7_75t_L g3460 ( 
.A(n_3168),
.B(n_3186),
.Y(n_3460)
);

INVx2_ASAP7_75t_SL g3461 ( 
.A(n_3243),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3183),
.B(n_183),
.Y(n_3462)
);

BUFx6f_ASAP7_75t_L g3463 ( 
.A(n_3414),
.Y(n_3463)
);

OAI21x1_ASAP7_75t_L g3464 ( 
.A1(n_3372),
.A2(n_3111),
.B(n_3130),
.Y(n_3464)
);

OAI22xp5_ASAP7_75t_L g3465 ( 
.A1(n_3329),
.A2(n_3251),
.B1(n_3164),
.B2(n_3191),
.Y(n_3465)
);

AND2x4_ASAP7_75t_L g3466 ( 
.A(n_3445),
.B(n_3381),
.Y(n_3466)
);

AOI21xp5_ASAP7_75t_L g3467 ( 
.A1(n_3327),
.A2(n_3130),
.B(n_3146),
.Y(n_3467)
);

INVx3_ASAP7_75t_L g3468 ( 
.A(n_3448),
.Y(n_3468)
);

NOR2xp33_ASAP7_75t_L g3469 ( 
.A(n_3388),
.B(n_3266),
.Y(n_3469)
);

AOI21x1_ASAP7_75t_L g3470 ( 
.A1(n_3426),
.A2(n_3418),
.B(n_3404),
.Y(n_3470)
);

AOI21x1_ASAP7_75t_L g3471 ( 
.A1(n_3422),
.A2(n_3218),
.B(n_3210),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3408),
.Y(n_3472)
);

NOR2xp33_ASAP7_75t_L g3473 ( 
.A(n_3393),
.B(n_3209),
.Y(n_3473)
);

OAI21x1_ASAP7_75t_L g3474 ( 
.A1(n_3343),
.A2(n_3160),
.B(n_3240),
.Y(n_3474)
);

OAI21x1_ASAP7_75t_SL g3475 ( 
.A1(n_3419),
.A2(n_3252),
.B(n_3248),
.Y(n_3475)
);

AND2x2_ASAP7_75t_L g3476 ( 
.A(n_3351),
.B(n_3243),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3301),
.Y(n_3477)
);

AO21x2_ASAP7_75t_L g3478 ( 
.A1(n_3435),
.A2(n_3174),
.B(n_3108),
.Y(n_3478)
);

OR2x6_ASAP7_75t_L g3479 ( 
.A(n_3319),
.B(n_3257),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3301),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3307),
.Y(n_3481)
);

OAI21x1_ASAP7_75t_L g3482 ( 
.A1(n_3457),
.A2(n_3268),
.B(n_3166),
.Y(n_3482)
);

HB1xp67_ASAP7_75t_L g3483 ( 
.A(n_3395),
.Y(n_3483)
);

OAI21x1_ASAP7_75t_L g3484 ( 
.A1(n_3313),
.A2(n_3161),
.B(n_3152),
.Y(n_3484)
);

OAI22xp5_ASAP7_75t_L g3485 ( 
.A1(n_3300),
.A2(n_3202),
.B1(n_3178),
.B2(n_3183),
.Y(n_3485)
);

OR2x6_ASAP7_75t_L g3486 ( 
.A(n_3392),
.B(n_3261),
.Y(n_3486)
);

AND2x4_ASAP7_75t_L g3487 ( 
.A(n_3389),
.B(n_3412),
.Y(n_3487)
);

OAI21x1_ASAP7_75t_L g3488 ( 
.A1(n_3302),
.A2(n_3229),
.B(n_3242),
.Y(n_3488)
);

NAND2x1p5_ASAP7_75t_L g3489 ( 
.A(n_3429),
.B(n_3146),
.Y(n_3489)
);

OAI21x1_ASAP7_75t_L g3490 ( 
.A1(n_3402),
.A2(n_3198),
.B(n_3196),
.Y(n_3490)
);

OAI22xp5_ASAP7_75t_SL g3491 ( 
.A1(n_3425),
.A2(n_3223),
.B1(n_3285),
.B2(n_3270),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_L g3492 ( 
.A1(n_3304),
.A2(n_3220),
.B1(n_3261),
.B2(n_3230),
.Y(n_3492)
);

INVx3_ASAP7_75t_L g3493 ( 
.A(n_3448),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3324),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3324),
.Y(n_3495)
);

A2O1A1Ixp33_ASAP7_75t_L g3496 ( 
.A1(n_3305),
.A2(n_3410),
.B(n_3398),
.C(n_3316),
.Y(n_3496)
);

XOR2xp5_ASAP7_75t_L g3497 ( 
.A(n_3362),
.B(n_3407),
.Y(n_3497)
);

BUFx2_ASAP7_75t_L g3498 ( 
.A(n_3377),
.Y(n_3498)
);

AND2x2_ASAP7_75t_SL g3499 ( 
.A(n_3322),
.B(n_3383),
.Y(n_3499)
);

HB1xp67_ASAP7_75t_L g3500 ( 
.A(n_3328),
.Y(n_3500)
);

O2A1O1Ixp33_ASAP7_75t_SL g3501 ( 
.A1(n_3326),
.A2(n_3258),
.B(n_3262),
.C(n_3249),
.Y(n_3501)
);

OAI21x1_ASAP7_75t_L g3502 ( 
.A1(n_3436),
.A2(n_3198),
.B(n_3196),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3328),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3355),
.Y(n_3504)
);

AOI21xp5_ASAP7_75t_L g3505 ( 
.A1(n_3428),
.A2(n_3269),
.B(n_3144),
.Y(n_3505)
);

OAI21x1_ASAP7_75t_L g3506 ( 
.A1(n_3314),
.A2(n_3244),
.B(n_3270),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3355),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3363),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3363),
.Y(n_3509)
);

AO21x2_ASAP7_75t_L g3510 ( 
.A1(n_3435),
.A2(n_3174),
.B(n_3108),
.Y(n_3510)
);

AOI21x1_ASAP7_75t_L g3511 ( 
.A1(n_3315),
.A2(n_3155),
.B(n_3245),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_3433),
.A2(n_3269),
.B(n_3188),
.Y(n_3512)
);

OA21x2_ASAP7_75t_L g3513 ( 
.A1(n_3318),
.A2(n_3173),
.B(n_3265),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_3370),
.Y(n_3514)
);

AO31x2_ASAP7_75t_L g3515 ( 
.A1(n_3439),
.A2(n_3263),
.A3(n_3281),
.B(n_3278),
.Y(n_3515)
);

CKINVDCx5p33_ASAP7_75t_R g3516 ( 
.A(n_3376),
.Y(n_3516)
);

INVx3_ASAP7_75t_L g3517 ( 
.A(n_3421),
.Y(n_3517)
);

OAI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_3317),
.A2(n_3411),
.B(n_3308),
.Y(n_3518)
);

AO21x2_ASAP7_75t_L g3519 ( 
.A1(n_3323),
.A2(n_3205),
.B(n_3201),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3370),
.Y(n_3520)
);

AOI21xp5_ASAP7_75t_L g3521 ( 
.A1(n_3437),
.A2(n_3260),
.B(n_3291),
.Y(n_3521)
);

OAI21x1_ASAP7_75t_L g3522 ( 
.A1(n_3331),
.A2(n_3282),
.B(n_3280),
.Y(n_3522)
);

NAND3xp33_ASAP7_75t_L g3523 ( 
.A(n_3416),
.B(n_3226),
.C(n_3263),
.Y(n_3523)
);

AND2x4_ASAP7_75t_L g3524 ( 
.A(n_3461),
.B(n_3170),
.Y(n_3524)
);

OAI21x1_ASAP7_75t_L g3525 ( 
.A1(n_3334),
.A2(n_3283),
.B(n_3286),
.Y(n_3525)
);

OAI21x1_ASAP7_75t_L g3526 ( 
.A1(n_3310),
.A2(n_3181),
.B(n_3232),
.Y(n_3526)
);

OR2x6_ASAP7_75t_L g3527 ( 
.A(n_3459),
.B(n_3291),
.Y(n_3527)
);

INVx2_ASAP7_75t_L g3528 ( 
.A(n_3380),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3380),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3384),
.Y(n_3530)
);

AOI221xp5_ASAP7_75t_L g3531 ( 
.A1(n_3396),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.C(n_189),
.Y(n_3531)
);

AND2x2_ASAP7_75t_L g3532 ( 
.A(n_3460),
.B(n_3203),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3336),
.Y(n_3533)
);

OAI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_3344),
.A2(n_3150),
.B(n_3295),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3342),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3387),
.Y(n_3536)
);

NAND2x1p5_ASAP7_75t_L g3537 ( 
.A(n_3429),
.B(n_3150),
.Y(n_3537)
);

AOI21xp5_ASAP7_75t_L g3538 ( 
.A1(n_3450),
.A2(n_3256),
.B(n_3295),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3391),
.Y(n_3539)
);

OAI21x1_ASAP7_75t_L g3540 ( 
.A1(n_3458),
.A2(n_3203),
.B(n_3122),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3303),
.Y(n_3541)
);

OAI21x1_ASAP7_75t_L g3542 ( 
.A1(n_3348),
.A2(n_3203),
.B(n_3122),
.Y(n_3542)
);

OR2x2_ASAP7_75t_L g3543 ( 
.A(n_3397),
.B(n_3122),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3353),
.Y(n_3544)
);

NAND3xp33_ASAP7_75t_L g3545 ( 
.A(n_3321),
.B(n_187),
.C(n_190),
.Y(n_3545)
);

AND2x4_ASAP7_75t_L g3546 ( 
.A(n_3427),
.B(n_3170),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3339),
.Y(n_3547)
);

NOR4xp25_ASAP7_75t_L g3548 ( 
.A(n_3335),
.B(n_190),
.C(n_191),
.D(n_192),
.Y(n_3548)
);

OR2x2_ASAP7_75t_L g3549 ( 
.A(n_3397),
.B(n_3455),
.Y(n_3549)
);

O2A1O1Ixp33_ASAP7_75t_SL g3550 ( 
.A1(n_3385),
.A2(n_191),
.B(n_192),
.C(n_195),
.Y(n_3550)
);

OAI21x1_ASAP7_75t_L g3551 ( 
.A1(n_3364),
.A2(n_3170),
.B(n_3180),
.Y(n_3551)
);

INVx1_ASAP7_75t_L g3552 ( 
.A(n_3346),
.Y(n_3552)
);

OAI22xp5_ASAP7_75t_L g3553 ( 
.A1(n_3424),
.A2(n_3276),
.B1(n_3233),
.B2(n_3110),
.Y(n_3553)
);

OAI21x1_ASAP7_75t_L g3554 ( 
.A1(n_3365),
.A2(n_3180),
.B(n_3233),
.Y(n_3554)
);

OAI21x1_ASAP7_75t_L g3555 ( 
.A1(n_3366),
.A2(n_3180),
.B(n_3233),
.Y(n_3555)
);

O2A1O1Ixp33_ASAP7_75t_L g3556 ( 
.A1(n_3358),
.A2(n_198),
.B(n_199),
.C(n_201),
.Y(n_3556)
);

CKINVDCx16_ASAP7_75t_R g3557 ( 
.A(n_3394),
.Y(n_3557)
);

INVx8_ASAP7_75t_L g3558 ( 
.A(n_3376),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3346),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3346),
.Y(n_3560)
);

OAI21x1_ASAP7_75t_L g3561 ( 
.A1(n_3373),
.A2(n_3110),
.B(n_3276),
.Y(n_3561)
);

NOR2xp33_ASAP7_75t_L g3562 ( 
.A(n_3388),
.B(n_198),
.Y(n_3562)
);

NOR2x1_ASAP7_75t_SL g3563 ( 
.A(n_3429),
.B(n_3110),
.Y(n_3563)
);

CKINVDCx6p67_ASAP7_75t_R g3564 ( 
.A(n_3451),
.Y(n_3564)
);

OAI22xp5_ASAP7_75t_L g3565 ( 
.A1(n_3420),
.A2(n_3350),
.B1(n_3347),
.B2(n_3371),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3367),
.Y(n_3566)
);

OAI21x1_ASAP7_75t_L g3567 ( 
.A1(n_3379),
.A2(n_3276),
.B(n_201),
.Y(n_3567)
);

OAI21x1_ASAP7_75t_L g3568 ( 
.A1(n_3406),
.A2(n_199),
.B(n_202),
.Y(n_3568)
);

INVx5_ASAP7_75t_L g3569 ( 
.A(n_3330),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3309),
.B(n_203),
.Y(n_3570)
);

INVxp67_ASAP7_75t_L g3571 ( 
.A(n_3322),
.Y(n_3571)
);

INVx2_ASAP7_75t_L g3572 ( 
.A(n_3311),
.Y(n_3572)
);

OAI21x1_ASAP7_75t_L g3573 ( 
.A1(n_3453),
.A2(n_203),
.B(n_204),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3382),
.Y(n_3574)
);

INVx1_ASAP7_75t_SL g3575 ( 
.A(n_3325),
.Y(n_3575)
);

AOI22x1_ASAP7_75t_L g3576 ( 
.A1(n_3444),
.A2(n_205),
.B1(n_206),
.B2(n_207),
.Y(n_3576)
);

AO22x2_ASAP7_75t_L g3577 ( 
.A1(n_3320),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_3577)
);

BUFx2_ASAP7_75t_SL g3578 ( 
.A(n_3378),
.Y(n_3578)
);

INVx1_ASAP7_75t_L g3579 ( 
.A(n_3359),
.Y(n_3579)
);

NOR2xp67_ASAP7_75t_L g3580 ( 
.A(n_3449),
.B(n_208),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3312),
.B(n_211),
.Y(n_3581)
);

BUFx2_ASAP7_75t_L g3582 ( 
.A(n_3415),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3375),
.Y(n_3583)
);

AO21x2_ASAP7_75t_L g3584 ( 
.A1(n_3462),
.A2(n_212),
.B(n_213),
.Y(n_3584)
);

OAI21xp5_ASAP7_75t_L g3585 ( 
.A1(n_3352),
.A2(n_212),
.B(n_214),
.Y(n_3585)
);

AO31x2_ASAP7_75t_L g3586 ( 
.A1(n_3440),
.A2(n_214),
.A3(n_217),
.B(n_218),
.Y(n_3586)
);

AOI221xp5_ASAP7_75t_L g3587 ( 
.A1(n_3409),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.C(n_225),
.Y(n_3587)
);

OA21x2_ASAP7_75t_L g3588 ( 
.A1(n_3345),
.A2(n_219),
.B(n_220),
.Y(n_3588)
);

OAI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3349),
.A2(n_226),
.B(n_227),
.Y(n_3589)
);

NAND2x1p5_ASAP7_75t_L g3590 ( 
.A(n_3430),
.B(n_1441),
.Y(n_3590)
);

BUFx2_ASAP7_75t_SL g3591 ( 
.A(n_3434),
.Y(n_3591)
);

NAND2x1p5_ASAP7_75t_L g3592 ( 
.A(n_3569),
.B(n_3325),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3500),
.Y(n_3593)
);

AO21x2_ASAP7_75t_L g3594 ( 
.A1(n_3571),
.A2(n_3357),
.B(n_3399),
.Y(n_3594)
);

OA21x2_ASAP7_75t_L g3595 ( 
.A1(n_3571),
.A2(n_3454),
.B(n_3452),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_SL g3596 ( 
.A1(n_3496),
.A2(n_3330),
.B(n_3390),
.Y(n_3596)
);

AOI211xp5_ASAP7_75t_L g3597 ( 
.A1(n_3518),
.A2(n_3338),
.B(n_3374),
.C(n_3403),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3500),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_3477),
.Y(n_3599)
);

AOI21xp5_ASAP7_75t_L g3600 ( 
.A1(n_3499),
.A2(n_3337),
.B(n_3405),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3518),
.A2(n_3360),
.B(n_3423),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3481),
.Y(n_3602)
);

BUFx8_ASAP7_75t_L g3603 ( 
.A(n_3463),
.Y(n_3603)
);

OA21x2_ASAP7_75t_L g3604 ( 
.A1(n_3552),
.A2(n_3369),
.B(n_3443),
.Y(n_3604)
);

BUFx4f_ASAP7_75t_SL g3605 ( 
.A(n_3564),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_SL g3606 ( 
.A(n_3557),
.B(n_3325),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3494),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3476),
.B(n_3442),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3543),
.A2(n_3438),
.B(n_3332),
.Y(n_3609)
);

OA21x2_ASAP7_75t_L g3610 ( 
.A1(n_3559),
.A2(n_3560),
.B(n_3583),
.Y(n_3610)
);

INVx6_ASAP7_75t_L g3611 ( 
.A(n_3558),
.Y(n_3611)
);

OAI21x1_ASAP7_75t_L g3612 ( 
.A1(n_3464),
.A2(n_3432),
.B(n_3354),
.Y(n_3612)
);

AOI21xp5_ASAP7_75t_L g3613 ( 
.A1(n_3565),
.A2(n_3456),
.B(n_3401),
.Y(n_3613)
);

INVx1_ASAP7_75t_SL g3614 ( 
.A(n_3591),
.Y(n_3614)
);

OAI21x1_ASAP7_75t_L g3615 ( 
.A1(n_3482),
.A2(n_3441),
.B(n_3400),
.Y(n_3615)
);

CKINVDCx16_ASAP7_75t_R g3616 ( 
.A(n_3463),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3495),
.Y(n_3617)
);

INVx1_ASAP7_75t_L g3618 ( 
.A(n_3503),
.Y(n_3618)
);

BUFx3_ASAP7_75t_L g3619 ( 
.A(n_3558),
.Y(n_3619)
);

OAI21x1_ASAP7_75t_L g3620 ( 
.A1(n_3561),
.A2(n_3375),
.B(n_3306),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3579),
.B(n_3375),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_3565),
.A2(n_3368),
.B(n_3306),
.Y(n_3622)
);

INVx2_ASAP7_75t_L g3623 ( 
.A(n_3480),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3504),
.Y(n_3624)
);

OAI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_3548),
.A2(n_3306),
.B(n_3333),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_3556),
.A2(n_3368),
.B(n_3333),
.Y(n_3626)
);

INVx1_ASAP7_75t_L g3627 ( 
.A(n_3507),
.Y(n_3627)
);

AO21x2_ASAP7_75t_L g3628 ( 
.A1(n_3563),
.A2(n_3368),
.B(n_3333),
.Y(n_3628)
);

OA21x2_ASAP7_75t_L g3629 ( 
.A1(n_3549),
.A2(n_3540),
.B(n_3474),
.Y(n_3629)
);

AND2x4_ASAP7_75t_L g3630 ( 
.A(n_3479),
.B(n_3386),
.Y(n_3630)
);

AND2x4_ASAP7_75t_L g3631 ( 
.A(n_3479),
.B(n_3386),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3542),
.A2(n_3386),
.B(n_3413),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3514),
.Y(n_3633)
);

NOR2xp33_ASAP7_75t_L g3634 ( 
.A(n_3470),
.B(n_3340),
.Y(n_3634)
);

AND2x4_ASAP7_75t_L g3635 ( 
.A(n_3479),
.B(n_3413),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3508),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3509),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3473),
.B(n_3417),
.Y(n_3638)
);

AO21x2_ASAP7_75t_L g3639 ( 
.A1(n_3475),
.A2(n_3446),
.B(n_3417),
.Y(n_3639)
);

INVx2_ASAP7_75t_L g3640 ( 
.A(n_3528),
.Y(n_3640)
);

AOI21x1_ASAP7_75t_L g3641 ( 
.A1(n_3582),
.A2(n_3471),
.B(n_3580),
.Y(n_3641)
);

BUFx6f_ASAP7_75t_L g3642 ( 
.A(n_3463),
.Y(n_3642)
);

AO31x2_ASAP7_75t_L g3643 ( 
.A1(n_3553),
.A2(n_3446),
.A3(n_3356),
.B(n_3447),
.Y(n_3643)
);

INVxp67_ASAP7_75t_L g3644 ( 
.A(n_3483),
.Y(n_3644)
);

OAI21x1_ASAP7_75t_L g3645 ( 
.A1(n_3489),
.A2(n_3446),
.B(n_3431),
.Y(n_3645)
);

AND2x2_ASAP7_75t_L g3646 ( 
.A(n_3498),
.B(n_3487),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3520),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3473),
.B(n_3547),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3489),
.A2(n_3447),
.B(n_3431),
.Y(n_3649)
);

NAND2x1p5_ASAP7_75t_L g3650 ( 
.A(n_3569),
.B(n_3340),
.Y(n_3650)
);

AO21x2_ASAP7_75t_L g3651 ( 
.A1(n_3538),
.A2(n_3356),
.B(n_3447),
.Y(n_3651)
);

AO31x2_ASAP7_75t_L g3652 ( 
.A1(n_3553),
.A2(n_3361),
.A3(n_3341),
.B(n_229),
.Y(n_3652)
);

INVxp67_ASAP7_75t_SL g3653 ( 
.A(n_3483),
.Y(n_3653)
);

INVx1_ASAP7_75t_L g3654 ( 
.A(n_3529),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3566),
.B(n_3341),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_3546),
.B(n_3341),
.Y(n_3656)
);

OAI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_3548),
.A2(n_3361),
.B(n_228),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3472),
.Y(n_3658)
);

HB1xp67_ASAP7_75t_L g3659 ( 
.A(n_3530),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3536),
.Y(n_3660)
);

INVx3_ASAP7_75t_L g3661 ( 
.A(n_3468),
.Y(n_3661)
);

AOI21xp33_ASAP7_75t_SL g3662 ( 
.A1(n_3497),
.A2(n_227),
.B(n_228),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3539),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3533),
.Y(n_3664)
);

BUFx3_ASAP7_75t_L g3665 ( 
.A(n_3516),
.Y(n_3665)
);

INVx2_ASAP7_75t_SL g3666 ( 
.A(n_3517),
.Y(n_3666)
);

AOI21x1_ASAP7_75t_L g3667 ( 
.A1(n_3570),
.A2(n_3361),
.B(n_231),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3502),
.A2(n_230),
.B(n_232),
.Y(n_3668)
);

INVx4_ASAP7_75t_L g3669 ( 
.A(n_3569),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_L g3670 ( 
.A(n_3541),
.B(n_232),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3535),
.Y(n_3671)
);

INVx3_ASAP7_75t_L g3672 ( 
.A(n_3468),
.Y(n_3672)
);

HB1xp67_ASAP7_75t_L g3673 ( 
.A(n_3588),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3466),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3544),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_3570),
.B(n_233),
.Y(n_3676)
);

OR2x2_ASAP7_75t_L g3677 ( 
.A(n_3466),
.B(n_233),
.Y(n_3677)
);

AO21x2_ASAP7_75t_L g3678 ( 
.A1(n_3538),
.A2(n_234),
.B(n_235),
.Y(n_3678)
);

INVx2_ASAP7_75t_L g3679 ( 
.A(n_3524),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3524),
.Y(n_3680)
);

A2O1A1Ixp33_ASAP7_75t_L g3681 ( 
.A1(n_3531),
.A2(n_236),
.B(n_237),
.C(n_238),
.Y(n_3681)
);

OA21x2_ASAP7_75t_L g3682 ( 
.A1(n_3467),
.A2(n_240),
.B(n_241),
.Y(n_3682)
);

INVx3_ASAP7_75t_L g3683 ( 
.A(n_3493),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3532),
.B(n_242),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3581),
.B(n_242),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3554),
.A2(n_243),
.B(n_244),
.Y(n_3686)
);

OAI21x1_ASAP7_75t_L g3687 ( 
.A1(n_3555),
.A2(n_243),
.B(n_244),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3487),
.B(n_245),
.Y(n_3688)
);

OA21x2_ASAP7_75t_L g3689 ( 
.A1(n_3467),
.A2(n_3488),
.B(n_3587),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3545),
.A2(n_245),
.B(n_246),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_3546),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3588),
.Y(n_3692)
);

OAI21x1_ASAP7_75t_L g3693 ( 
.A1(n_3551),
.A2(n_247),
.B(n_248),
.Y(n_3693)
);

INVx1_ASAP7_75t_L g3694 ( 
.A(n_3493),
.Y(n_3694)
);

BUFx3_ASAP7_75t_L g3695 ( 
.A(n_3517),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3575),
.B(n_247),
.Y(n_3696)
);

AOI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_3545),
.A2(n_248),
.B(n_249),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3572),
.B(n_249),
.Y(n_3698)
);

NAND2x1p5_ASAP7_75t_L g3699 ( 
.A(n_3569),
.B(n_250),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_3578),
.Y(n_3700)
);

A2O1A1Ixp33_ASAP7_75t_L g3701 ( 
.A1(n_3531),
.A2(n_251),
.B(n_255),
.C(n_256),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_L g3702 ( 
.A(n_3575),
.B(n_251),
.Y(n_3702)
);

AOI21xp5_ASAP7_75t_L g3703 ( 
.A1(n_3492),
.A2(n_256),
.B(n_257),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3584),
.Y(n_3704)
);

AOI21xp33_ASAP7_75t_L g3705 ( 
.A1(n_3587),
.A2(n_258),
.B(n_260),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3465),
.B(n_260),
.Y(n_3706)
);

AND2x4_ASAP7_75t_L g3707 ( 
.A(n_3515),
.B(n_261),
.Y(n_3707)
);

INVx3_ASAP7_75t_L g3708 ( 
.A(n_3537),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_L g3709 ( 
.A(n_3465),
.B(n_261),
.Y(n_3709)
);

INVx4_ASAP7_75t_R g3710 ( 
.A(n_3614),
.Y(n_3710)
);

OAI21xp5_ASAP7_75t_SL g3711 ( 
.A1(n_3705),
.A2(n_3492),
.B(n_3589),
.Y(n_3711)
);

NOR2x1_ASAP7_75t_L g3712 ( 
.A(n_3606),
.B(n_3469),
.Y(n_3712)
);

OAI21xp33_ASAP7_75t_L g3713 ( 
.A1(n_3625),
.A2(n_3589),
.B(n_3534),
.Y(n_3713)
);

AOI22xp33_ASAP7_75t_L g3714 ( 
.A1(n_3622),
.A2(n_3491),
.B1(n_3486),
.B2(n_3576),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3659),
.Y(n_3715)
);

BUFx5_ASAP7_75t_L g3716 ( 
.A(n_3707),
.Y(n_3716)
);

INVx1_ASAP7_75t_L g3717 ( 
.A(n_3659),
.Y(n_3717)
);

OAI22xp5_ASAP7_75t_L g3718 ( 
.A1(n_3626),
.A2(n_3486),
.B1(n_3577),
.B2(n_3523),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3638),
.B(n_3584),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3599),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3595),
.B(n_3581),
.Y(n_3721)
);

AOI22xp33_ASAP7_75t_L g3722 ( 
.A1(n_3706),
.A2(n_3486),
.B1(n_3534),
.B2(n_3523),
.Y(n_3722)
);

AND2x2_ASAP7_75t_L g3723 ( 
.A(n_3646),
.B(n_3574),
.Y(n_3723)
);

BUFx3_ASAP7_75t_L g3724 ( 
.A(n_3603),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3669),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3669),
.Y(n_3726)
);

BUFx12f_ASAP7_75t_L g3727 ( 
.A(n_3603),
.Y(n_3727)
);

OAI22xp5_ASAP7_75t_L g3728 ( 
.A1(n_3681),
.A2(n_3577),
.B1(n_3527),
.B2(n_3505),
.Y(n_3728)
);

INVx3_ASAP7_75t_L g3729 ( 
.A(n_3642),
.Y(n_3729)
);

CKINVDCx8_ASAP7_75t_R g3730 ( 
.A(n_3616),
.Y(n_3730)
);

INVx1_ASAP7_75t_L g3731 ( 
.A(n_3602),
.Y(n_3731)
);

AOI22xp33_ASAP7_75t_L g3732 ( 
.A1(n_3709),
.A2(n_3513),
.B1(n_3577),
.B2(n_3485),
.Y(n_3732)
);

BUFx2_ASAP7_75t_L g3733 ( 
.A(n_3700),
.Y(n_3733)
);

AOI22xp33_ASAP7_75t_L g3734 ( 
.A1(n_3600),
.A2(n_3513),
.B1(n_3485),
.B2(n_3512),
.Y(n_3734)
);

AOI22xp33_ASAP7_75t_L g3735 ( 
.A1(n_3606),
.A2(n_3512),
.B1(n_3585),
.B2(n_3505),
.Y(n_3735)
);

OAI21xp5_ASAP7_75t_SL g3736 ( 
.A1(n_3703),
.A2(n_3585),
.B(n_3562),
.Y(n_3736)
);

AOI22xp5_ASAP7_75t_L g3737 ( 
.A1(n_3681),
.A2(n_3550),
.B1(n_3501),
.B2(n_3527),
.Y(n_3737)
);

NOR2xp33_ASAP7_75t_L g3738 ( 
.A(n_3605),
.B(n_3611),
.Y(n_3738)
);

AOI22xp33_ASAP7_75t_L g3739 ( 
.A1(n_3689),
.A2(n_3639),
.B1(n_3678),
.B2(n_3697),
.Y(n_3739)
);

OAI22xp5_ASAP7_75t_L g3740 ( 
.A1(n_3701),
.A2(n_3596),
.B1(n_3601),
.B2(n_3700),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3607),
.Y(n_3741)
);

AOI22xp33_ASAP7_75t_L g3742 ( 
.A1(n_3689),
.A2(n_3527),
.B1(n_3573),
.B2(n_3519),
.Y(n_3742)
);

OAI22xp5_ASAP7_75t_L g3743 ( 
.A1(n_3701),
.A2(n_3537),
.B1(n_3590),
.B2(n_3521),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_L g3744 ( 
.A1(n_3689),
.A2(n_3519),
.B1(n_3490),
.B2(n_3568),
.Y(n_3744)
);

AOI22xp33_ASAP7_75t_L g3745 ( 
.A1(n_3639),
.A2(n_3521),
.B1(n_3478),
.B2(n_3510),
.Y(n_3745)
);

OAI21xp5_ASAP7_75t_SL g3746 ( 
.A1(n_3690),
.A2(n_3511),
.B(n_3590),
.Y(n_3746)
);

AOI22xp33_ASAP7_75t_SL g3747 ( 
.A1(n_3657),
.A2(n_3567),
.B1(n_3478),
.B2(n_3510),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3617),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3618),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3678),
.A2(n_3594),
.B1(n_3651),
.B2(n_3628),
.Y(n_3750)
);

OAI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3673),
.A2(n_3586),
.B1(n_3515),
.B2(n_3525),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3624),
.Y(n_3752)
);

AOI22xp33_ASAP7_75t_SL g3753 ( 
.A1(n_3628),
.A2(n_3586),
.B1(n_3484),
.B2(n_3506),
.Y(n_3753)
);

INVxp67_ASAP7_75t_L g3754 ( 
.A(n_3673),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3627),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3594),
.A2(n_3522),
.B1(n_3526),
.B2(n_3586),
.Y(n_3756)
);

INVx1_ASAP7_75t_L g3757 ( 
.A(n_3636),
.Y(n_3757)
);

OAI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3597),
.A2(n_263),
.B1(n_264),
.B2(n_266),
.Y(n_3758)
);

OAI22xp33_ASAP7_75t_L g3759 ( 
.A1(n_3699),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_3759)
);

AND2x2_ASAP7_75t_L g3760 ( 
.A(n_3674),
.B(n_267),
.Y(n_3760)
);

OAI22xp5_ASAP7_75t_L g3761 ( 
.A1(n_3613),
.A2(n_1529),
.B1(n_356),
.B2(n_359),
.Y(n_3761)
);

AOI22xp33_ASAP7_75t_L g3762 ( 
.A1(n_3651),
.A2(n_1496),
.B1(n_1495),
.B2(n_1491),
.Y(n_3762)
);

OAI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3699),
.A2(n_350),
.B1(n_360),
.B2(n_361),
.Y(n_3763)
);

AOI22xp33_ASAP7_75t_L g3764 ( 
.A1(n_3595),
.A2(n_1497),
.B1(n_1496),
.B2(n_1495),
.Y(n_3764)
);

AOI22xp33_ASAP7_75t_L g3765 ( 
.A1(n_3595),
.A2(n_1497),
.B1(n_1496),
.B2(n_1495),
.Y(n_3765)
);

OAI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3641),
.A2(n_365),
.B(n_368),
.Y(n_3766)
);

INVx1_ASAP7_75t_L g3767 ( 
.A(n_3637),
.Y(n_3767)
);

OAI22xp5_ASAP7_75t_L g3768 ( 
.A1(n_3648),
.A2(n_371),
.B1(n_372),
.B2(n_375),
.Y(n_3768)
);

OAI22xp5_ASAP7_75t_L g3769 ( 
.A1(n_3684),
.A2(n_376),
.B1(n_380),
.B2(n_381),
.Y(n_3769)
);

CKINVDCx5p33_ASAP7_75t_R g3770 ( 
.A(n_3603),
.Y(n_3770)
);

OAI22xp33_ASAP7_75t_L g3771 ( 
.A1(n_3662),
.A2(n_391),
.B1(n_392),
.B2(n_394),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3634),
.B(n_398),
.Y(n_3772)
);

OAI22xp5_ASAP7_75t_L g3773 ( 
.A1(n_3611),
.A2(n_400),
.B1(n_402),
.B2(n_405),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3679),
.Y(n_3774)
);

OAI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3692),
.A2(n_3667),
.B1(n_3642),
.B2(n_3605),
.Y(n_3775)
);

AOI22xp33_ASAP7_75t_SL g3776 ( 
.A1(n_3676),
.A2(n_408),
.B1(n_410),
.B2(n_412),
.Y(n_3776)
);

AOI22xp33_ASAP7_75t_L g3777 ( 
.A1(n_3630),
.A2(n_1496),
.B1(n_1495),
.B2(n_1491),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3630),
.A2(n_1496),
.B1(n_1495),
.B2(n_1491),
.Y(n_3778)
);

AND2x2_ASAP7_75t_L g3779 ( 
.A(n_3695),
.B(n_414),
.Y(n_3779)
);

AOI22xp33_ASAP7_75t_L g3780 ( 
.A1(n_3630),
.A2(n_1497),
.B1(n_1491),
.B2(n_1490),
.Y(n_3780)
);

OAI22xp5_ASAP7_75t_L g3781 ( 
.A1(n_3611),
.A2(n_418),
.B1(n_421),
.B2(n_424),
.Y(n_3781)
);

BUFx2_ASAP7_75t_L g3782 ( 
.A(n_3695),
.Y(n_3782)
);

INVx4_ASAP7_75t_L g3783 ( 
.A(n_3642),
.Y(n_3783)
);

HB1xp67_ASAP7_75t_L g3784 ( 
.A(n_3610),
.Y(n_3784)
);

BUFx4f_ASAP7_75t_SL g3785 ( 
.A(n_3665),
.Y(n_3785)
);

OAI21xp33_ASAP7_75t_L g3786 ( 
.A1(n_3631),
.A2(n_427),
.B(n_430),
.Y(n_3786)
);

AOI22xp33_ASAP7_75t_SL g3787 ( 
.A1(n_3676),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3656),
.B(n_3708),
.Y(n_3788)
);

CKINVDCx5p33_ASAP7_75t_R g3789 ( 
.A(n_3665),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3619),
.B(n_3642),
.Y(n_3790)
);

OAI21xp5_ASAP7_75t_L g3791 ( 
.A1(n_3634),
.A2(n_434),
.B(n_436),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3680),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3654),
.Y(n_3793)
);

AOI22xp33_ASAP7_75t_L g3794 ( 
.A1(n_3631),
.A2(n_1497),
.B1(n_1491),
.B2(n_1490),
.Y(n_3794)
);

AOI22xp33_ASAP7_75t_L g3795 ( 
.A1(n_3631),
.A2(n_3635),
.B1(n_3619),
.B2(n_3692),
.Y(n_3795)
);

OAI21xp5_ASAP7_75t_SL g3796 ( 
.A1(n_3685),
.A2(n_441),
.B(n_442),
.Y(n_3796)
);

AOI22xp33_ASAP7_75t_SL g3797 ( 
.A1(n_3685),
.A2(n_443),
.B1(n_1497),
.B2(n_1490),
.Y(n_3797)
);

OAI22xp5_ASAP7_75t_L g3798 ( 
.A1(n_3592),
.A2(n_1490),
.B1(n_1442),
.B2(n_1448),
.Y(n_3798)
);

OAI22xp33_ASAP7_75t_L g3799 ( 
.A1(n_3704),
.A2(n_1441),
.B1(n_1442),
.B2(n_1448),
.Y(n_3799)
);

AOI22xp33_ASAP7_75t_L g3800 ( 
.A1(n_3682),
.A2(n_1441),
.B1(n_1442),
.B2(n_1448),
.Y(n_3800)
);

CKINVDCx20_ASAP7_75t_R g3801 ( 
.A(n_3608),
.Y(n_3801)
);

CKINVDCx5p33_ASAP7_75t_R g3802 ( 
.A(n_3688),
.Y(n_3802)
);

HB1xp67_ASAP7_75t_L g3803 ( 
.A(n_3610),
.Y(n_3803)
);

BUFx12f_ASAP7_75t_L g3804 ( 
.A(n_3677),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_L g3805 ( 
.A1(n_3682),
.A2(n_3704),
.B1(n_3691),
.B2(n_3675),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3682),
.A2(n_1467),
.B1(n_1482),
.B2(n_1489),
.Y(n_3806)
);

HB1xp67_ASAP7_75t_L g3807 ( 
.A(n_3610),
.Y(n_3807)
);

BUFx12f_ASAP7_75t_L g3808 ( 
.A(n_3698),
.Y(n_3808)
);

OAI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3650),
.A2(n_1467),
.B1(n_1482),
.B2(n_1489),
.Y(n_3809)
);

OAI22xp33_ASAP7_75t_L g3810 ( 
.A1(n_3670),
.A2(n_1467),
.B1(n_1482),
.B2(n_1489),
.Y(n_3810)
);

AOI22xp5_ASAP7_75t_L g3811 ( 
.A1(n_3655),
.A2(n_1443),
.B1(n_3621),
.B2(n_3707),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3647),
.Y(n_3812)
);

INVx5_ASAP7_75t_SL g3813 ( 
.A(n_3693),
.Y(n_3813)
);

OAI22xp33_ASAP7_75t_L g3814 ( 
.A1(n_3650),
.A2(n_1443),
.B1(n_3702),
.B2(n_3696),
.Y(n_3814)
);

OAI21xp33_ASAP7_75t_L g3815 ( 
.A1(n_3620),
.A2(n_1443),
.B(n_3632),
.Y(n_3815)
);

INVx1_ASAP7_75t_SL g3816 ( 
.A(n_3666),
.Y(n_3816)
);

AO21x2_ASAP7_75t_L g3817 ( 
.A1(n_3754),
.A2(n_3653),
.B(n_3632),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3716),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3712),
.B(n_3652),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_SL g3820 ( 
.A1(n_3740),
.A2(n_3653),
.B(n_3644),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3720),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3731),
.Y(n_3822)
);

INVx2_ASAP7_75t_L g3823 ( 
.A(n_3716),
.Y(n_3823)
);

INVx3_ASAP7_75t_L g3824 ( 
.A(n_3730),
.Y(n_3824)
);

BUFx3_ASAP7_75t_L g3825 ( 
.A(n_3727),
.Y(n_3825)
);

INVx1_ASAP7_75t_L g3826 ( 
.A(n_3741),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3721),
.B(n_3719),
.Y(n_3827)
);

OA21x2_ASAP7_75t_L g3828 ( 
.A1(n_3750),
.A2(n_3644),
.B(n_3645),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3722),
.B(n_3652),
.Y(n_3829)
);

OA21x2_ASAP7_75t_L g3830 ( 
.A1(n_3739),
.A2(n_3754),
.B(n_3713),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3748),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_3716),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3788),
.B(n_3782),
.Y(n_3833)
);

OA21x2_ASAP7_75t_L g3834 ( 
.A1(n_3784),
.A2(n_3649),
.B(n_3593),
.Y(n_3834)
);

INVxp67_ASAP7_75t_L g3835 ( 
.A(n_3733),
.Y(n_3835)
);

HB1xp67_ASAP7_75t_L g3836 ( 
.A(n_3715),
.Y(n_3836)
);

BUFx3_ASAP7_75t_L g3837 ( 
.A(n_3724),
.Y(n_3837)
);

INVx2_ASAP7_75t_L g3838 ( 
.A(n_3716),
.Y(n_3838)
);

INVxp67_ASAP7_75t_SL g3839 ( 
.A(n_3775),
.Y(n_3839)
);

HB1xp67_ASAP7_75t_L g3840 ( 
.A(n_3717),
.Y(n_3840)
);

OR2x6_ASAP7_75t_L g3841 ( 
.A(n_3725),
.B(n_3687),
.Y(n_3841)
);

BUFx2_ASAP7_75t_L g3842 ( 
.A(n_3783),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_3716),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_3726),
.B(n_3652),
.Y(n_3844)
);

INVx3_ASAP7_75t_L g3845 ( 
.A(n_3783),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3749),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3752),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3716),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3784),
.Y(n_3849)
);

INVx1_ASAP7_75t_L g3850 ( 
.A(n_3755),
.Y(n_3850)
);

INVx1_ASAP7_75t_L g3851 ( 
.A(n_3757),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3767),
.Y(n_3852)
);

INVx3_ASAP7_75t_L g3853 ( 
.A(n_3729),
.Y(n_3853)
);

AO21x2_ASAP7_75t_L g3854 ( 
.A1(n_3803),
.A2(n_3649),
.B(n_3686),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3793),
.Y(n_3855)
);

OAI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3747),
.A2(n_3718),
.B(n_3711),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3812),
.Y(n_3857)
);

INVx1_ASAP7_75t_L g3858 ( 
.A(n_3803),
.Y(n_3858)
);

INVx2_ASAP7_75t_L g3859 ( 
.A(n_3807),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3807),
.Y(n_3860)
);

OR2x6_ASAP7_75t_L g3861 ( 
.A(n_3766),
.B(n_3668),
.Y(n_3861)
);

AND2x4_ASAP7_75t_L g3862 ( 
.A(n_3729),
.B(n_3652),
.Y(n_3862)
);

AND2x2_ASAP7_75t_L g3863 ( 
.A(n_3774),
.B(n_3661),
.Y(n_3863)
);

HB1xp67_ASAP7_75t_L g3864 ( 
.A(n_3816),
.Y(n_3864)
);

AO21x2_ASAP7_75t_L g3865 ( 
.A1(n_3775),
.A2(n_3598),
.B(n_3694),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3792),
.B(n_3683),
.Y(n_3866)
);

NOR2xp33_ASAP7_75t_L g3867 ( 
.A(n_3785),
.B(n_3663),
.Y(n_3867)
);

HB1xp67_ASAP7_75t_L g3868 ( 
.A(n_3751),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3795),
.B(n_3683),
.Y(n_3869)
);

BUFx3_ASAP7_75t_L g3870 ( 
.A(n_3770),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_3813),
.Y(n_3871)
);

OR2x2_ASAP7_75t_L g3872 ( 
.A(n_3805),
.B(n_3643),
.Y(n_3872)
);

INVx2_ASAP7_75t_L g3873 ( 
.A(n_3813),
.Y(n_3873)
);

INVx2_ASAP7_75t_L g3874 ( 
.A(n_3813),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3760),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3723),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3811),
.B(n_3734),
.Y(n_3877)
);

INVx1_ASAP7_75t_L g3878 ( 
.A(n_3710),
.Y(n_3878)
);

OAI21x1_ASAP7_75t_L g3879 ( 
.A1(n_3745),
.A2(n_3629),
.B(n_3661),
.Y(n_3879)
);

OAI211xp5_ASAP7_75t_SL g3880 ( 
.A1(n_3714),
.A2(n_3660),
.B(n_3671),
.C(n_3664),
.Y(n_3880)
);

INVx1_ASAP7_75t_L g3881 ( 
.A(n_3790),
.Y(n_3881)
);

INVxp67_ASAP7_75t_L g3882 ( 
.A(n_3737),
.Y(n_3882)
);

BUFx3_ASAP7_75t_L g3883 ( 
.A(n_3789),
.Y(n_3883)
);

OR2x6_ASAP7_75t_L g3884 ( 
.A(n_3728),
.B(n_3758),
.Y(n_3884)
);

OR2x2_ASAP7_75t_L g3885 ( 
.A(n_3732),
.B(n_3643),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3804),
.Y(n_3886)
);

INVx3_ASAP7_75t_L g3887 ( 
.A(n_3808),
.Y(n_3887)
);

NAND2x1p5_ASAP7_75t_L g3888 ( 
.A(n_3738),
.B(n_3615),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_3736),
.A2(n_3629),
.B(n_3609),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3814),
.Y(n_3890)
);

OR2x2_ASAP7_75t_L g3891 ( 
.A(n_3742),
.B(n_3643),
.Y(n_3891)
);

NOR2xp33_ASAP7_75t_L g3892 ( 
.A(n_3801),
.B(n_3664),
.Y(n_3892)
);

OR2x2_ASAP7_75t_L g3893 ( 
.A(n_3744),
.B(n_3643),
.Y(n_3893)
);

INVx1_ASAP7_75t_SL g3894 ( 
.A(n_3802),
.Y(n_3894)
);

INVx1_ASAP7_75t_L g3895 ( 
.A(n_3814),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3743),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3779),
.Y(n_3897)
);

NAND2xp33_ASAP7_75t_SL g3898 ( 
.A(n_3735),
.B(n_3772),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3753),
.B(n_3672),
.Y(n_3899)
);

AND2x2_ASAP7_75t_L g3900 ( 
.A(n_3753),
.B(n_3672),
.Y(n_3900)
);

BUFx12f_ASAP7_75t_L g3901 ( 
.A(n_3759),
.Y(n_3901)
);

BUFx6f_ASAP7_75t_L g3902 ( 
.A(n_3759),
.Y(n_3902)
);

INVx2_ASAP7_75t_L g3903 ( 
.A(n_3809),
.Y(n_3903)
);

OR2x2_ASAP7_75t_L g3904 ( 
.A(n_3756),
.B(n_3658),
.Y(n_3904)
);

INVx2_ASAP7_75t_L g3905 ( 
.A(n_3798),
.Y(n_3905)
);

HB1xp67_ASAP7_75t_L g3906 ( 
.A(n_3746),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3761),
.Y(n_3907)
);

INVx2_ASAP7_75t_L g3908 ( 
.A(n_3763),
.Y(n_3908)
);

INVx1_ASAP7_75t_SL g3909 ( 
.A(n_3747),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3810),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3810),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3815),
.Y(n_3912)
);

BUFx2_ASAP7_75t_L g3913 ( 
.A(n_3791),
.Y(n_3913)
);

AOI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3771),
.A2(n_3796),
.B1(n_3797),
.B2(n_3786),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3769),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3764),
.Y(n_3916)
);

BUFx4f_ASAP7_75t_SL g3917 ( 
.A(n_3776),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3849),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3842),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3849),
.Y(n_3920)
);

HB1xp67_ASAP7_75t_L g3921 ( 
.A(n_3864),
.Y(n_3921)
);

NOR2xp33_ASAP7_75t_L g3922 ( 
.A(n_3824),
.B(n_3771),
.Y(n_3922)
);

BUFx3_ASAP7_75t_L g3923 ( 
.A(n_3825),
.Y(n_3923)
);

HB1xp67_ASAP7_75t_L g3924 ( 
.A(n_3842),
.Y(n_3924)
);

INVx2_ASAP7_75t_L g3925 ( 
.A(n_3817),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3901),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3878),
.B(n_3629),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3859),
.Y(n_3928)
);

HB1xp67_ASAP7_75t_L g3929 ( 
.A(n_3835),
.Y(n_3929)
);

AND2x2_ASAP7_75t_L g3930 ( 
.A(n_3878),
.B(n_3640),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3859),
.Y(n_3931)
);

INVx3_ASAP7_75t_L g3932 ( 
.A(n_3865),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3858),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3902),
.B(n_3765),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3817),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3833),
.B(n_3824),
.Y(n_3936)
);

INVxp67_ASAP7_75t_SL g3937 ( 
.A(n_3824),
.Y(n_3937)
);

OR2x2_ASAP7_75t_SL g3938 ( 
.A(n_3902),
.B(n_3623),
.Y(n_3938)
);

OR2x2_ASAP7_75t_SL g3939 ( 
.A(n_3902),
.B(n_3623),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3860),
.Y(n_3940)
);

INVx1_ASAP7_75t_SL g3941 ( 
.A(n_3825),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3833),
.B(n_3633),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3817),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3865),
.Y(n_3944)
);

OA21x2_ASAP7_75t_L g3945 ( 
.A1(n_3856),
.A2(n_3800),
.B(n_3806),
.Y(n_3945)
);

BUFx3_ASAP7_75t_L g3946 ( 
.A(n_3901),
.Y(n_3946)
);

INVx1_ASAP7_75t_L g3947 ( 
.A(n_3836),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3840),
.Y(n_3948)
);

INVx1_ASAP7_75t_L g3949 ( 
.A(n_3821),
.Y(n_3949)
);

AO21x2_ASAP7_75t_L g3950 ( 
.A1(n_3820),
.A2(n_3799),
.B(n_3768),
.Y(n_3950)
);

OR2x2_ASAP7_75t_L g3951 ( 
.A(n_3872),
.B(n_3778),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3865),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3834),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3819),
.B(n_3869),
.Y(n_3954)
);

NAND2x1p5_ASAP7_75t_L g3955 ( 
.A(n_3913),
.B(n_3612),
.Y(n_3955)
);

OAI211xp5_ASAP7_75t_L g3956 ( 
.A1(n_3820),
.A2(n_3776),
.B(n_3787),
.C(n_3762),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3834),
.Y(n_3957)
);

INVx1_ASAP7_75t_L g3958 ( 
.A(n_3821),
.Y(n_3958)
);

OR2x2_ASAP7_75t_L g3959 ( 
.A(n_3872),
.B(n_3780),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3853),
.Y(n_3960)
);

INVx3_ASAP7_75t_L g3961 ( 
.A(n_3902),
.Y(n_3961)
);

NOR2xp33_ASAP7_75t_L g3962 ( 
.A(n_3870),
.B(n_3787),
.Y(n_3962)
);

OAI21x1_ASAP7_75t_L g3963 ( 
.A1(n_3879),
.A2(n_3888),
.B(n_3889),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3852),
.Y(n_3964)
);

AND2x2_ASAP7_75t_L g3965 ( 
.A(n_3819),
.B(n_3777),
.Y(n_3965)
);

OR2x2_ASAP7_75t_L g3966 ( 
.A(n_3827),
.B(n_3794),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3902),
.B(n_3604),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3869),
.B(n_3612),
.Y(n_3968)
);

INVx3_ASAP7_75t_L g3969 ( 
.A(n_3834),
.Y(n_3969)
);

AND2x2_ASAP7_75t_L g3970 ( 
.A(n_3899),
.B(n_3604),
.Y(n_3970)
);

AND2x4_ASAP7_75t_L g3971 ( 
.A(n_3845),
.B(n_3799),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3839),
.B(n_3604),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3875),
.B(n_3882),
.Y(n_3973)
);

OR2x2_ASAP7_75t_L g3974 ( 
.A(n_3827),
.B(n_3773),
.Y(n_3974)
);

AOI21xp33_ASAP7_75t_L g3975 ( 
.A1(n_3909),
.A2(n_3781),
.B(n_3884),
.Y(n_3975)
);

INVxp67_ASAP7_75t_L g3976 ( 
.A(n_3892),
.Y(n_3976)
);

AOI22xp33_ASAP7_75t_L g3977 ( 
.A1(n_3917),
.A2(n_3884),
.B1(n_3913),
.B2(n_3898),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3852),
.Y(n_3978)
);

AND2x2_ASAP7_75t_L g3979 ( 
.A(n_3899),
.B(n_3900),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3900),
.B(n_3845),
.Y(n_3980)
);

NAND2x1_ASAP7_75t_L g3981 ( 
.A(n_3830),
.B(n_3828),
.Y(n_3981)
);

AO21x2_ASAP7_75t_L g3982 ( 
.A1(n_3868),
.A2(n_3885),
.B(n_3829),
.Y(n_3982)
);

INVx1_ASAP7_75t_L g3983 ( 
.A(n_3855),
.Y(n_3983)
);

HB1xp67_ASAP7_75t_L g3984 ( 
.A(n_3853),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3845),
.B(n_3863),
.Y(n_3985)
);

OR2x2_ASAP7_75t_L g3986 ( 
.A(n_3910),
.B(n_3911),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3863),
.B(n_3866),
.Y(n_3987)
);

HB1xp67_ASAP7_75t_L g3988 ( 
.A(n_3853),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3866),
.B(n_3881),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3876),
.B(n_3844),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3876),
.B(n_3844),
.Y(n_3991)
);

BUFx2_ASAP7_75t_SL g3992 ( 
.A(n_3883),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3854),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3854),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3855),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3871),
.B(n_3873),
.Y(n_3996)
);

BUFx6f_ASAP7_75t_L g3997 ( 
.A(n_3870),
.Y(n_3997)
);

HB1xp67_ASAP7_75t_L g3998 ( 
.A(n_3841),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3854),
.Y(n_3999)
);

AND2x2_ASAP7_75t_L g4000 ( 
.A(n_3871),
.B(n_3873),
.Y(n_4000)
);

INVx1_ASAP7_75t_SL g4001 ( 
.A(n_3883),
.Y(n_4001)
);

BUFx6f_ASAP7_75t_L g4002 ( 
.A(n_3837),
.Y(n_4002)
);

INVx1_ASAP7_75t_L g4003 ( 
.A(n_3857),
.Y(n_4003)
);

AND2x4_ASAP7_75t_L g4004 ( 
.A(n_3818),
.B(n_3823),
.Y(n_4004)
);

OAI33xp33_ASAP7_75t_L g4005 ( 
.A1(n_3885),
.A2(n_3893),
.A3(n_3891),
.B1(n_3895),
.B2(n_3890),
.B3(n_3896),
.Y(n_4005)
);

AND2x2_ASAP7_75t_L g4006 ( 
.A(n_3874),
.B(n_3903),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3822),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3826),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3874),
.B(n_3903),
.Y(n_4009)
);

NAND2xp5_ASAP7_75t_L g4010 ( 
.A(n_3916),
.B(n_3912),
.Y(n_4010)
);

INVx2_ASAP7_75t_L g4011 ( 
.A(n_3932),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3921),
.B(n_3830),
.Y(n_4012)
);

HB1xp67_ASAP7_75t_L g4013 ( 
.A(n_3952),
.Y(n_4013)
);

AND2x4_ASAP7_75t_SL g4014 ( 
.A(n_4002),
.B(n_3887),
.Y(n_4014)
);

INVx2_ASAP7_75t_SL g4015 ( 
.A(n_3932),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3932),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3924),
.Y(n_4017)
);

AND2x4_ASAP7_75t_SL g4018 ( 
.A(n_4002),
.B(n_3887),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3932),
.Y(n_4019)
);

AND2x4_ASAP7_75t_L g4020 ( 
.A(n_3952),
.B(n_3862),
.Y(n_4020)
);

AND2x2_ASAP7_75t_L g4021 ( 
.A(n_3936),
.B(n_3830),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3952),
.Y(n_4022)
);

BUFx2_ASAP7_75t_L g4023 ( 
.A(n_3944),
.Y(n_4023)
);

BUFx2_ASAP7_75t_L g4024 ( 
.A(n_3944),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_3936),
.B(n_3884),
.Y(n_4025)
);

NOR2x1_ASAP7_75t_L g4026 ( 
.A(n_3961),
.B(n_3884),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_3950),
.B(n_3818),
.Y(n_4027)
);

OR2x2_ASAP7_75t_L g4028 ( 
.A(n_3981),
.B(n_3893),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3969),
.Y(n_4029)
);

INVx1_ASAP7_75t_L g4030 ( 
.A(n_3981),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3950),
.B(n_3823),
.Y(n_4031)
);

HB1xp67_ASAP7_75t_L g4032 ( 
.A(n_3961),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3925),
.Y(n_4033)
);

NOR2xp33_ASAP7_75t_SL g4034 ( 
.A(n_3926),
.B(n_3837),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3950),
.B(n_3848),
.Y(n_4035)
);

HB1xp67_ASAP7_75t_L g4036 ( 
.A(n_3961),
.Y(n_4036)
);

AND2x2_ASAP7_75t_L g4037 ( 
.A(n_3980),
.B(n_3848),
.Y(n_4037)
);

AOI22xp33_ASAP7_75t_L g4038 ( 
.A1(n_3926),
.A2(n_3906),
.B1(n_3898),
.B2(n_3877),
.Y(n_4038)
);

INVx2_ASAP7_75t_L g4039 ( 
.A(n_3969),
.Y(n_4039)
);

INVx1_ASAP7_75t_L g4040 ( 
.A(n_3925),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3925),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3918),
.Y(n_4042)
);

BUFx2_ASAP7_75t_L g4043 ( 
.A(n_3938),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_3980),
.B(n_3843),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_3937),
.B(n_3843),
.Y(n_4045)
);

HB1xp67_ASAP7_75t_L g4046 ( 
.A(n_3961),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3935),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3929),
.B(n_3847),
.Y(n_4048)
);

NOR2x1_ASAP7_75t_SL g4049 ( 
.A(n_3956),
.B(n_3861),
.Y(n_4049)
);

AND2x2_ASAP7_75t_L g4050 ( 
.A(n_3954),
.B(n_3838),
.Y(n_4050)
);

AND2x2_ASAP7_75t_SL g4051 ( 
.A(n_3977),
.B(n_3887),
.Y(n_4051)
);

INVx2_ASAP7_75t_L g4052 ( 
.A(n_3969),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3982),
.B(n_3846),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3954),
.B(n_3832),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3985),
.B(n_3832),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_3969),
.Y(n_4056)
);

OR2x2_ASAP7_75t_L g4057 ( 
.A(n_3938),
.B(n_3891),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3985),
.B(n_3838),
.Y(n_4058)
);

INVx2_ASAP7_75t_L g4059 ( 
.A(n_3939),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3939),
.Y(n_4060)
);

INVx2_ASAP7_75t_L g4061 ( 
.A(n_3935),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3987),
.B(n_3828),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3935),
.Y(n_4063)
);

INVx2_ASAP7_75t_L g4064 ( 
.A(n_3943),
.Y(n_4064)
);

INVx4_ASAP7_75t_L g4065 ( 
.A(n_4014),
.Y(n_4065)
);

HB1xp67_ASAP7_75t_L g4066 ( 
.A(n_4032),
.Y(n_4066)
);

AND2x2_ASAP7_75t_L g4067 ( 
.A(n_4025),
.B(n_3923),
.Y(n_4067)
);

NOR2xp33_ASAP7_75t_L g4068 ( 
.A(n_4034),
.B(n_3941),
.Y(n_4068)
);

INVx3_ASAP7_75t_L g4069 ( 
.A(n_4014),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_4025),
.B(n_3923),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_4023),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_4032),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_L g4073 ( 
.A(n_4025),
.B(n_3946),
.Y(n_4073)
);

NOR2xp33_ASAP7_75t_SL g4074 ( 
.A(n_4034),
.B(n_4001),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_SL g4075 ( 
.A(n_4026),
.B(n_4002),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_4043),
.Y(n_4076)
);

INVx2_ASAP7_75t_SL g4077 ( 
.A(n_4036),
.Y(n_4077)
);

INVxp67_ASAP7_75t_SL g4078 ( 
.A(n_4036),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_4014),
.B(n_3923),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_4046),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_4023),
.Y(n_4081)
);

AND2x2_ASAP7_75t_L g4082 ( 
.A(n_4014),
.B(n_3992),
.Y(n_4082)
);

INVx1_ASAP7_75t_L g4083 ( 
.A(n_4023),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_4046),
.Y(n_4084)
);

AND2x4_ASAP7_75t_SL g4085 ( 
.A(n_4017),
.B(n_4002),
.Y(n_4085)
);

AND2x2_ASAP7_75t_L g4086 ( 
.A(n_4018),
.B(n_3992),
.Y(n_4086)
);

AND2x2_ASAP7_75t_L g4087 ( 
.A(n_4018),
.B(n_3946),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_4043),
.Y(n_4088)
);

OAI22xp5_ASAP7_75t_L g4089 ( 
.A1(n_4038),
.A2(n_3946),
.B1(n_3914),
.B2(n_3922),
.Y(n_4089)
);

OR2x2_ASAP7_75t_L g4090 ( 
.A(n_4012),
.B(n_3919),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_SL g4091 ( 
.A(n_4026),
.B(n_4002),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_4043),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_4012),
.B(n_3919),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_4018),
.B(n_3997),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4038),
.B(n_3989),
.Y(n_4095)
);

HB1xp67_ASAP7_75t_L g4096 ( 
.A(n_4059),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_4049),
.B(n_3989),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_4049),
.B(n_3979),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_4029),
.Y(n_4099)
);

AND2x4_ASAP7_75t_L g4100 ( 
.A(n_4018),
.B(n_3997),
.Y(n_4100)
);

OAI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_4057),
.A2(n_3962),
.B1(n_3861),
.B2(n_3934),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_4049),
.B(n_3979),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_L g4103 ( 
.A(n_4017),
.B(n_3976),
.Y(n_4103)
);

NAND2x1p5_ASAP7_75t_L g4104 ( 
.A(n_4024),
.B(n_3997),
.Y(n_4104)
);

AND2x4_ASAP7_75t_SL g4105 ( 
.A(n_4045),
.B(n_3997),
.Y(n_4105)
);

NOR2xp67_ASAP7_75t_L g4106 ( 
.A(n_4059),
.B(n_3984),
.Y(n_4106)
);

OR2x2_ASAP7_75t_L g4107 ( 
.A(n_4059),
.B(n_3947),
.Y(n_4107)
);

HB1xp67_ASAP7_75t_L g4108 ( 
.A(n_4059),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_4051),
.B(n_3997),
.Y(n_4109)
);

AND2x4_ASAP7_75t_SL g4110 ( 
.A(n_4045),
.B(n_3886),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4051),
.B(n_4006),
.Y(n_4111)
);

NAND3xp33_ASAP7_75t_L g4112 ( 
.A(n_4021),
.B(n_3975),
.C(n_3967),
.Y(n_4112)
);

AND2x2_ASAP7_75t_L g4113 ( 
.A(n_4051),
.B(n_3987),
.Y(n_4113)
);

OR2x2_ASAP7_75t_L g4114 ( 
.A(n_4060),
.B(n_3947),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4029),
.Y(n_4115)
);

INVx2_ASAP7_75t_L g4116 ( 
.A(n_4024),
.Y(n_4116)
);

OR2x2_ASAP7_75t_L g4117 ( 
.A(n_4076),
.B(n_4057),
.Y(n_4117)
);

AND2x2_ASAP7_75t_L g4118 ( 
.A(n_4067),
.B(n_4051),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4066),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4072),
.Y(n_4120)
);

OR2x2_ASAP7_75t_L g4121 ( 
.A(n_4076),
.B(n_4057),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_4067),
.B(n_3996),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_4070),
.B(n_4113),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4070),
.B(n_3996),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4078),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_4113),
.B(n_4000),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4077),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4109),
.B(n_4000),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_4109),
.B(n_4006),
.Y(n_4129)
);

HB1xp67_ASAP7_75t_L g4130 ( 
.A(n_4106),
.Y(n_4130)
);

AND2x2_ASAP7_75t_L g4131 ( 
.A(n_4110),
.B(n_4087),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_4110),
.B(n_4009),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4077),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_4104),
.Y(n_4134)
);

HB1xp67_ASAP7_75t_L g4135 ( 
.A(n_4104),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4116),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_4116),
.Y(n_4137)
);

BUFx2_ASAP7_75t_L g4138 ( 
.A(n_4104),
.Y(n_4138)
);

AND2x4_ASAP7_75t_L g4139 ( 
.A(n_4100),
.B(n_4030),
.Y(n_4139)
);

OR2x2_ASAP7_75t_L g4140 ( 
.A(n_4088),
.B(n_4060),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4071),
.Y(n_4141)
);

BUFx3_ASAP7_75t_L g4142 ( 
.A(n_4100),
.Y(n_4142)
);

OR2x2_ASAP7_75t_L g4143 ( 
.A(n_4088),
.B(n_4060),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4092),
.Y(n_4144)
);

AND2x2_ASAP7_75t_L g4145 ( 
.A(n_4087),
.B(n_4009),
.Y(n_4145)
);

OR2x2_ASAP7_75t_L g4146 ( 
.A(n_4092),
.B(n_4060),
.Y(n_4146)
);

NAND2xp5_ASAP7_75t_L g4147 ( 
.A(n_4085),
.B(n_3948),
.Y(n_4147)
);

OR2x2_ASAP7_75t_L g4148 ( 
.A(n_4096),
.B(n_4028),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_4108),
.B(n_4028),
.Y(n_4149)
);

INVx1_ASAP7_75t_SL g4150 ( 
.A(n_4082),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4082),
.B(n_4086),
.Y(n_4151)
);

AND2x2_ASAP7_75t_L g4152 ( 
.A(n_4086),
.B(n_4079),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4071),
.Y(n_4153)
);

AND2x4_ASAP7_75t_SL g4154 ( 
.A(n_4100),
.B(n_3948),
.Y(n_4154)
);

BUFx3_ASAP7_75t_L g4155 ( 
.A(n_4069),
.Y(n_4155)
);

AND2x2_ASAP7_75t_L g4156 ( 
.A(n_4123),
.B(n_4079),
.Y(n_4156)
);

NAND2xp5_ASAP7_75t_L g4157 ( 
.A(n_4123),
.B(n_4085),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4122),
.B(n_4094),
.Y(n_4158)
);

OR2x2_ASAP7_75t_L g4159 ( 
.A(n_4148),
.B(n_4090),
.Y(n_4159)
);

OR2x2_ASAP7_75t_L g4160 ( 
.A(n_4148),
.B(n_4090),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4149),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_4122),
.B(n_4094),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_4149),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4140),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_4142),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_4124),
.B(n_4105),
.Y(n_4166)
);

AND2x2_ASAP7_75t_L g4167 ( 
.A(n_4124),
.B(n_4105),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4140),
.Y(n_4168)
);

INVxp67_ASAP7_75t_L g4169 ( 
.A(n_4132),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_4142),
.Y(n_4170)
);

NAND2xp5_ASAP7_75t_L g4171 ( 
.A(n_4126),
.B(n_4068),
.Y(n_4171)
);

INVx2_ASAP7_75t_L g4172 ( 
.A(n_4142),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4143),
.Y(n_4173)
);

HB1xp67_ASAP7_75t_L g4174 ( 
.A(n_4155),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_4155),
.Y(n_4175)
);

INVx1_ASAP7_75t_SL g4176 ( 
.A(n_4132),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4126),
.B(n_4069),
.Y(n_4177)
);

NAND2xp5_ASAP7_75t_L g4178 ( 
.A(n_4118),
.B(n_4111),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_4118),
.B(n_4069),
.Y(n_4179)
);

AND2x2_ASAP7_75t_L g4180 ( 
.A(n_4145),
.B(n_4065),
.Y(n_4180)
);

OR2x2_ASAP7_75t_L g4181 ( 
.A(n_4117),
.B(n_4093),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_4156),
.B(n_4145),
.Y(n_4182)
);

AND2x2_ASAP7_75t_L g4183 ( 
.A(n_4156),
.B(n_4129),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4179),
.B(n_4129),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_4174),
.Y(n_4185)
);

INVx2_ASAP7_75t_L g4186 ( 
.A(n_4181),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4179),
.B(n_4128),
.Y(n_4187)
);

BUFx2_ASAP7_75t_L g4188 ( 
.A(n_4164),
.Y(n_4188)
);

NAND2x1_ASAP7_75t_L g4189 ( 
.A(n_4177),
.B(n_4065),
.Y(n_4189)
);

AND2x4_ASAP7_75t_L g4190 ( 
.A(n_4165),
.B(n_4155),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4164),
.Y(n_4191)
);

AND2x4_ASAP7_75t_L g4192 ( 
.A(n_4165),
.B(n_4154),
.Y(n_4192)
);

AOI22xp33_ASAP7_75t_L g4193 ( 
.A1(n_4171),
.A2(n_4005),
.B1(n_4089),
.B2(n_4112),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4181),
.Y(n_4194)
);

OR2x2_ASAP7_75t_L g4195 ( 
.A(n_4159),
.B(n_4117),
.Y(n_4195)
);

AND2x2_ASAP7_75t_L g4196 ( 
.A(n_4177),
.B(n_4128),
.Y(n_4196)
);

INVxp67_ASAP7_75t_SL g4197 ( 
.A(n_4159),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_4158),
.B(n_4152),
.Y(n_4198)
);

OR2x6_ASAP7_75t_L g4199 ( 
.A(n_4170),
.B(n_4144),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4168),
.Y(n_4200)
);

AND2x2_ASAP7_75t_L g4201 ( 
.A(n_4158),
.B(n_4152),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_4195),
.Y(n_4202)
);

AND2x2_ASAP7_75t_L g4203 ( 
.A(n_4201),
.B(n_4162),
.Y(n_4203)
);

INVx1_ASAP7_75t_SL g4204 ( 
.A(n_4195),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4199),
.Y(n_4205)
);

AND2x2_ASAP7_75t_L g4206 ( 
.A(n_4201),
.B(n_4162),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_4199),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4188),
.Y(n_4208)
);

INVxp67_ASAP7_75t_SL g4209 ( 
.A(n_4197),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4188),
.Y(n_4210)
);

INVxp67_ASAP7_75t_L g4211 ( 
.A(n_4199),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4199),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4184),
.B(n_4151),
.Y(n_4213)
);

INVx2_ASAP7_75t_L g4214 ( 
.A(n_4192),
.Y(n_4214)
);

AOI22xp5_ASAP7_75t_L g4215 ( 
.A1(n_4193),
.A2(n_4074),
.B1(n_4101),
.B2(n_4095),
.Y(n_4215)
);

HB1xp67_ASAP7_75t_L g4216 ( 
.A(n_4192),
.Y(n_4216)
);

INVx1_ASAP7_75t_L g4217 ( 
.A(n_4192),
.Y(n_4217)
);

O2A1O1Ixp33_ASAP7_75t_L g4218 ( 
.A1(n_4186),
.A2(n_4130),
.B(n_4091),
.C(n_4075),
.Y(n_4218)
);

INVx2_ASAP7_75t_L g4219 ( 
.A(n_4202),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4203),
.B(n_4184),
.Y(n_4220)
);

OR2x2_ASAP7_75t_L g4221 ( 
.A(n_4204),
.B(n_4198),
.Y(n_4221)
);

AOI22xp5_ASAP7_75t_L g4222 ( 
.A1(n_4206),
.A2(n_4182),
.B1(n_4150),
.B2(n_4102),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4216),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_4202),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_4216),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_4214),
.B(n_4182),
.Y(n_4226)
);

OR2x6_ASAP7_75t_L g4227 ( 
.A(n_4213),
.B(n_4186),
.Y(n_4227)
);

INVxp67_ASAP7_75t_L g4228 ( 
.A(n_4209),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_4217),
.B(n_4187),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4209),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4220),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4226),
.Y(n_4232)
);

NOR2xp33_ASAP7_75t_L g4233 ( 
.A(n_4222),
.B(n_4073),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4223),
.Y(n_4234)
);

INVxp67_ASAP7_75t_L g4235 ( 
.A(n_4227),
.Y(n_4235)
);

OAI322xp33_ASAP7_75t_L g4236 ( 
.A1(n_4228),
.A2(n_4215),
.A3(n_4121),
.B1(n_4160),
.B2(n_4093),
.C1(n_4125),
.C2(n_4169),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4225),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4229),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4232),
.B(n_4183),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4236),
.Y(n_4240)
);

AOI322xp5_ASAP7_75t_L g4241 ( 
.A1(n_4233),
.A2(n_4098),
.A3(n_4176),
.B1(n_4103),
.B2(n_4097),
.C1(n_4183),
.C2(n_4125),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4235),
.B(n_4187),
.Y(n_4242)
);

OR2x2_ASAP7_75t_L g4243 ( 
.A(n_4237),
.B(n_4160),
.Y(n_4243)
);

BUFx2_ASAP7_75t_L g4244 ( 
.A(n_4234),
.Y(n_4244)
);

OAI22xp5_ASAP7_75t_L g4245 ( 
.A1(n_4231),
.A2(n_4157),
.B1(n_4178),
.B2(n_4221),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4238),
.Y(n_4246)
);

AO22x1_ASAP7_75t_L g4247 ( 
.A1(n_4233),
.A2(n_4190),
.B1(n_4194),
.B2(n_4208),
.Y(n_4247)
);

OAI222xp33_ASAP7_75t_L g4248 ( 
.A1(n_4235),
.A2(n_4189),
.B1(n_4065),
.B2(n_4227),
.C1(n_4121),
.C2(n_4194),
.Y(n_4248)
);

AOI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4233),
.A2(n_4196),
.B1(n_4151),
.B2(n_4167),
.Y(n_4249)
);

AND2x2_ASAP7_75t_L g4250 ( 
.A(n_4232),
.B(n_4196),
.Y(n_4250)
);

NOR2xp33_ASAP7_75t_L g4251 ( 
.A(n_4236),
.B(n_4131),
.Y(n_4251)
);

AOI22xp5_ASAP7_75t_L g4252 ( 
.A1(n_4251),
.A2(n_4166),
.B1(n_4167),
.B2(n_4131),
.Y(n_4252)
);

OR2x2_ASAP7_75t_L g4253 ( 
.A(n_4243),
.B(n_4170),
.Y(n_4253)
);

AOI32xp33_ASAP7_75t_L g4254 ( 
.A1(n_4239),
.A2(n_4180),
.A3(n_4166),
.B1(n_4154),
.B2(n_4161),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4249),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_4250),
.Y(n_4256)
);

OR2x2_ASAP7_75t_L g4257 ( 
.A(n_4247),
.B(n_4172),
.Y(n_4257)
);

AOI21xp33_ASAP7_75t_L g4258 ( 
.A1(n_4242),
.A2(n_4218),
.B(n_4163),
.Y(n_4258)
);

OAI22xp5_ASAP7_75t_L g4259 ( 
.A1(n_4240),
.A2(n_4147),
.B1(n_4172),
.B2(n_4185),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_4241),
.B(n_4190),
.Y(n_4260)
);

OR2x2_ASAP7_75t_L g4261 ( 
.A(n_4245),
.B(n_4161),
.Y(n_4261)
);

INVx1_ASAP7_75t_L g4262 ( 
.A(n_4244),
.Y(n_4262)
);

OAI211xp5_ASAP7_75t_SL g4263 ( 
.A1(n_4246),
.A2(n_4230),
.B(n_4219),
.C(n_4224),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4248),
.Y(n_4264)
);

AOI32xp33_ASAP7_75t_SL g4265 ( 
.A1(n_4251),
.A2(n_4127),
.A3(n_4133),
.B1(n_4120),
.B2(n_4119),
.Y(n_4265)
);

HB1xp67_ASAP7_75t_L g4266 ( 
.A(n_4243),
.Y(n_4266)
);

AND2x2_ASAP7_75t_L g4267 ( 
.A(n_4250),
.B(n_4180),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4249),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_4241),
.B(n_4190),
.Y(n_4269)
);

OAI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_4249),
.A2(n_4163),
.B(n_4210),
.Y(n_4270)
);

AND2x4_ASAP7_75t_SL g4271 ( 
.A(n_4239),
.B(n_4175),
.Y(n_4271)
);

O2A1O1Ixp33_ASAP7_75t_SL g4272 ( 
.A1(n_4248),
.A2(n_4168),
.B(n_4173),
.C(n_4211),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_4241),
.B(n_4175),
.Y(n_4273)
);

AOI221xp5_ASAP7_75t_L g4274 ( 
.A1(n_4258),
.A2(n_4127),
.B1(n_4133),
.B2(n_4119),
.C(n_4120),
.Y(n_4274)
);

OAI221xp5_ASAP7_75t_L g4275 ( 
.A1(n_4254),
.A2(n_4173),
.B1(n_4135),
.B2(n_4138),
.C(n_4211),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_L g4276 ( 
.A(n_4267),
.B(n_4154),
.Y(n_4276)
);

AOI21xp33_ASAP7_75t_L g4277 ( 
.A1(n_4266),
.A2(n_4253),
.B(n_4261),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_4272),
.A2(n_4212),
.B(n_4205),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4271),
.B(n_4144),
.Y(n_4279)
);

NAND2x1p5_ASAP7_75t_L g4280 ( 
.A(n_4257),
.B(n_4207),
.Y(n_4280)
);

AOI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_4270),
.A2(n_4205),
.B(n_4200),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_4260),
.A2(n_4191),
.B(n_4134),
.Y(n_4282)
);

AND2x2_ASAP7_75t_L g4283 ( 
.A(n_4252),
.B(n_4144),
.Y(n_4283)
);

OAI211xp5_ASAP7_75t_SL g4284 ( 
.A1(n_4255),
.A2(n_4136),
.B(n_4137),
.C(n_4143),
.Y(n_4284)
);

OAI211xp5_ASAP7_75t_L g4285 ( 
.A1(n_4269),
.A2(n_4138),
.B(n_4136),
.C(n_4137),
.Y(n_4285)
);

AOI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4259),
.A2(n_4139),
.B1(n_4080),
.B2(n_4084),
.Y(n_4286)
);

INVx1_ASAP7_75t_L g4287 ( 
.A(n_4273),
.Y(n_4287)
);

AOI21xp5_ASAP7_75t_L g4288 ( 
.A1(n_4262),
.A2(n_4134),
.B(n_4146),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_4256),
.Y(n_4289)
);

O2A1O1Ixp33_ASAP7_75t_L g4290 ( 
.A1(n_4263),
.A2(n_4146),
.B(n_4153),
.C(n_4141),
.Y(n_4290)
);

NOR3xp33_ASAP7_75t_L g4291 ( 
.A(n_4268),
.B(n_4141),
.C(n_4153),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_4264),
.Y(n_4292)
);

OAI21xp33_ASAP7_75t_L g4293 ( 
.A1(n_4265),
.A2(n_4114),
.B(n_4107),
.Y(n_4293)
);

AOI221xp5_ASAP7_75t_L g4294 ( 
.A1(n_4258),
.A2(n_4139),
.B1(n_4134),
.B2(n_4081),
.C(n_4083),
.Y(n_4294)
);

AOI221xp5_ASAP7_75t_L g4295 ( 
.A1(n_4258),
.A2(n_4139),
.B1(n_4081),
.B2(n_4083),
.C(n_4030),
.Y(n_4295)
);

OAI221xp5_ASAP7_75t_L g4296 ( 
.A1(n_4254),
.A2(n_4114),
.B1(n_4107),
.B2(n_4030),
.C(n_4115),
.Y(n_4296)
);

AOI22xp5_ASAP7_75t_L g4297 ( 
.A1(n_4252),
.A2(n_4139),
.B1(n_4099),
.B2(n_4021),
.Y(n_4297)
);

AOI211xp5_ASAP7_75t_L g4298 ( 
.A1(n_4258),
.A2(n_4021),
.B(n_4048),
.C(n_4013),
.Y(n_4298)
);

OAI22xp33_ASAP7_75t_L g4299 ( 
.A1(n_4252),
.A2(n_4028),
.B1(n_4024),
.B2(n_4015),
.Y(n_4299)
);

O2A1O1Ixp5_ASAP7_75t_L g4300 ( 
.A1(n_4285),
.A2(n_4022),
.B(n_4039),
.C(n_4029),
.Y(n_4300)
);

AND2x2_ASAP7_75t_L g4301 ( 
.A(n_4283),
.B(n_4048),
.Y(n_4301)
);

AOI211xp5_ASAP7_75t_SL g4302 ( 
.A1(n_4277),
.A2(n_4013),
.B(n_4042),
.C(n_4016),
.Y(n_4302)
);

AOI211xp5_ASAP7_75t_L g4303 ( 
.A1(n_4275),
.A2(n_4053),
.B(n_4042),
.C(n_4016),
.Y(n_4303)
);

OAI21xp33_ASAP7_75t_L g4304 ( 
.A1(n_4276),
.A2(n_4045),
.B(n_4015),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_4288),
.A2(n_4053),
.B(n_4022),
.Y(n_4305)
);

NAND3xp33_ASAP7_75t_L g4306 ( 
.A(n_4274),
.B(n_4022),
.C(n_4016),
.Y(n_4306)
);

OAI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_4297),
.A2(n_4010),
.B1(n_3986),
.B2(n_3973),
.Y(n_4307)
);

NOR3x1_ASAP7_75t_L g4308 ( 
.A(n_4296),
.B(n_4015),
.C(n_4041),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_4294),
.B(n_3894),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4278),
.A2(n_4022),
.B(n_4011),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_SL g4311 ( 
.A(n_4298),
.B(n_4029),
.Y(n_4311)
);

AOI211xp5_ASAP7_75t_L g4312 ( 
.A1(n_4299),
.A2(n_4035),
.B(n_4031),
.C(n_4027),
.Y(n_4312)
);

AOI222xp33_ASAP7_75t_L g4313 ( 
.A1(n_4293),
.A2(n_4019),
.B1(n_4011),
.B2(n_4047),
.C1(n_4041),
.C2(n_4040),
.Y(n_4313)
);

NAND2xp5_ASAP7_75t_L g4314 ( 
.A(n_4286),
.B(n_3933),
.Y(n_4314)
);

OAI22xp5_ASAP7_75t_L g4315 ( 
.A1(n_4292),
.A2(n_3986),
.B1(n_3933),
.B2(n_3940),
.Y(n_4315)
);

AOI322xp5_ASAP7_75t_L g4316 ( 
.A1(n_4287),
.A2(n_4035),
.A3(n_4027),
.B1(n_4031),
.B2(n_4019),
.C1(n_4011),
.C2(n_4052),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_4295),
.B(n_4039),
.Y(n_4317)
);

OAI22xp5_ASAP7_75t_L g4318 ( 
.A1(n_4289),
.A2(n_3940),
.B1(n_4052),
.B2(n_4039),
.Y(n_4318)
);

O2A1O1Ixp33_ASAP7_75t_L g4319 ( 
.A1(n_4290),
.A2(n_4019),
.B(n_4011),
.C(n_3982),
.Y(n_4319)
);

NAND4xp25_ASAP7_75t_SL g4320 ( 
.A(n_4282),
.B(n_4033),
.C(n_4040),
.D(n_4041),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4291),
.B(n_3982),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_4281),
.A2(n_4019),
.B(n_4039),
.Y(n_4322)
);

AOI211x1_ASAP7_75t_SL g4323 ( 
.A1(n_4284),
.A2(n_4052),
.B(n_4056),
.C(n_4061),
.Y(n_4323)
);

NOR2xp67_ASAP7_75t_L g4324 ( 
.A(n_4320),
.B(n_4279),
.Y(n_4324)
);

NOR3x1_ASAP7_75t_L g4325 ( 
.A(n_4309),
.B(n_4280),
.C(n_4040),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4318),
.Y(n_4326)
);

NAND4xp25_ASAP7_75t_SL g4327 ( 
.A(n_4312),
.B(n_4303),
.C(n_4316),
.D(n_4313),
.Y(n_4327)
);

AOI221xp5_ASAP7_75t_L g4328 ( 
.A1(n_4315),
.A2(n_4033),
.B1(n_4047),
.B2(n_4052),
.C(n_4056),
.Y(n_4328)
);

NAND4xp75_ASAP7_75t_L g4329 ( 
.A(n_4308),
.B(n_4317),
.C(n_4310),
.D(n_4311),
.Y(n_4329)
);

OAI221xp5_ASAP7_75t_L g4330 ( 
.A1(n_4304),
.A2(n_4056),
.B1(n_4033),
.B2(n_4047),
.C(n_4064),
.Y(n_4330)
);

NOR4xp25_ASAP7_75t_L g4331 ( 
.A(n_4306),
.B(n_4321),
.C(n_4319),
.D(n_4314),
.Y(n_4331)
);

A2O1A1Ixp33_ASAP7_75t_L g4332 ( 
.A1(n_4300),
.A2(n_4056),
.B(n_4020),
.C(n_4061),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4301),
.Y(n_4333)
);

A2O1A1Ixp33_ASAP7_75t_L g4334 ( 
.A1(n_4302),
.A2(n_4020),
.B(n_4063),
.C(n_4061),
.Y(n_4334)
);

BUFx6f_ASAP7_75t_SL g4335 ( 
.A(n_4323),
.Y(n_4335)
);

AOI32xp33_ASAP7_75t_L g4336 ( 
.A1(n_4307),
.A2(n_4035),
.A3(n_4031),
.B1(n_4027),
.B2(n_4020),
.Y(n_4336)
);

AOI22xp33_ASAP7_75t_L g4337 ( 
.A1(n_4322),
.A2(n_4020),
.B1(n_4044),
.B2(n_4037),
.Y(n_4337)
);

A2O1A1Ixp33_ASAP7_75t_L g4338 ( 
.A1(n_4305),
.A2(n_4020),
.B(n_4063),
.C(n_4061),
.Y(n_4338)
);

AOI222xp33_ASAP7_75t_L g4339 ( 
.A1(n_4304),
.A2(n_4064),
.B1(n_4063),
.B2(n_4020),
.C1(n_3999),
.C2(n_3994),
.Y(n_4339)
);

NOR3xp33_ASAP7_75t_SL g4340 ( 
.A(n_4304),
.B(n_3972),
.C(n_3928),
.Y(n_4340)
);

NOR2xp33_ASAP7_75t_L g4341 ( 
.A(n_4333),
.B(n_4063),
.Y(n_4341)
);

NAND3xp33_ASAP7_75t_L g4342 ( 
.A(n_4326),
.B(n_4064),
.C(n_3931),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_4337),
.B(n_3918),
.Y(n_4343)
);

NOR3xp33_ASAP7_75t_L g4344 ( 
.A(n_4327),
.B(n_4064),
.C(n_3920),
.Y(n_4344)
);

INVx3_ASAP7_75t_L g4345 ( 
.A(n_4329),
.Y(n_4345)
);

NOR3xp33_ASAP7_75t_L g4346 ( 
.A(n_4324),
.B(n_3931),
.C(n_3928),
.Y(n_4346)
);

AOI211xp5_ASAP7_75t_SL g4347 ( 
.A1(n_4330),
.A2(n_3998),
.B(n_4062),
.C(n_4037),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_4340),
.B(n_4336),
.Y(n_4348)
);

NAND2xp5_ASAP7_75t_SL g4349 ( 
.A(n_4328),
.B(n_3920),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_L g4350 ( 
.A(n_4334),
.B(n_4325),
.Y(n_4350)
);

AOI22xp33_ASAP7_75t_L g4351 ( 
.A1(n_4335),
.A2(n_4037),
.B1(n_4044),
.B2(n_4055),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4332),
.B(n_4007),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4335),
.Y(n_4353)
);

AOI21xp5_ASAP7_75t_L g4354 ( 
.A1(n_4331),
.A2(n_3994),
.B(n_3999),
.Y(n_4354)
);

NAND2xp5_ASAP7_75t_L g4355 ( 
.A(n_4338),
.B(n_4007),
.Y(n_4355)
);

NOR4xp25_ASAP7_75t_L g4356 ( 
.A(n_4353),
.B(n_4339),
.C(n_3943),
.D(n_3993),
.Y(n_4356)
);

NOR2x1_ASAP7_75t_L g4357 ( 
.A(n_4350),
.B(n_4341),
.Y(n_4357)
);

AOI221xp5_ASAP7_75t_SL g4358 ( 
.A1(n_4354),
.A2(n_3993),
.B1(n_3943),
.B2(n_4062),
.C(n_3953),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_4347),
.B(n_4008),
.Y(n_4359)
);

NAND4xp25_ASAP7_75t_L g4360 ( 
.A(n_4344),
.B(n_4044),
.C(n_4062),
.D(n_4055),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_4351),
.B(n_4008),
.Y(n_4361)
);

O2A1O1Ixp33_ASAP7_75t_L g4362 ( 
.A1(n_4348),
.A2(n_3988),
.B(n_3957),
.C(n_3953),
.Y(n_4362)
);

AND2x2_ASAP7_75t_L g4363 ( 
.A(n_4345),
.B(n_4055),
.Y(n_4363)
);

NOR2x1_ASAP7_75t_L g4364 ( 
.A(n_4345),
.B(n_3949),
.Y(n_4364)
);

AND4x1_ASAP7_75t_L g4365 ( 
.A(n_4342),
.B(n_4058),
.C(n_4054),
.D(n_4050),
.Y(n_4365)
);

NOR4xp25_ASAP7_75t_L g4366 ( 
.A(n_4349),
.B(n_3957),
.C(n_3953),
.D(n_4058),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_4346),
.B(n_4003),
.Y(n_4367)
);

INVx2_ASAP7_75t_SL g4368 ( 
.A(n_4343),
.Y(n_4368)
);

AND2x4_ASAP7_75t_L g4369 ( 
.A(n_4355),
.B(n_3960),
.Y(n_4369)
);

AOI211xp5_ASAP7_75t_L g4370 ( 
.A1(n_4352),
.A2(n_4058),
.B(n_4050),
.C(n_4054),
.Y(n_4370)
);

AOI221x1_ASAP7_75t_L g4371 ( 
.A1(n_4353),
.A2(n_3957),
.B1(n_4054),
.B2(n_4050),
.C(n_3960),
.Y(n_4371)
);

NOR2x1_ASAP7_75t_L g4372 ( 
.A(n_4353),
.B(n_3964),
.Y(n_4372)
);

NOR2x1_ASAP7_75t_L g4373 ( 
.A(n_4353),
.B(n_3964),
.Y(n_4373)
);

CKINVDCx20_ASAP7_75t_R g4374 ( 
.A(n_4363),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4369),
.Y(n_4375)
);

NOR2x1_ASAP7_75t_L g4376 ( 
.A(n_4364),
.B(n_3995),
.Y(n_4376)
);

INVx1_ASAP7_75t_L g4377 ( 
.A(n_4372),
.Y(n_4377)
);

HB1xp67_ASAP7_75t_L g4378 ( 
.A(n_4373),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4362),
.Y(n_4379)
);

NOR2x1_ASAP7_75t_L g4380 ( 
.A(n_4357),
.B(n_3995),
.Y(n_4380)
);

HB1xp67_ASAP7_75t_L g4381 ( 
.A(n_4359),
.Y(n_4381)
);

AND2x4_ASAP7_75t_L g4382 ( 
.A(n_4369),
.B(n_4003),
.Y(n_4382)
);

AND2x2_ASAP7_75t_L g4383 ( 
.A(n_4370),
.B(n_3990),
.Y(n_4383)
);

INVxp67_ASAP7_75t_SL g4384 ( 
.A(n_4361),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4367),
.Y(n_4385)
);

OR2x2_ASAP7_75t_L g4386 ( 
.A(n_4360),
.B(n_4366),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4368),
.Y(n_4387)
);

NOR2xp67_ASAP7_75t_L g4388 ( 
.A(n_4356),
.B(n_3958),
.Y(n_4388)
);

INVx1_ASAP7_75t_SL g4389 ( 
.A(n_4365),
.Y(n_4389)
);

AOI22xp5_ASAP7_75t_L g4390 ( 
.A1(n_4358),
.A2(n_3991),
.B1(n_3990),
.B2(n_3983),
.Y(n_4390)
);

AND4x1_ASAP7_75t_L g4391 ( 
.A(n_4387),
.B(n_4371),
.C(n_3991),
.D(n_3965),
.Y(n_4391)
);

NOR2xp33_ASAP7_75t_L g4392 ( 
.A(n_4389),
.B(n_3978),
.Y(n_4392)
);

NOR2x1p5_ASAP7_75t_L g4393 ( 
.A(n_4384),
.B(n_3949),
.Y(n_4393)
);

NOR3xp33_ASAP7_75t_L g4394 ( 
.A(n_4379),
.B(n_3963),
.C(n_3983),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4376),
.Y(n_4395)
);

NAND4xp75_ASAP7_75t_L g4396 ( 
.A(n_4380),
.B(n_3927),
.C(n_3978),
.D(n_3958),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4383),
.Y(n_4397)
);

OAI211xp5_ASAP7_75t_SL g4398 ( 
.A1(n_4386),
.A2(n_3959),
.B(n_3951),
.C(n_3974),
.Y(n_4398)
);

NOR2x1p5_ASAP7_75t_L g4399 ( 
.A(n_4375),
.B(n_3974),
.Y(n_4399)
);

NOR4xp25_ASAP7_75t_L g4400 ( 
.A(n_4377),
.B(n_3927),
.C(n_3970),
.D(n_3951),
.Y(n_4400)
);

NAND4xp25_ASAP7_75t_L g4401 ( 
.A(n_4388),
.B(n_4385),
.C(n_4390),
.D(n_4382),
.Y(n_4401)
);

NAND3xp33_ASAP7_75t_L g4402 ( 
.A(n_4392),
.B(n_4378),
.C(n_4381),
.Y(n_4402)
);

NOR4xp75_ASAP7_75t_L g4403 ( 
.A(n_4396),
.B(n_4374),
.C(n_3970),
.D(n_3965),
.Y(n_4403)
);

OAI211xp5_ASAP7_75t_SL g4404 ( 
.A1(n_4397),
.A2(n_3959),
.B(n_3966),
.C(n_3915),
.Y(n_4404)
);

AOI322xp5_ASAP7_75t_L g4405 ( 
.A1(n_4395),
.A2(n_4004),
.A3(n_3971),
.B1(n_3968),
.B2(n_3877),
.C1(n_3930),
.C2(n_3867),
.Y(n_4405)
);

NOR2x1_ASAP7_75t_L g4406 ( 
.A(n_4401),
.B(n_3971),
.Y(n_4406)
);

NOR2x1_ASAP7_75t_L g4407 ( 
.A(n_4393),
.B(n_4399),
.Y(n_4407)
);

AND4x2_ASAP7_75t_L g4408 ( 
.A(n_4406),
.B(n_4391),
.C(n_4398),
.D(n_4400),
.Y(n_4408)
);

NAND2x1_ASAP7_75t_L g4409 ( 
.A(n_4407),
.B(n_4394),
.Y(n_4409)
);

NOR3xp33_ASAP7_75t_L g4410 ( 
.A(n_4402),
.B(n_3963),
.C(n_3880),
.Y(n_4410)
);

OAI22xp33_ASAP7_75t_L g4411 ( 
.A1(n_4409),
.A2(n_4403),
.B1(n_4404),
.B2(n_4405),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4408),
.Y(n_4412)
);

OAI211xp5_ASAP7_75t_L g4413 ( 
.A1(n_4412),
.A2(n_4410),
.B(n_3945),
.C(n_3828),
.Y(n_4413)
);

AOI22x1_ASAP7_75t_L g4414 ( 
.A1(n_4413),
.A2(n_4411),
.B1(n_3955),
.B2(n_4004),
.Y(n_4414)
);

OAI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_4414),
.A2(n_4004),
.B1(n_3966),
.B2(n_3968),
.Y(n_4415)
);

OAI21x1_ASAP7_75t_L g4416 ( 
.A1(n_4415),
.A2(n_3930),
.B(n_3888),
.Y(n_4416)
);

OAI21xp33_ASAP7_75t_L g4417 ( 
.A1(n_4416),
.A2(n_4004),
.B(n_3971),
.Y(n_4417)
);

INVx1_ASAP7_75t_L g4418 ( 
.A(n_4417),
.Y(n_4418)
);

XNOR2xp5_ASAP7_75t_L g4419 ( 
.A(n_4418),
.B(n_3945),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4419),
.Y(n_4420)
);

NOR2xp33_ASAP7_75t_L g4421 ( 
.A(n_4420),
.B(n_3897),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4421),
.Y(n_4422)
);

OAI21x1_ASAP7_75t_L g4423 ( 
.A1(n_4422),
.A2(n_3888),
.B(n_3942),
.Y(n_4423)
);

AOI221xp5_ASAP7_75t_L g4424 ( 
.A1(n_4423),
.A2(n_3862),
.B1(n_3831),
.B2(n_3850),
.C(n_3851),
.Y(n_4424)
);

AOI21xp33_ASAP7_75t_L g4425 ( 
.A1(n_4424),
.A2(n_3945),
.B(n_3908),
.Y(n_4425)
);

AOI211xp5_ASAP7_75t_L g4426 ( 
.A1(n_4425),
.A2(n_3905),
.B(n_3904),
.C(n_3907),
.Y(n_4426)
);


endmodule