module real_jpeg_1423_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_1),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_2),
.A2(n_20),
.B1(n_21),
.B2(n_37),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_37),
.B1(n_55),
.B2(n_57),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_37),
.B1(n_44),
.B2(n_45),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_3),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_34),
.B1(n_55),
.B2(n_57),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_3),
.B(n_26),
.C(n_30),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_28),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_3),
.B(n_41),
.C(n_45),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_3),
.B(n_100),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_3),
.B(n_53),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_3),
.B(n_54),
.C(n_57),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_3),
.B(n_47),
.Y(n_237)
);

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_6),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_6),
.A2(n_24),
.B1(n_44),
.B2(n_45),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_6),
.A2(n_24),
.B1(n_55),
.B2(n_57),
.Y(n_162)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_10),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_49),
.B1(n_55),
.B2(n_57),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_85),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_83),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_69),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_15),
.B(n_69),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_62),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_35),
.C(n_50),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_17),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_17),
.A2(n_71),
.B1(n_106),
.B2(n_108),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_17),
.A2(n_71),
.B1(n_146),
.B2(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_17),
.B(n_146),
.C(n_156),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B1(n_28),
.B2(n_33),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_19),
.A2(n_64),
.B(n_66),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_26),
.Y(n_27)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_21),
.B(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_25),
.B(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_25),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_30),
.B(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_33),
.B(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_35),
.A2(n_50),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_35),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_35)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_38),
.A2(n_47),
.B1(n_107),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_39),
.B(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_39),
.A2(n_43),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

AOI22x1_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_45),
.B1(n_54),
.B2(n_58),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_45),
.B(n_230),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g106 ( 
.A1(n_47),
.A2(n_81),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_76),
.C(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_50),
.A2(n_75),
.B1(n_78),
.B2(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_59),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_52),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_52),
.A2(n_59),
.B1(n_95),
.B2(n_96),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_52),
.A2(n_59),
.B(n_96),
.Y(n_172)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_53),
.A2(n_61),
.B1(n_118),
.B2(n_145),
.Y(n_144)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_57),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_64),
.B(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.C(n_77),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_70),
.A2(n_76),
.B1(n_129),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_70),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_71),
.B(n_91),
.C(n_106),
.Y(n_149)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_76),
.A2(n_129),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_76),
.A2(n_128),
.B1(n_129),
.B2(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_76),
.A2(n_129),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_77),
.B(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_78),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_260),
.B(n_277),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_150),
.B(n_259),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_130),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_89),
.B(n_130),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_109),
.C(n_120),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_90),
.B(n_109),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_104),
.B2(n_105),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_93),
.A2(n_94),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_93),
.A2(n_94),
.B1(n_210),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_94),
.B(n_205),
.C(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_94),
.B(n_161),
.C(n_237),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_100),
.B1(n_125),
.B2(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_102),
.B(n_124),
.Y(n_123)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_102),
.A2(n_124),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_129),
.C(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_106),
.A2(n_108),
.B1(n_172),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_106),
.A2(n_108),
.B1(n_126),
.B2(n_127),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_106),
.B(n_126),
.C(n_245),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_113),
.B1(n_114),
.B2(n_119),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_114),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_119),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_112),
.B(n_125),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_119),
.A2(n_134),
.B(n_141),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_120),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_128),
.C(n_129),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_121),
.A2(n_122),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_123),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_126),
.A2(n_127),
.B1(n_229),
.B2(n_231),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_126),
.B(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_149),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_142),
.B2(n_143),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_133),
.B(n_142),
.C(n_149),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B(n_148),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_146),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_180),
.C(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_164),
.B1(n_206),
.B2(n_209),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_148),
.A2(n_264),
.B1(n_265),
.B2(n_269),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_148),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_254),
.B(n_258),
.Y(n_150)
);

OAI211xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_183),
.B(n_197),
.C(n_198),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_173),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_165),
.B2(n_166),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_168),
.C(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_163),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_158),
.B1(n_160),
.B2(n_161),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_160),
.A2(n_161),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_161),
.B(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_225),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_178),
.C(n_179),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_179),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_181),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_199),
.C(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_186),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_187),
.B(n_189),
.C(n_195),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_216),
.B(n_253),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_202),
.B(n_204),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_210),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_247),
.B(n_252),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_241),
.B(n_246),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_233),
.B(n_240),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B(n_232),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_224),
.B(n_226),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_239),
.Y(n_240)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_243),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_256),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_272),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_271),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_271),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_269),
.C(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_276),
.Y(n_279)
);


endmodule