module fake_netlist_1_5451_n_570 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_570);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_570;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_476;
wire n_384;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_77), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
INVxp67_ASAP7_75t_L g82 ( .A(n_40), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_9), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_33), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
BUFx10_ASAP7_75t_L g86 ( .A(n_67), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_50), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_5), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_27), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_49), .Y(n_91) );
BUFx5_ASAP7_75t_L g92 ( .A(n_37), .Y(n_92) );
OR2x2_ASAP7_75t_L g93 ( .A(n_9), .B(n_79), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_16), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_15), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_5), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_25), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_19), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_47), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_60), .Y(n_101) );
CKINVDCx14_ASAP7_75t_R g102 ( .A(n_13), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_56), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_3), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_38), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_57), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_20), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_36), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_18), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_39), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_59), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_51), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_3), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_70), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_55), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_28), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_86), .Y(n_120) );
BUFx3_ASAP7_75t_L g121 ( .A(n_92), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_102), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_122) );
NOR2xp33_ASAP7_75t_L g123 ( .A(n_80), .B(n_0), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_102), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_90), .B(n_2), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_92), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_97), .B(n_4), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
XOR2xp5_ASAP7_75t_L g136 ( .A(n_114), .B(n_6), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_113), .B(n_6), .Y(n_137) );
NOR2x1_ASAP7_75t_L g138 ( .A(n_85), .B(n_7), .Y(n_138) );
XOR2xp5_ASAP7_75t_L g139 ( .A(n_114), .B(n_7), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_99), .Y(n_140) );
OAI22xp5_ASAP7_75t_SL g141 ( .A1(n_88), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_87), .Y(n_142) );
INVx2_ASAP7_75t_SL g143 ( .A(n_120), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_120), .B(n_109), .Y(n_144) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_126), .A2(n_104), .B1(n_109), .B2(n_116), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_120), .B(n_82), .Y(n_146) );
BUFx10_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
BUFx10_ASAP7_75t_L g148 ( .A(n_133), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_132), .Y(n_149) );
NAND2xp33_ASAP7_75t_L g150 ( .A(n_135), .B(n_92), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_119), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_119), .Y(n_152) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_134), .A2(n_93), .B1(n_117), .B2(n_115), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_120), .A2(n_118), .B1(n_94), .B2(n_100), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_134), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_135), .A2(n_105), .B1(n_107), .B2(n_91), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx4_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
BUFx4f_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_125), .B(n_103), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_132), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_119), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_136), .Y(n_166) );
INVx1_ASAP7_75t_SL g167 ( .A(n_125), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_125), .B(n_101), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_147), .B(n_129), .Y(n_171) );
NAND2xp33_ASAP7_75t_L g172 ( .A(n_167), .B(n_92), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_147), .B(n_129), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_147), .B(n_129), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g175 ( .A1(n_155), .A2(n_148), .B1(n_163), .B2(n_149), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_148), .B(n_129), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_148), .A2(n_142), .B1(n_121), .B2(n_123), .Y(n_177) );
OAI22xp33_ASAP7_75t_L g178 ( .A1(n_145), .A2(n_122), .B1(n_127), .B2(n_137), .Y(n_178) );
NAND2xp33_ASAP7_75t_L g179 ( .A(n_143), .B(n_92), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_144), .B(n_142), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_162), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_166), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_169), .B(n_121), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_153), .A2(n_141), .B1(n_138), .B2(n_131), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_154), .A2(n_138), .B1(n_131), .B2(n_128), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_146), .B(n_128), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_162), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_143), .B(n_131), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_160), .B(n_130), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_159), .B(n_130), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_163), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_159), .B(n_108), .Y(n_192) );
BUFx4f_ASAP7_75t_SL g193 ( .A(n_166), .Y(n_193) );
INVx1_ASAP7_75t_SL g194 ( .A(n_162), .Y(n_194) );
NAND3xp33_ASAP7_75t_L g195 ( .A(n_156), .B(n_106), .C(n_95), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_159), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
NOR2xp67_ASAP7_75t_SL g198 ( .A(n_158), .B(n_111), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_158), .B(n_112), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_158), .B(n_110), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_161), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_150), .B(n_98), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_165), .B(n_96), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_165), .B(n_139), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_204), .B(n_136), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_180), .A2(n_139), .B1(n_124), .B2(n_140), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_178), .A2(n_92), .B1(n_124), .B2(n_140), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_175), .B(n_140), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_171), .B(n_124), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_170), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_170), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_191), .Y(n_212) );
OAI21xp33_ASAP7_75t_L g213 ( .A1(n_177), .A2(n_124), .B(n_140), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_124), .B1(n_140), .B2(n_168), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_191), .Y(n_215) );
OA22x2_ASAP7_75t_L g216 ( .A1(n_185), .A2(n_182), .B1(n_197), .B2(n_194), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_189), .B(n_140), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_SL g218 ( .A1(n_198), .A2(n_164), .B(n_157), .C(n_152), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_204), .B(n_8), .Y(n_219) );
OR2x6_ASAP7_75t_SL g220 ( .A(n_182), .B(n_10), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_195), .B(n_11), .Y(n_221) );
CKINVDCx8_ASAP7_75t_R g222 ( .A(n_193), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_173), .B(n_12), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_174), .B(n_161), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_176), .B(n_161), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_186), .A2(n_168), .B1(n_164), .B2(n_157), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_181), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_181), .B(n_152), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_187), .A2(n_151), .B1(n_161), .B2(n_12), .Y(n_231) );
INVx3_ASAP7_75t_SL g232 ( .A(n_181), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_200), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_199), .B(n_13), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_196), .B(n_151), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_201), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_196), .A2(n_161), .B1(n_17), .B2(n_21), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_202), .B(n_14), .Y(n_238) );
OR2x6_ASAP7_75t_L g239 ( .A(n_196), .B(n_22), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_210), .Y(n_240) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_213), .A2(n_183), .B(n_203), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_235), .A2(n_179), .B(n_172), .Y(n_242) );
AND2x4_ASAP7_75t_L g243 ( .A(n_225), .B(n_233), .Y(n_243) );
AO31x2_ASAP7_75t_L g244 ( .A1(n_237), .A2(n_201), .A3(n_192), .B(n_179), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_212), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_205), .B(n_198), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_237), .A2(n_172), .B(n_201), .Y(n_247) );
AO31x2_ASAP7_75t_L g248 ( .A1(n_231), .A2(n_78), .A3(n_24), .B(n_26), .Y(n_248) );
NAND2xp33_ASAP7_75t_SL g249 ( .A(n_206), .B(n_23), .Y(n_249) );
AOI221x1_ASAP7_75t_L g250 ( .A1(n_231), .A2(n_29), .B1(n_31), .B2(n_32), .C(n_34), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_227), .B(n_35), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_208), .A2(n_41), .B(n_42), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g253 ( .A1(n_234), .A2(n_43), .B(n_44), .C(n_46), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_217), .A2(n_48), .B(n_52), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_239), .B(n_53), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_215), .B(n_54), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_207), .A2(n_61), .B(n_62), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_230), .A2(n_63), .B(n_64), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_219), .B(n_65), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_230), .A2(n_66), .B(n_68), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_224), .A2(n_69), .B(n_71), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_73), .B(n_74), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_236), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_206), .B(n_75), .Y(n_265) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_214), .A2(n_76), .B(n_228), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_232), .B(n_211), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_209), .A2(n_218), .B(n_228), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_240), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_243), .Y(n_270) );
AO31x2_ASAP7_75t_L g271 ( .A1(n_250), .A2(n_238), .A3(n_223), .B(n_229), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_265), .A2(n_221), .B(n_216), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_243), .B(n_216), .Y(n_273) );
AOI21x1_ASAP7_75t_L g274 ( .A1(n_241), .A2(n_239), .B(n_221), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
NOR2x1_ASAP7_75t_SL g276 ( .A(n_262), .B(n_239), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_243), .B(n_220), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_240), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_264), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_245), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_245), .Y(n_281) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_268), .A2(n_236), .B(n_222), .Y(n_282) );
AOI21x1_ASAP7_75t_L g283 ( .A1(n_241), .A2(n_236), .B(n_266), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_255), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_242), .A2(n_241), .B(n_249), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_256), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_246), .B(n_267), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_256), .B(n_264), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_259), .B(n_251), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_247), .B(n_244), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_292), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_287), .A2(n_257), .B(n_252), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_292), .Y(n_295) );
BUFx12f_ASAP7_75t_L g296 ( .A(n_270), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_269), .B(n_248), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_269), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_285), .B(n_249), .Y(n_299) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_289), .A2(n_253), .B1(n_260), .B2(n_258), .C(n_261), .Y(n_300) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_283), .A2(n_252), .B(n_254), .Y(n_301) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_278), .B(n_248), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_292), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_292), .Y(n_304) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_283), .A2(n_254), .B(n_247), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_274), .A2(n_263), .B(n_244), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_278), .Y(n_307) );
AOI21x1_ASAP7_75t_L g308 ( .A1(n_274), .A2(n_244), .B(n_248), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_280), .B(n_248), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_286), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_284), .B(n_244), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_311), .B(n_284), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_311), .B(n_286), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_311), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_298), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_313), .B(n_273), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_298), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_315), .B(n_272), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_293), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_307), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_307), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_297), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_315), .B(n_290), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_313), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_293), .B(n_277), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_299), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_293), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_312), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_295), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_303), .B(n_276), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_312), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_312), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_302), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_303), .B(n_290), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_335), .B(n_299), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_327), .B(n_304), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_318), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_329), .B(n_304), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_329), .B(n_304), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_333), .B(n_302), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_319), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_321), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_327), .B(n_308), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_308), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_328), .B(n_277), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_306), .Y(n_359) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_343), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
OR2x2_ASAP7_75t_L g362 ( .A(n_330), .B(n_314), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_341), .Y(n_364) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_333), .B(n_314), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_333), .Y(n_366) );
INVx3_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_326), .B(n_306), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_324), .B(n_310), .Y(n_369) );
INVx3_ASAP7_75t_L g370 ( .A(n_345), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_342), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_319), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_326), .B(n_306), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_325), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_325), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_320), .A2(n_305), .B(n_301), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_339), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_326), .B(n_305), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_330), .B(n_305), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_317), .B(n_270), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_345), .B(n_276), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_334), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_345), .B(n_305), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_338), .B(n_279), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_338), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_346), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_334), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_331), .B(n_346), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_345), .B(n_301), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_388), .B(n_344), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_388), .B(n_387), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_387), .B(n_331), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_378), .B(n_316), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_371), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_374), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_378), .B(n_316), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_390), .B(n_332), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_356), .B(n_336), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_361), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_356), .B(n_344), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_350), .B(n_337), .Y(n_407) );
INVx2_ASAP7_75t_SL g408 ( .A(n_364), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_361), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
AND2x2_ASAP7_75t_SL g411 ( .A(n_366), .B(n_332), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_348), .B(n_323), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_358), .B(n_332), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_348), .B(n_323), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_363), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_359), .B(n_336), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_363), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_381), .B(n_296), .Y(n_418) );
BUFx2_ASAP7_75t_L g419 ( .A(n_366), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_372), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_349), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_372), .Y(n_422) );
BUFx2_ASAP7_75t_L g423 ( .A(n_366), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_359), .B(n_332), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_357), .B(n_337), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
BUFx2_ASAP7_75t_SL g427 ( .A(n_366), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_374), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_377), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_357), .B(n_340), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_350), .B(n_335), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_380), .B(n_340), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_382), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_352), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_380), .B(n_340), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_375), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_379), .B(n_340), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_365), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_379), .B(n_301), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_368), .B(n_301), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_375), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_368), .B(n_294), .Y(n_442) );
INVx2_ASAP7_75t_SL g443 ( .A(n_365), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_370), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_373), .B(n_294), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_395), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_430), .B(n_352), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_406), .B(n_351), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_L g449 ( .A1(n_410), .A2(n_347), .B(n_386), .C(n_383), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_399), .B(n_373), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_408), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_429), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_399), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_430), .B(n_352), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_411), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_406), .B(n_351), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_408), .B(n_362), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_425), .B(n_362), .Y(n_458) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_411), .A2(n_391), .B(n_385), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_404), .B(n_391), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_431), .B(n_369), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_392), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_438), .B(n_370), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_392), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_432), .B(n_352), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_409), .Y(n_467) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_427), .B(n_370), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_432), .B(n_370), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_419), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_425), .B(n_404), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_417), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_417), .Y(n_475) );
AND2x4_ASAP7_75t_L g476 ( .A(n_423), .B(n_391), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_402), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_429), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_423), .A2(n_383), .B1(n_367), .B2(n_296), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_434), .B(n_391), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_431), .B(n_377), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_397), .B(n_401), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_407), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_427), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_405), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_415), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_394), .Y(n_487) );
OAI32xp33_ASAP7_75t_L g488 ( .A1(n_424), .A2(n_383), .A3(n_367), .B1(n_349), .B2(n_353), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_435), .B(n_367), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_426), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_435), .B(n_385), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_455), .A2(n_434), .B1(n_413), .B2(n_403), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_472), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_449), .A2(n_443), .B(n_438), .Y(n_495) );
NAND3xp33_ASAP7_75t_SL g496 ( .A(n_449), .B(n_418), .C(n_393), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_455), .A2(n_443), .B1(n_396), .B2(n_414), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_472), .B(n_440), .Y(n_498) );
OAI221xp5_ASAP7_75t_SL g499 ( .A1(n_459), .A2(n_437), .B1(n_416), .B2(n_445), .C(n_442), .Y(n_499) );
AOI32xp33_ASAP7_75t_L g500 ( .A1(n_455), .A2(n_414), .A3(n_412), .B1(n_437), .B2(n_416), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_483), .B(n_440), .Y(n_501) );
NAND2xp33_ASAP7_75t_L g502 ( .A(n_484), .B(n_412), .Y(n_502) );
AOI22x1_ASAP7_75t_L g503 ( .A1(n_470), .A2(n_296), .B1(n_444), .B2(n_385), .Y(n_503) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_453), .B(n_441), .C(n_420), .Y(n_504) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_462), .A2(n_445), .B(n_442), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_451), .B(n_393), .Y(n_506) );
NAND4xp25_ASAP7_75t_SL g507 ( .A(n_468), .B(n_407), .C(n_439), .D(n_436), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_480), .A2(n_385), .B1(n_439), .B2(n_444), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_453), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_483), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_463), .Y(n_511) );
NAND3x2_ASAP7_75t_L g512 ( .A(n_480), .B(n_441), .C(n_420), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_479), .A2(n_422), .B1(n_428), .B2(n_400), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_448), .B(n_456), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_446), .B(n_422), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_467), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_473), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_474), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_475), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_458), .B(n_400), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_482), .B(n_428), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_495), .A2(n_479), .B(n_462), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_515), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_495), .A2(n_464), .B(n_476), .C(n_480), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_496), .A2(n_476), .B1(n_457), .B2(n_460), .Y(n_527) );
OAI211xp5_ASAP7_75t_SL g528 ( .A1(n_500), .A2(n_450), .B(n_461), .C(n_485), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g529 ( .A1(n_505), .A2(n_476), .B1(n_471), .B2(n_481), .Y(n_529) );
XNOR2x1_ASAP7_75t_L g530 ( .A(n_497), .B(n_447), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_512), .A2(n_488), .B(n_460), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_501), .B(n_487), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_510), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_502), .A2(n_454), .B(n_466), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_511), .Y(n_535) );
NAND3xp33_ASAP7_75t_SL g536 ( .A(n_509), .B(n_469), .C(n_489), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_493), .A2(n_491), .B1(n_492), .B2(n_490), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_493), .A2(n_486), .B1(n_478), .B2(n_452), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_514), .B(n_478), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_SL g540 ( .A1(n_494), .A2(n_498), .B(n_513), .C(n_504), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_516), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_517), .Y(n_542) );
AOI21xp5_ASAP7_75t_SL g543 ( .A1(n_507), .A2(n_487), .B(n_452), .Y(n_543) );
NOR2x1_ASAP7_75t_L g544 ( .A(n_505), .B(n_398), .Y(n_544) );
NAND4xp75_ASAP7_75t_L g545 ( .A(n_506), .B(n_282), .C(n_398), .D(n_394), .Y(n_545) );
AOI211xp5_ASAP7_75t_L g546 ( .A1(n_499), .A2(n_389), .B(n_384), .C(n_300), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_523), .B(n_376), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_522), .B(n_376), .Y(n_548) );
OAI221xp5_ASAP7_75t_L g549 ( .A1(n_508), .A2(n_389), .B1(n_384), .B2(n_291), .C(n_353), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_503), .A2(n_288), .B1(n_376), .B2(n_271), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_518), .B(n_288), .C(n_271), .Y(n_551) );
NAND5xp2_ASAP7_75t_L g552 ( .A(n_519), .B(n_244), .C(n_271), .D(n_294), .E(n_520), .Y(n_552) );
NOR3xp33_ASAP7_75t_SL g553 ( .A(n_528), .B(n_526), .C(n_524), .Y(n_553) );
NOR5xp2_ASAP7_75t_L g554 ( .A(n_529), .B(n_531), .C(n_533), .D(n_540), .E(n_549), .Y(n_554) );
AOI221xp5_ASAP7_75t_SL g555 ( .A1(n_531), .A2(n_547), .B1(n_534), .B2(n_552), .C(n_525), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_543), .A2(n_527), .B1(n_538), .B2(n_548), .C(n_536), .Y(n_556) );
NAND4xp75_ASAP7_75t_L g557 ( .A(n_544), .B(n_537), .C(n_539), .D(n_541), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_556), .A2(n_530), .B(n_542), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_553), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_557), .B(n_545), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_559), .A2(n_555), .B1(n_554), .B2(n_550), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_560), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_562), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_561), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_564), .A2(n_558), .B(n_535), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_565), .Y(n_566) );
XNOR2xp5_ASAP7_75t_L g567 ( .A(n_566), .B(n_563), .Y(n_567) );
XNOR2xp5_ASAP7_75t_L g568 ( .A(n_567), .B(n_546), .Y(n_568) );
AO21x2_ASAP7_75t_L g569 ( .A1(n_568), .A2(n_551), .B(n_532), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_569), .A2(n_271), .B1(n_521), .B2(n_559), .Y(n_570) );
endmodule