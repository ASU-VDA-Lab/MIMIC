module real_aes_8426_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g171 ( .A1(n_0), .A2(n_172), .B(n_173), .C(n_177), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_1), .B(n_166), .Y(n_179) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_3), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_4), .A2(n_160), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_5), .A2(n_140), .B(n_157), .C(n_513), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_6), .A2(n_160), .B(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_7), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_8), .B(n_166), .Y(n_475) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_9), .A2(n_132), .B(n_254), .Y(n_253) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_10), .A2(n_445), .B1(n_715), .B2(n_718), .C1(n_722), .C2(n_723), .Y(n_444) );
AND2x6_ASAP7_75t_L g157 ( .A(n_11), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_12), .A2(n_140), .B(n_157), .C(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g566 ( .A(n_13), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_14), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_14), .B(n_40), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_15), .B(n_176), .Y(n_515) );
INVx1_ASAP7_75t_L g137 ( .A(n_16), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_17), .B(n_151), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_18), .A2(n_152), .B(n_524), .C(n_526), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_19), .B(n_166), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_20), .B(n_194), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_21), .A2(n_140), .B(n_186), .C(n_193), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_22), .A2(n_175), .B(n_228), .C(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_23), .B(n_176), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_24), .B(n_176), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_25), .Y(n_493) );
INVx1_ASAP7_75t_L g463 ( .A(n_26), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_27), .A2(n_140), .B(n_193), .C(n_257), .Y(n_256) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_28), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_29), .Y(n_511) );
INVx1_ASAP7_75t_L g487 ( .A(n_30), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_31), .A2(n_160), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g142 ( .A(n_32), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_33), .A2(n_155), .B(n_209), .C(n_210), .Y(n_208) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_34), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_35), .A2(n_175), .B(n_472), .C(n_474), .Y(n_471) );
INVxp67_ASAP7_75t_L g488 ( .A(n_36), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_37), .B(n_259), .Y(n_258) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_38), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_39), .A2(n_140), .B(n_193), .C(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_41), .A2(n_177), .B(n_564), .C(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_42), .B(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_43), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_44), .B(n_151), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_45), .B(n_160), .Y(n_255) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_46), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_47), .Y(n_484) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_48), .A2(n_155), .B(n_209), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g174 ( .A(n_49), .Y(n_174) );
INVx1_ASAP7_75t_L g238 ( .A(n_50), .Y(n_238) );
INVx1_ASAP7_75t_L g531 ( .A(n_51), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_52), .B(n_160), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_53), .A2(n_102), .B1(n_114), .B2(n_728), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_54), .A2(n_71), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_54), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_55), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g562 ( .A(n_56), .Y(n_562) );
INVx1_ASAP7_75t_L g158 ( .A(n_57), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_58), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_59), .B(n_166), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_60), .A2(n_147), .B(n_192), .C(n_249), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_61), .A2(n_70), .B1(n_716), .B2(n_717), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_61), .Y(n_716) );
INVx1_ASAP7_75t_L g136 ( .A(n_62), .Y(n_136) );
INVx1_ASAP7_75t_SL g473 ( .A(n_63), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_64), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_65), .B(n_151), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_66), .B(n_166), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_67), .B(n_152), .Y(n_225) );
INVx1_ASAP7_75t_L g496 ( .A(n_68), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_69), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_70), .Y(n_717) );
INVx1_ASAP7_75t_L g124 ( .A(n_71), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_72), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_73), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_74), .Y(n_247) );
INVx1_ASAP7_75t_L g110 ( .A(n_75), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_76), .A2(n_160), .B(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_77), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_78), .A2(n_160), .B(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_79), .A2(n_184), .B(n_483), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_80), .Y(n_460) );
INVx1_ASAP7_75t_L g522 ( .A(n_81), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_82), .B(n_190), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_83), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_84), .A2(n_160), .B(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g525 ( .A(n_85), .Y(n_525) );
INVx2_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g514 ( .A(n_87), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_88), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_89), .B(n_176), .Y(n_226) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_90), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g436 ( .A(n_90), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g449 ( .A(n_90), .B(n_438), .Y(n_449) );
INVx2_ASAP7_75t_L g714 ( .A(n_90), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_91), .A2(n_140), .B(n_155), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_92), .B(n_160), .Y(n_207) );
INVx1_ASAP7_75t_L g211 ( .A(n_93), .Y(n_211) );
INVxp67_ASAP7_75t_L g250 ( .A(n_94), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_95), .B(n_132), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_96), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
INVx1_ASAP7_75t_L g221 ( .A(n_98), .Y(n_221) );
INVx2_ASAP7_75t_L g534 ( .A(n_99), .Y(n_534) );
AND2x2_ASAP7_75t_L g240 ( .A(n_100), .B(n_196), .Y(n_240) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_SL g730 ( .A(n_104), .Y(n_730) );
AND2x2_ASAP7_75t_SL g104 ( .A(n_105), .B(n_111), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g438 ( .A(n_107), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_443), .Y(n_114) );
BUFx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g727 ( .A(n_118), .Y(n_727) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_435), .B(n_440), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx1_ASAP7_75t_L g446 ( .A(n_125), .Y(n_446) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_125), .A2(n_451), .B1(n_719), .B2(n_720), .Y(n_718) );
OR3x1_ASAP7_75t_L g125 ( .A(n_126), .B(n_343), .C(n_392), .Y(n_125) );
NAND5xp2_ASAP7_75t_L g126 ( .A(n_127), .B(n_277), .C(n_306), .D(n_314), .E(n_329), .Y(n_126) );
O2A1O1Ixp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_200), .B(n_216), .C(n_261), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_180), .Y(n_128) );
AND2x2_ASAP7_75t_L g272 ( .A(n_129), .B(n_269), .Y(n_272) );
AND2x2_ASAP7_75t_L g305 ( .A(n_129), .B(n_181), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_129), .B(n_204), .Y(n_398) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
INVx2_ASAP7_75t_L g203 ( .A(n_130), .Y(n_203) );
BUFx2_ASAP7_75t_L g372 ( .A(n_130), .Y(n_372) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_163), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_131), .B(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_131), .B(n_215), .Y(n_214) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_131), .A2(n_220), .B(n_230), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_131), .B(n_466), .Y(n_465) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_131), .A2(n_492), .B(n_499), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_131), .B(n_517), .Y(n_516) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_132), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_132), .A2(n_255), .B(n_256), .Y(n_254) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g232 ( .A(n_133), .Y(n_232) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g196 ( .A(n_134), .B(n_135), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_159), .Y(n_138) );
INVx5_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
BUFx3_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx1_ASAP7_75t_L g229 ( .A(n_142), .Y(n_229) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_144), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_144), .B(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx1_ASAP7_75t_L g259 ( .A(n_144), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_148), .A2(n_151), .B1(n_487), .B2(n_488), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_148), .B(n_525), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_148), .B(n_534), .Y(n_533) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
INVx2_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_151), .B(n_250), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g462 ( .A1(n_151), .A2(n_191), .B(n_463), .C(n_464), .Y(n_462) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_152), .B(n_566), .Y(n_565) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g474 ( .A(n_154), .Y(n_474) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_156), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_156), .A2(n_170), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_156), .A2(n_170), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_156), .A2(n_170), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g521 ( .A1(n_156), .A2(n_170), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_SL g530 ( .A1(n_156), .A2(n_170), .B(n_531), .C(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_SL g561 ( .A1(n_156), .A2(n_170), .B(n_562), .C(n_563), .Y(n_561) );
INVx4_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g160 ( .A(n_157), .B(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
NAND2x1p5_ASAP7_75t_L g222 ( .A(n_157), .B(n_161), .Y(n_222) );
BUFx2_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx1_ASAP7_75t_L g192 ( .A(n_162), .Y(n_192) );
AND2x2_ASAP7_75t_L g180 ( .A(n_165), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g270 ( .A(n_165), .Y(n_270) );
AND2x2_ASAP7_75t_L g356 ( .A(n_165), .B(n_269), .Y(n_356) );
AND2x2_ASAP7_75t_L g411 ( .A(n_165), .B(n_203), .Y(n_411) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_179), .Y(n_165) );
INVx2_ASAP7_75t_L g209 ( .A(n_170), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_175), .B(n_473), .Y(n_472) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g564 ( .A(n_176), .Y(n_564) );
INVx2_ASAP7_75t_L g498 ( .A(n_177), .Y(n_498) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
INVx1_ASAP7_75t_L g526 ( .A(n_178), .Y(n_526) );
INVx1_ASAP7_75t_L g328 ( .A(n_180), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_180), .B(n_204), .Y(n_375) );
INVx5_ASAP7_75t_L g269 ( .A(n_181), .Y(n_269) );
AND2x4_ASAP7_75t_L g290 ( .A(n_181), .B(n_270), .Y(n_290) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_181), .Y(n_312) );
AND2x2_ASAP7_75t_L g387 ( .A(n_181), .B(n_372), .Y(n_387) );
AND2x2_ASAP7_75t_L g390 ( .A(n_181), .B(n_205), .Y(n_390) );
OR2x6_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
AOI21xp5_ASAP7_75t_SL g182 ( .A1(n_183), .A2(n_185), .B(n_194), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_191), .Y(n_186) );
INVx2_ASAP7_75t_L g190 ( .A(n_188), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_190), .A2(n_211), .B(n_212), .C(n_213), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g237 ( .A1(n_190), .A2(n_213), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_190), .A2(n_496), .B(n_497), .C(n_498), .Y(n_495) );
O2A1O1Ixp5_ASAP7_75t_L g513 ( .A1(n_190), .A2(n_498), .B(n_514), .C(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_192), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_195), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_196), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_196), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_196), .A2(n_235), .B(n_236), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g459 ( .A1(n_196), .A2(n_222), .B(n_460), .C(n_461), .Y(n_459) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_196), .A2(n_560), .B(n_567), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_199), .A2(n_510), .B(n_516), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_200), .B(n_270), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_200), .B(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
AND2x2_ASAP7_75t_L g295 ( .A(n_202), .B(n_270), .Y(n_295) );
AND2x2_ASAP7_75t_L g313 ( .A(n_202), .B(n_205), .Y(n_313) );
INVx1_ASAP7_75t_L g333 ( .A(n_202), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_202), .B(n_269), .Y(n_378) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_202), .Y(n_420) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_203), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_204), .B(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_204), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g325 ( .A1(n_204), .A2(n_265), .B(n_326), .C(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g332 ( .A(n_204), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g341 ( .A(n_204), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g345 ( .A(n_204), .B(n_269), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_204), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g360 ( .A(n_204), .B(n_270), .Y(n_360) );
AND2x2_ASAP7_75t_L g410 ( .A(n_204), .B(n_411), .Y(n_410) );
INVx5_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
BUFx2_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
AND2x2_ASAP7_75t_L g315 ( .A(n_205), .B(n_268), .Y(n_315) );
AND2x2_ASAP7_75t_L g327 ( .A(n_205), .B(n_302), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_205), .B(n_356), .Y(n_374) );
OR2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_214), .Y(n_205) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_241), .Y(n_216) );
INVx1_ASAP7_75t_L g263 ( .A(n_217), .Y(n_263) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_233), .Y(n_217) );
OR2x2_ASAP7_75t_L g265 ( .A(n_218), .B(n_233), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_218), .B(n_272), .C(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_218), .B(n_243), .Y(n_282) );
OR2x2_ASAP7_75t_L g297 ( .A(n_218), .B(n_285), .Y(n_297) );
AND2x2_ASAP7_75t_L g303 ( .A(n_218), .B(n_252), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_218), .B(n_434), .Y(n_433) );
INVx5_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_219), .B(n_243), .Y(n_300) );
AND2x2_ASAP7_75t_L g339 ( .A(n_219), .B(n_253), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_219), .B(n_252), .Y(n_367) );
OR2x2_ASAP7_75t_L g370 ( .A(n_219), .B(n_252), .Y(n_370) );
OAI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_223), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_222), .A2(n_493), .B(n_494), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_222), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_227), .A2(n_258), .B(n_260), .Y(n_257) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g481 ( .A(n_232), .Y(n_481) );
INVx5_ASAP7_75t_SL g285 ( .A(n_233), .Y(n_285) );
OR2x2_ASAP7_75t_L g291 ( .A(n_233), .B(n_242), .Y(n_291) );
AND2x2_ASAP7_75t_L g307 ( .A(n_233), .B(n_308), .Y(n_307) );
AOI321xp33_ASAP7_75t_L g314 ( .A1(n_233), .A2(n_315), .A3(n_316), .B1(n_317), .B2(n_323), .C(n_325), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_233), .B(n_241), .Y(n_324) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_233), .Y(n_337) );
OR2x2_ASAP7_75t_L g384 ( .A(n_233), .B(n_282), .Y(n_384) );
AND2x2_ASAP7_75t_L g406 ( .A(n_233), .B(n_303), .Y(n_406) );
AND2x2_ASAP7_75t_L g425 ( .A(n_233), .B(n_243), .Y(n_425) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
INVx1_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_252), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_243), .B(n_252), .Y(n_266) );
AND2x2_ASAP7_75t_L g275 ( .A(n_243), .B(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g302 ( .A(n_243), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_243), .B(n_303), .Y(n_308) );
INVxp67_ASAP7_75t_L g338 ( .A(n_243), .Y(n_338) );
OR2x2_ASAP7_75t_L g380 ( .A(n_243), .B(n_285), .Y(n_380) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_244), .A2(n_468), .B(n_475), .Y(n_467) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_244), .A2(n_520), .B(n_527), .Y(n_519) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_244), .A2(n_529), .B(n_535), .Y(n_528) );
OR2x2_ASAP7_75t_L g262 ( .A(n_252), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_SL g276 ( .A(n_252), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g309 ( .A(n_252), .B(n_265), .Y(n_309) );
AND2x2_ASAP7_75t_L g358 ( .A(n_252), .B(n_302), .Y(n_358) );
AND2x2_ASAP7_75t_L g396 ( .A(n_252), .B(n_285), .Y(n_396) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_253), .B(n_285), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_264), .B(n_267), .C(n_271), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_262), .A2(n_264), .B1(n_389), .B2(n_391), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_264), .A2(n_287), .B1(n_342), .B2(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_SL g416 ( .A(n_265), .Y(n_416) );
INVx1_ASAP7_75t_SL g316 ( .A(n_266), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_268), .B(n_288), .Y(n_318) );
AOI222xp33_ASAP7_75t_L g329 ( .A1(n_268), .A2(n_309), .B1(n_316), .B2(n_330), .C1(n_334), .C2(n_340), .Y(n_329) );
AND2x2_ASAP7_75t_L g419 ( .A(n_268), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g294 ( .A(n_269), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_269), .B(n_289), .Y(n_364) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_269), .Y(n_401) );
AND2x2_ASAP7_75t_L g404 ( .A(n_269), .B(n_313), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_269), .B(n_420), .Y(n_430) );
INVx1_ASAP7_75t_L g321 ( .A(n_270), .Y(n_321) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_270), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g412 ( .A1(n_272), .A2(n_413), .B(n_414), .C(n_417), .Y(n_412) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g335 ( .A(n_274), .B(n_336), .C(n_339), .Y(n_335) );
OR2x2_ASAP7_75t_L g363 ( .A(n_274), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_274), .B(n_290), .Y(n_391) );
OR2x2_ASAP7_75t_L g296 ( .A(n_276), .B(n_297), .Y(n_296) );
AOI211xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B(n_286), .C(n_298), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_279), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g385 ( .A(n_280), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_281), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g299 ( .A(n_284), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_285), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g353 ( .A(n_285), .B(n_303), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_285), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_285), .B(n_302), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B1(n_292), .B2(n_296), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_288), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_290), .B(n_332), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g354 ( .A1(n_291), .A2(n_355), .B1(n_357), .B2(n_359), .C(n_361), .Y(n_354) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AND2x2_ASAP7_75t_L g409 ( .A(n_294), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g422 ( .A(n_294), .B(n_411), .Y(n_422) );
INVx1_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
INVx1_ASAP7_75t_L g413 ( .A(n_296), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_297), .A2(n_380), .B(n_403), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_304), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI21xp5_ASAP7_75t_SL g306 ( .A1(n_307), .A2(n_309), .B(n_310), .Y(n_306) );
INVx1_ASAP7_75t_L g346 ( .A(n_307), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_308), .A2(n_394), .B1(n_397), .B2(n_399), .C(n_402), .Y(n_393) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_316), .A2(n_406), .B1(n_407), .B2(n_409), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g382 ( .A(n_318), .Y(n_382) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp67_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g386 ( .A(n_322), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g351 ( .A(n_327), .Y(n_351) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_332), .B(n_356), .Y(n_408) );
INVxp67_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_338), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_339), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g431 ( .A(n_339), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI211xp5_ASAP7_75t_SL g343 ( .A1(n_344), .A2(n_346), .B(n_347), .C(n_381), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_350), .B(n_354), .C(n_373), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g434 ( .A(n_358), .Y(n_434) );
AND2x2_ASAP7_75t_L g371 ( .A(n_360), .B(n_372), .Y(n_371) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_369), .B2(n_371), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
OR2x2_ASAP7_75t_L g379 ( .A(n_367), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g432 ( .A(n_368), .Y(n_432) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AOI31xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .A3(n_376), .B(n_379), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_385), .C(n_388), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g389 ( .A(n_390), .Y(n_389) );
NAND5xp2_ASAP7_75t_L g392 ( .A(n_393), .B(n_405), .C(n_412), .D(n_426), .E(n_429), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_404), .A2(n_430), .B1(n_431), .B2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_SL g428 ( .A(n_406), .Y(n_428) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B(n_423), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_436), .Y(n_442) );
NOR2x2_ASAP7_75t_L g725 ( .A(n_437), .B(n_714), .Y(n_725) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
OR2x2_ASAP7_75t_L g713 ( .A(n_438), .B(n_714), .Y(n_713) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_440), .B(n_444), .C(n_726), .Y(n_443) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g445 ( .A1(n_446), .A2(n_447), .B1(n_450), .B2(n_713), .Y(n_445) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g719 ( .A(n_448), .Y(n_719) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR3x1_ASAP7_75t_L g451 ( .A(n_452), .B(n_624), .C(n_671), .Y(n_451) );
NAND3xp33_ASAP7_75t_SL g452 ( .A(n_453), .B(n_570), .C(n_595), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_508), .B1(n_536), .B2(n_539), .C(n_547), .Y(n_453) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_476), .B(n_501), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_456), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_456), .B(n_552), .Y(n_668) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_467), .Y(n_456) );
AND2x2_ASAP7_75t_L g538 ( .A(n_457), .B(n_507), .Y(n_538) );
AND2x2_ASAP7_75t_L g588 ( .A(n_457), .B(n_506), .Y(n_588) );
AND2x2_ASAP7_75t_L g609 ( .A(n_457), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g614 ( .A(n_457), .B(n_581), .Y(n_614) );
OR2x2_ASAP7_75t_L g622 ( .A(n_457), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g694 ( .A(n_457), .B(n_490), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_457), .B(n_643), .Y(n_708) );
INVx3_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g553 ( .A(n_458), .B(n_467), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_458), .B(n_490), .Y(n_554) );
AND2x4_ASAP7_75t_L g576 ( .A(n_458), .B(n_507), .Y(n_576) );
AND2x2_ASAP7_75t_L g606 ( .A(n_458), .B(n_478), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_458), .B(n_605), .Y(n_615) );
AND2x2_ASAP7_75t_L g631 ( .A(n_458), .B(n_491), .Y(n_631) );
OR2x2_ASAP7_75t_L g640 ( .A(n_458), .B(n_623), .Y(n_640) );
AND2x2_ASAP7_75t_L g646 ( .A(n_458), .B(n_581), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_458), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g660 ( .A(n_458), .B(n_503), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_458), .B(n_549), .Y(n_670) );
NAND2xp5_ASAP7_75t_SL g699 ( .A(n_458), .B(n_610), .Y(n_699) );
OR2x6_ASAP7_75t_L g458 ( .A(n_459), .B(n_465), .Y(n_458) );
INVx2_ASAP7_75t_L g507 ( .A(n_467), .Y(n_507) );
AND2x2_ASAP7_75t_L g605 ( .A(n_467), .B(n_490), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_467), .B(n_491), .Y(n_610) );
INVx1_ASAP7_75t_L g666 ( .A(n_467), .Y(n_666) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g575 ( .A(n_477), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_478), .B(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
OR2x2_ASAP7_75t_L g623 ( .A(n_478), .B(n_490), .Y(n_623) );
OR2x2_ASAP7_75t_L g684 ( .A(n_478), .B(n_591), .Y(n_684) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_482), .B(n_489), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_480), .A2(n_504), .B(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g504 ( .A(n_482), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_489), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_490), .B(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g643 ( .A(n_490), .B(n_503), .Y(n_643) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g582 ( .A(n_491), .Y(n_582) );
INVx1_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_502), .A2(n_688), .B1(n_692), .B2(n_695), .C(n_696), .Y(n_687) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
INVx1_ASAP7_75t_SL g550 ( .A(n_503), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_503), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_503), .B(n_538), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_506), .B(n_552), .Y(n_674) );
AND2x2_ASAP7_75t_L g581 ( .A(n_507), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_SL g585 ( .A(n_508), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_508), .B(n_591), .Y(n_621) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
AND2x2_ASAP7_75t_L g546 ( .A(n_509), .B(n_519), .Y(n_546) );
INVx4_ASAP7_75t_L g558 ( .A(n_509), .Y(n_558) );
BUFx3_ASAP7_75t_L g601 ( .A(n_509), .Y(n_601) );
AND3x2_ASAP7_75t_L g616 ( .A(n_509), .B(n_617), .C(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g698 ( .A(n_518), .B(n_612), .Y(n_698) );
AND2x2_ASAP7_75t_L g706 ( .A(n_518), .B(n_591), .Y(n_706) );
INVx1_ASAP7_75t_SL g711 ( .A(n_518), .Y(n_711) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
INVx1_ASAP7_75t_SL g569 ( .A(n_519), .Y(n_569) );
AND2x2_ASAP7_75t_L g592 ( .A(n_519), .B(n_558), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_519), .B(n_542), .Y(n_594) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_519), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_519), .B(n_558), .Y(n_639) );
INVx2_ASAP7_75t_L g544 ( .A(n_528), .Y(n_544) );
AND2x2_ASAP7_75t_L g579 ( .A(n_528), .B(n_559), .Y(n_579) );
OR2x2_ASAP7_75t_L g599 ( .A(n_528), .B(n_559), .Y(n_599) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_528), .Y(n_619) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_537), .A2(n_578), .B(n_670), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g705 ( .A1(n_539), .A2(n_549), .A3(n_576), .B1(n_706), .B2(n_707), .C1(n_709), .C2(n_712), .Y(n_705) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_541), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_542), .B(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g568 ( .A(n_543), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g636 ( .A(n_544), .B(n_558), .Y(n_636) );
AND2x2_ASAP7_75t_L g703 ( .A(n_544), .B(n_559), .Y(n_703) );
INVx1_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g644 ( .A(n_546), .B(n_598), .Y(n_644) );
AOI31xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_551), .A3(n_554), .B(n_555), .Y(n_547) );
AND2x2_ASAP7_75t_L g603 ( .A(n_549), .B(n_581), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_549), .B(n_573), .Y(n_685) );
AND2x2_ASAP7_75t_L g704 ( .A(n_549), .B(n_609), .Y(n_704) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_552), .B(n_581), .Y(n_593) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_552), .B(n_610), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_552), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_552), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_553), .B(n_610), .Y(n_642) );
INVx1_ASAP7_75t_L g686 ( .A(n_553), .Y(n_686) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_568), .Y(n_556) );
INVxp67_ASAP7_75t_L g638 ( .A(n_557), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_558), .B(n_569), .Y(n_574) );
INVx1_ASAP7_75t_L g680 ( .A(n_558), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_558), .B(n_657), .Y(n_691) );
BUFx3_ASAP7_75t_L g591 ( .A(n_559), .Y(n_591) );
AND2x2_ASAP7_75t_L g617 ( .A(n_559), .B(n_569), .Y(n_617) );
INVx2_ASAP7_75t_L g657 ( .A(n_559), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_568), .B(n_690), .Y(n_689) );
AOI211xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_575), .B(n_577), .C(n_586), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g620 ( .A1(n_572), .A2(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_573), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_573), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g653 ( .A(n_574), .B(n_599), .Y(n_653) );
INVx3_ASAP7_75t_L g584 ( .A(n_576), .Y(n_584) );
OAI22xp5_ASAP7_75t_SL g577 ( .A1(n_578), .A2(n_580), .B1(n_583), .B2(n_585), .Y(n_577) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_579), .A2(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g628 ( .A(n_579), .B(n_592), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_579), .B(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g583 ( .A(n_582), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g652 ( .A(n_582), .Y(n_652) );
OAI21xp5_ASAP7_75t_SL g596 ( .A1(n_583), .A2(n_597), .B(n_602), .Y(n_596) );
OAI22xp33_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_589), .B1(n_593), .B2(n_594), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_588), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_591), .B(n_634), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_607), .C(n_620), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g662 ( .A1(n_597), .A2(n_663), .B1(n_667), .B2(n_668), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g667 ( .A(n_599), .B(n_600), .Y(n_667) );
AND2x2_ASAP7_75t_L g675 ( .A(n_600), .B(n_656), .Y(n_675) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_601), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_SL g683 ( .A1(n_601), .A2(n_684), .B(n_685), .C(n_686), .Y(n_683) );
OR2x2_ASAP7_75t_L g710 ( .A(n_601), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_611), .B(n_613), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g645 ( .A1(n_609), .A2(n_646), .B(n_647), .C(n_650), .Y(n_645) );
OAI21xp33_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_615), .B(n_616), .Y(n_613) );
AND2x2_ASAP7_75t_L g678 ( .A(n_617), .B(n_636), .Y(n_678) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g656 ( .A(n_619), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_645), .C(n_658), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B(n_629), .C(n_637), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
INVx1_ASAP7_75t_L g695 ( .A(n_632), .Y(n_695) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_634), .B(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B(n_640), .C(n_641), .Y(n_637) );
INVx2_ASAP7_75t_SL g649 ( .A(n_639), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_640), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_650) );
OAI21xp33_ASAP7_75t_SL g641 ( .A1(n_642), .A2(n_643), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_661), .B(n_662), .C(n_669), .Y(n_658) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVxp33_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g712 ( .A(n_666), .Y(n_712) );
NAND4xp25_ASAP7_75t_L g671 ( .A(n_672), .B(n_687), .C(n_700), .D(n_705), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_676), .C(n_683), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_681), .Y(n_676) );
AOI21xp33_ASAP7_75t_L g696 ( .A1(n_677), .A2(n_697), .B(n_699), .Y(n_696) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_684), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g721 ( .A(n_713), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_715), .Y(n_722) );
INVx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
INVx3_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
endmodule