module fake_netlist_5_1330_n_1446 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1446);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1446;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_759;
wire n_806;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_968;
wire n_912;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_1050;
wire n_841;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_176),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_106),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_73),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_23),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_161),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_175),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_50),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_84),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_240),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_59),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_114),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_184),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_45),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_197),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g344 ( 
.A(n_49),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_19),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_4),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_178),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_316),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_293),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_186),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_77),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_110),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_196),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_78),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_247),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_30),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_188),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_43),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_17),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_111),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_166),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_16),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_86),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_282),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_259),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_85),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_45),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_214),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_126),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_66),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_26),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_206),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_89),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_79),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_292),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_142),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_30),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_160),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_269),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_151),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_319),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_217),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_104),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_156),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_288),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_177),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g390 ( 
.A(n_123),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_54),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_24),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_50),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_241),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_210),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_24),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_42),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_265),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_213),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_21),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_135),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_39),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_315),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_164),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_117),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_239),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_81),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_174),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_100),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_250),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_279),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_202),
.Y(n_412)
);

CKINVDCx12_ASAP7_75t_R g413 ( 
.A(n_9),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_91),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_194),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_41),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_246),
.Y(n_417)
);

BUFx2_ASAP7_75t_SL g418 ( 
.A(n_69),
.Y(n_418)
);

BUFx10_ASAP7_75t_L g419 ( 
.A(n_273),
.Y(n_419)
);

CKINVDCx14_ASAP7_75t_R g420 ( 
.A(n_183),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_19),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_271),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_201),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_43),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_18),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_134),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_172),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_41),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_291),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_304),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_289),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_108),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_260),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_7),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_228),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_237),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_171),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_270),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_224),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_252),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_3),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_243),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_234),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_32),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_38),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_267),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_261),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_0),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_52),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_28),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_147),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_70),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_94),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_44),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_119),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_195),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_105),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_153),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_93),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_162),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_131),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_216),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_308),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_39),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_248),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_102),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_154),
.Y(n_467)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_51),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_249),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_208),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_87),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_180),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_90),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_231),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_258),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_98),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_64),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_143),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_109),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_286),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_276),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_185),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_139),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_80),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_7),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_12),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_57),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g488 ( 
.A(n_294),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_125),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_51),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_6),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_55),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_173),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_2),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_74),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_116),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_170),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_5),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_320),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_21),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_14),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_124),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_6),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_15),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_107),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_204),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_127),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_132),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_2),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_168),
.Y(n_510)
);

BUFx10_ASAP7_75t_L g511 ( 
.A(n_11),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_62),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_150),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_181),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_302),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_33),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_314),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_11),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_344),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_484),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_481),
.B(n_0),
.Y(n_521)
);

BUFx12f_ASAP7_75t_L g522 ( 
.A(n_511),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_1),
.Y(n_523)
);

BUFx12f_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_340),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_445),
.B(n_1),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_340),
.B(n_3),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_484),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_484),
.Y(n_530)
);

BUFx8_ASAP7_75t_SL g531 ( 
.A(n_392),
.Y(n_531)
);

INVx6_ASAP7_75t_L g532 ( 
.A(n_366),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_467),
.B(n_4),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_516),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_391),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_392),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_420),
.B(n_5),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_347),
.B(n_8),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_488),
.B(n_8),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_484),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_391),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_505),
.B(n_9),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_518),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_505),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_357),
.B(n_10),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_467),
.B(n_344),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_329),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_391),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_468),
.B(n_417),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

INVx5_ASAP7_75t_L g552 ( 
.A(n_366),
.Y(n_552)
);

INVx5_ASAP7_75t_L g553 ( 
.A(n_366),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_499),
.B(n_10),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_330),
.B(n_12),
.Y(n_555)
);

BUFx12f_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_353),
.B(n_13),
.Y(n_557)
);

BUFx12f_ASAP7_75t_L g558 ( 
.A(n_419),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_419),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_428),
.B(n_13),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_335),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_395),
.B(n_14),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_330),
.Y(n_563)
);

BUFx12f_ASAP7_75t_L g564 ( 
.A(n_419),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_375),
.B(n_15),
.Y(n_565)
);

BUFx8_ASAP7_75t_SL g566 ( 
.A(n_448),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_375),
.B(n_16),
.Y(n_567)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_518),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_338),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_333),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_408),
.B(n_17),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_348),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_408),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_427),
.B(n_18),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_427),
.B(n_20),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g576 ( 
.A(n_331),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_334),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_342),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_447),
.B(n_20),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_345),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_336),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_390),
.B(n_22),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_337),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_459),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_346),
.B(n_22),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_351),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_360),
.B(n_23),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_363),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_339),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_354),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_448),
.B(n_25),
.Y(n_593)
);

BUFx8_ASAP7_75t_SL g594 ( 
.A(n_485),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_364),
.B(n_370),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_371),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_341),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_390),
.B(n_25),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_413),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_372),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_381),
.B(n_26),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_435),
.B(n_27),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_359),
.B(n_27),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_398),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_348),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_373),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_396),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_352),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_397),
.B(n_28),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_424),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_399),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_332),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_407),
.B(n_411),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_349),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_414),
.B(n_422),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_450),
.B(n_29),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_423),
.B(n_426),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_433),
.B(n_29),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_368),
.B(n_31),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_453),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_452),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_454),
.B(n_31),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_457),
.B(n_32),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_492),
.B(n_33),
.Y(n_624)
);

BUFx8_ASAP7_75t_SL g625 ( 
.A(n_485),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_349),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_494),
.B(n_34),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_512),
.Y(n_628)
);

BUFx8_ASAP7_75t_L g629 ( 
.A(n_463),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_469),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_471),
.Y(n_631)
);

BUFx8_ASAP7_75t_SL g632 ( 
.A(n_343),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_474),
.B(n_34),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_550),
.B(n_350),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_541),
.Y(n_635)
);

OA22x2_ASAP7_75t_L g636 ( 
.A1(n_519),
.A2(n_393),
.B1(n_400),
.B2(n_380),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_SL g637 ( 
.A1(n_584),
.A2(n_356),
.B1(n_358),
.B2(n_343),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_548),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_548),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_532),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_554),
.A2(n_416),
.B1(n_421),
.B2(n_402),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_537),
.A2(n_356),
.B1(n_405),
.B2(n_358),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_539),
.A2(n_405),
.B1(n_446),
.B2(n_412),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_548),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_549),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_554),
.A2(n_434),
.B1(n_441),
.B2(n_425),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_549),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_549),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_576),
.B(n_350),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_523),
.B(n_412),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_552),
.B(n_446),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_535),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_SL g653 ( 
.A1(n_593),
.A2(n_444),
.B1(n_477),
.B2(n_464),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_593),
.A2(n_490),
.B1(n_491),
.B2(n_486),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_520),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_520),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_598),
.A2(n_461),
.B1(n_470),
.B2(n_498),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_532),
.A2(n_501),
.B1(n_503),
.B2(n_500),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_521),
.A2(n_504),
.B1(n_509),
.B2(n_487),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_533),
.A2(n_461),
.B1(n_470),
.B2(n_517),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_520),
.Y(n_661)
);

AO22x2_ASAP7_75t_L g662 ( 
.A1(n_527),
.A2(n_418),
.B1(n_479),
.B2(n_476),
.Y(n_662)
);

OAI22xp33_ASAP7_75t_L g663 ( 
.A1(n_533),
.A2(n_517),
.B1(n_432),
.B2(n_495),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_529),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_560),
.A2(n_432),
.B1(n_496),
.B2(n_480),
.Y(n_665)
);

AO22x2_ASAP7_75t_L g666 ( 
.A1(n_527),
.A2(n_542),
.B1(n_526),
.B2(n_545),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_529),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_632),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_538),
.A2(n_361),
.B1(n_362),
.B2(n_355),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_546),
.A2(n_506),
.B1(n_508),
.B2(n_497),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_557),
.A2(n_367),
.B1(n_369),
.B2(n_365),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_602),
.A2(n_376),
.B1(n_377),
.B2(n_374),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_560),
.A2(n_513),
.B1(n_514),
.B2(n_510),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_562),
.A2(n_379),
.B1(n_382),
.B2(n_378),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_528),
.B(n_35),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_578),
.B(n_515),
.Y(n_676)
);

BUFx6f_ASAP7_75t_SL g677 ( 
.A(n_542),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_562),
.A2(n_384),
.B1(n_385),
.B2(n_383),
.Y(n_678)
);

OA22x2_ASAP7_75t_L g679 ( 
.A1(n_519),
.A2(n_387),
.B1(n_388),
.B2(n_386),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_SL g680 ( 
.A1(n_546),
.A2(n_394),
.B1(n_401),
.B2(n_389),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_529),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_612),
.B(n_403),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_572),
.B(n_404),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_583),
.B(n_406),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_530),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_530),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_572),
.B(n_409),
.Y(n_687)
);

OAI22xp33_ASAP7_75t_L g688 ( 
.A1(n_567),
.A2(n_507),
.B1(n_502),
.B2(n_493),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_567),
.A2(n_489),
.B1(n_483),
.B2(n_482),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_568),
.A2(n_443),
.B1(n_475),
.B2(n_473),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_530),
.Y(n_691)
);

AO22x2_ASAP7_75t_L g692 ( 
.A1(n_555),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_534),
.A2(n_478),
.B1(n_472),
.B2(n_466),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_603),
.A2(n_465),
.B1(n_462),
.B2(n_460),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_525),
.B(n_410),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_547),
.B(n_415),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_540),
.Y(n_697)
);

AO22x2_ASAP7_75t_L g698 ( 
.A1(n_555),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_619),
.A2(n_458),
.B1(n_456),
.B2(n_455),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_575),
.A2(n_451),
.B1(n_442),
.B2(n_440),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_543),
.A2(n_439),
.B1(n_438),
.B2(n_437),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_570),
.B(n_429),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_540),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_575),
.A2(n_436),
.B1(n_431),
.B2(n_430),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_580),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_552),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_707)
);

OA22x2_ASAP7_75t_L g708 ( 
.A1(n_551),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_558),
.A2(n_564),
.B1(n_559),
.B2(n_524),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_585),
.B(n_75),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_580),
.A2(n_553),
.B1(n_552),
.B2(n_587),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_522),
.A2(n_48),
.B1(n_49),
.B2(n_52),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_544),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_552),
.A2(n_553),
.B1(n_589),
.B2(n_587),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_544),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_553),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_608),
.B(n_76),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_544),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_591),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_553),
.B(n_82),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_597),
.B(n_56),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_563),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_696),
.B(n_702),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_635),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_720),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_722),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_722),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_656),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_652),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_656),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_661),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_642),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_661),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_641),
.B(n_605),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_691),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_688),
.B(n_565),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_691),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_634),
.B(n_599),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_703),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_649),
.B(n_599),
.Y(n_740)
);

INVxp67_ASAP7_75t_SL g741 ( 
.A(n_715),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_703),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_706),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_666),
.A2(n_613),
.B(n_595),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_664),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_706),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_715),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_643),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_667),
.Y(n_749)
);

INVxp33_ASAP7_75t_L g750 ( 
.A(n_657),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_667),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_681),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_685),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_676),
.B(n_605),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_695),
.B(n_599),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_686),
.Y(n_756)
);

INVx4_ASAP7_75t_SL g757 ( 
.A(n_677),
.Y(n_757)
);

XOR2xp5_ASAP7_75t_L g758 ( 
.A(n_668),
.B(n_531),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_682),
.B(n_599),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_697),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_646),
.B(n_605),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_689),
.B(n_565),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_654),
.B(n_605),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_678),
.B(n_614),
.Y(n_764)
);

XOR2xp5_ASAP7_75t_L g765 ( 
.A(n_709),
.B(n_637),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_713),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_718),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_647),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_638),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_639),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_644),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_645),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_648),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_678),
.B(n_614),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_655),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_655),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_655),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_676),
.B(n_614),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_666),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_675),
.B(n_551),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_693),
.B(n_614),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_694),
.A2(n_615),
.B(n_613),
.Y(n_783)
);

AND2x2_ASAP7_75t_SL g784 ( 
.A(n_650),
.B(n_571),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_640),
.B(n_595),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_701),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_700),
.B(n_626),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_704),
.B(n_663),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_687),
.B(n_617),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_677),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_699),
.A2(n_617),
.B(n_601),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_R g792 ( 
.A(n_684),
.B(n_601),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_710),
.A2(n_633),
.B(n_623),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_717),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_684),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_651),
.B(n_626),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_679),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_690),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_683),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_662),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_680),
.B(n_571),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_660),
.B(n_626),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_670),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_636),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_672),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_674),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_708),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_692),
.Y(n_808)
);

INVxp33_ASAP7_75t_L g809 ( 
.A(n_659),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_724),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_724),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_729),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_789),
.B(n_692),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_729),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_784),
.B(n_698),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_784),
.B(n_698),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_793),
.B(n_669),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_795),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_807),
.B(n_623),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_785),
.Y(n_820)
);

BUFx4f_ASAP7_75t_L g821 ( 
.A(n_803),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_807),
.B(n_633),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_780),
.Y(n_823)
);

OR2x2_ASAP7_75t_SL g824 ( 
.A(n_723),
.B(n_653),
.Y(n_824)
);

NAND2x1p5_ASAP7_75t_L g825 ( 
.A(n_796),
.B(n_797),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_799),
.B(n_671),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_781),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_776),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_783),
.B(n_628),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_806),
.B(n_721),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_740),
.B(n_628),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_759),
.B(n_574),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_794),
.B(n_574),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_808),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_791),
.B(n_569),
.Y(n_835)
);

INVx4_ASAP7_75t_L g836 ( 
.A(n_725),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_786),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_745),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_738),
.B(n_600),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_804),
.B(n_600),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_776),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_809),
.B(n_763),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_745),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_764),
.B(n_536),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_769),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_736),
.A2(n_762),
.B(n_744),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_800),
.B(n_788),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_732),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_769),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_726),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_727),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_801),
.B(n_561),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_728),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_730),
.Y(n_854)
);

BUFx2_ASAP7_75t_R g855 ( 
.A(n_736),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_788),
.B(n_579),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_731),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_763),
.B(n_658),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_725),
.B(n_626),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_762),
.A2(n_665),
.B(n_673),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_734),
.A2(n_618),
.B1(n_719),
.B2(n_705),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_733),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_725),
.B(n_764),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_775),
.A2(n_711),
.B(n_714),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_775),
.B(n_582),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_755),
.B(n_590),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_735),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_737),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_801),
.B(n_606),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_734),
.B(n_761),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_748),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_739),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_761),
.B(n_607),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_742),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_743),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_802),
.B(n_610),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_766),
.B(n_621),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_802),
.B(n_618),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_767),
.B(n_589),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_746),
.Y(n_880)
);

AND2x6_ASAP7_75t_L g881 ( 
.A(n_787),
.B(n_712),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_R g882 ( 
.A(n_792),
.B(n_556),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_787),
.A2(n_782),
.B(n_779),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_725),
.B(n_563),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_782),
.B(n_566),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_779),
.B(n_609),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_741),
.B(n_609),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_752),
.B(n_616),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_768),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_770),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_753),
.B(n_616),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_756),
.Y(n_892)
);

INVx1_ASAP7_75t_SL g893 ( 
.A(n_758),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_725),
.B(n_563),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_760),
.B(n_622),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_771),
.B(n_622),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_772),
.B(n_773),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_774),
.B(n_624),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_754),
.B(n_624),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_747),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_777),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_749),
.Y(n_902)
);

AND2x2_ASAP7_75t_SL g903 ( 
.A(n_750),
.B(n_627),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_751),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_842),
.B(n_757),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_887),
.B(n_725),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_837),
.B(n_805),
.Y(n_907)
);

OR2x2_ASAP7_75t_L g908 ( 
.A(n_827),
.B(n_790),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_843),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_SL g910 ( 
.A(n_855),
.B(n_594),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_831),
.B(n_757),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_887),
.B(n_778),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_831),
.B(n_757),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_848),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_843),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_873),
.B(n_798),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_886),
.B(n_573),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_843),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_818),
.B(n_627),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_818),
.B(n_83),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_829),
.B(n_707),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_886),
.B(n_829),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_882),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_825),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_870),
.B(n_573),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_824),
.B(n_765),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_870),
.B(n_573),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_826),
.B(n_625),
.Y(n_928)
);

CKINVDCx14_ASAP7_75t_R g929 ( 
.A(n_871),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_818),
.B(n_88),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_810),
.Y(n_931)
);

CKINVDCx14_ASAP7_75t_R g932 ( 
.A(n_871),
.Y(n_932)
);

BUFx4f_ASAP7_75t_L g933 ( 
.A(n_825),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_834),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_823),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_847),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_835),
.B(n_581),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_820),
.B(n_92),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_820),
.B(n_95),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_834),
.Y(n_940)
);

OR2x6_ASAP7_75t_L g941 ( 
.A(n_815),
.B(n_792),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_847),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_815),
.B(n_816),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_SL g944 ( 
.A(n_830),
.B(n_716),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_SL g945 ( 
.A(n_844),
.B(n_629),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_856),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_856),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_823),
.B(n_96),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_865),
.B(n_899),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_823),
.B(n_852),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_845),
.Y(n_951)
);

NAND2x1_ASAP7_75t_L g952 ( 
.A(n_836),
.B(n_581),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_845),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_865),
.B(n_586),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_836),
.B(n_586),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_845),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_840),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_849),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_824),
.B(n_588),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_852),
.B(n_97),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_852),
.B(n_99),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_849),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_816),
.B(n_588),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_899),
.B(n_586),
.Y(n_964)
);

AND2x6_ASAP7_75t_L g965 ( 
.A(n_863),
.B(n_588),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_853),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_SL g967 ( 
.A(n_885),
.B(n_629),
.Y(n_967)
);

CKINVDCx6p67_ASAP7_75t_R g968 ( 
.A(n_903),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_813),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_828),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_811),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_893),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_899),
.B(n_592),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_811),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_878),
.B(n_592),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_853),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_SL g977 ( 
.A(n_903),
.B(n_592),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_878),
.B(n_596),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_840),
.Y(n_979)
);

BUFx6f_ASAP7_75t_SL g980 ( 
.A(n_934),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_940),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_935),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_970),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_971),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_971),
.Y(n_985)
);

BUFx2_ASAP7_75t_SL g986 ( 
.A(n_972),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_935),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_922),
.A2(n_881),
.B1(n_860),
.B2(n_903),
.Y(n_988)
);

BUFx6f_ASAP7_75t_SL g989 ( 
.A(n_941),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_974),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_935),
.Y(n_991)
);

BUFx4f_ASAP7_75t_SL g992 ( 
.A(n_914),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_950),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_909),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_950),
.Y(n_995)
);

INVx5_ASAP7_75t_L g996 ( 
.A(n_920),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_909),
.Y(n_997)
);

CKINVDCx16_ASAP7_75t_R g998 ( 
.A(n_910),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_943),
.Y(n_999)
);

BUFx3_ASAP7_75t_L g1000 ( 
.A(n_957),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_924),
.Y(n_1001)
);

INVx8_ASAP7_75t_L g1002 ( 
.A(n_943),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_979),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_920),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_936),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_908),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_924),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_916),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_933),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_915),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_933),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_946),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_942),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_930),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_974),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_942),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_960),
.B(n_852),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_930),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_929),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_947),
.B(n_858),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_926),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_969),
.B(n_873),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_960),
.Y(n_1023)
);

INVx5_ASAP7_75t_SL g1024 ( 
.A(n_963),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_931),
.Y(n_1025)
);

BUFx3_ASAP7_75t_L g1026 ( 
.A(n_942),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_975),
.B(n_876),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_970),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_948),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_932),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_923),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_938),
.Y(n_1032)
);

INVx2_ASAP7_75t_SL g1033 ( 
.A(n_938),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_948),
.Y(n_1034)
);

BUFx8_ASAP7_75t_L g1035 ( 
.A(n_911),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_939),
.Y(n_1036)
);

BUFx2_ASAP7_75t_L g1037 ( 
.A(n_963),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_941),
.Y(n_1038)
);

INVx6_ASAP7_75t_L g1039 ( 
.A(n_939),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_915),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_961),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_919),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_918),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_961),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_913),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_988),
.A2(n_881),
.B1(n_944),
.B2(n_968),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_992),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_981),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_988),
.A2(n_881),
.B1(n_817),
.B2(n_921),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_1030),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1025),
.Y(n_1051)
);

CKINVDCx11_ASAP7_75t_R g1052 ( 
.A(n_1030),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_1008),
.B(n_1022),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_986),
.Y(n_1054)
);

BUFx8_ASAP7_75t_L g1055 ( 
.A(n_980),
.Y(n_1055)
);

INVxp67_ASAP7_75t_SL g1056 ( 
.A(n_1014),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_984),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_985),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_990),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1017),
.A2(n_881),
.B1(n_883),
.B2(n_821),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_1017),
.A2(n_881),
.B1(n_821),
.B2(n_864),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1023),
.A2(n_821),
.B1(n_949),
.B2(n_906),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_994),
.Y(n_1063)
);

INVx6_ASAP7_75t_L g1064 ( 
.A(n_1035),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_1001),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1020),
.B(n_919),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1023),
.A2(n_996),
.B1(n_1004),
.B2(n_1039),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_1031),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_994),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1023),
.A2(n_836),
.B(n_846),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_996),
.A2(n_978),
.B1(n_927),
.B2(n_925),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_997),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1021),
.A2(n_928),
.B1(n_907),
.B2(n_881),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1020),
.B(n_876),
.Y(n_1074)
);

CKINVDCx11_ASAP7_75t_R g1075 ( 
.A(n_1031),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_1019),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_992),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1017),
.A2(n_881),
.B1(n_813),
.B2(n_861),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_997),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_1038),
.A2(n_861),
.B1(n_959),
.B2(n_869),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_989),
.A2(n_869),
.B1(n_977),
.B2(n_905),
.Y(n_1081)
);

INVx6_ASAP7_75t_L g1082 ( 
.A(n_1035),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_983),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_996),
.A2(n_912),
.B1(n_954),
.B2(n_917),
.Y(n_1084)
);

BUFx8_ASAP7_75t_L g1085 ( 
.A(n_980),
.Y(n_1085)
);

CKINVDCx6p67_ASAP7_75t_R g1086 ( 
.A(n_980),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_981),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_996),
.A2(n_836),
.B1(n_825),
.B2(n_937),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_989),
.A2(n_879),
.B1(n_832),
.B2(n_833),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1010),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1015),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_989),
.A2(n_879),
.B1(n_832),
.B2(n_833),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_1006),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1000),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_1000),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_983),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1010),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_SL g1098 ( 
.A1(n_1024),
.A2(n_967),
.B1(n_945),
.B2(n_866),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1042),
.A2(n_879),
.B1(n_866),
.B2(n_839),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1003),
.Y(n_1100)
);

OAI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1027),
.A2(n_850),
.B1(n_867),
.B2(n_851),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1040),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1042),
.A2(n_879),
.B1(n_839),
.B2(n_888),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_999),
.A2(n_888),
.B1(n_896),
.B2(n_895),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1040),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1004),
.A2(n_958),
.B1(n_962),
.B2(n_872),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1004),
.A2(n_862),
.B1(n_872),
.B2(n_867),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_SL g1108 ( 
.A1(n_1024),
.A2(n_896),
.B1(n_895),
.B2(n_898),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_SL g1109 ( 
.A(n_1003),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_SL g1110 ( 
.A1(n_1024),
.A2(n_1035),
.B1(n_1002),
.B2(n_998),
.Y(n_1110)
);

INVxp67_ASAP7_75t_SL g1111 ( 
.A(n_1014),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1073),
.A2(n_1045),
.B1(n_1018),
.B2(n_1029),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1049),
.B(n_973),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1064),
.A2(n_1082),
.B1(n_1085),
.B2(n_1055),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1063),
.B(n_1043),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1046),
.A2(n_1108),
.B1(n_1061),
.B2(n_1066),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1060),
.A2(n_1005),
.B1(n_1045),
.B2(n_1044),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_SL g1118 ( 
.A1(n_1064),
.A2(n_1002),
.B1(n_1018),
.B2(n_1014),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_L g1119 ( 
.A1(n_1078),
.A2(n_1005),
.B1(n_1044),
.B2(n_1041),
.Y(n_1119)
);

CKINVDCx11_ASAP7_75t_R g1120 ( 
.A(n_1068),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_1048),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1074),
.B(n_964),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1083),
.Y(n_1123)
);

OAI222xp33_ASAP7_75t_L g1124 ( 
.A1(n_1080),
.A2(n_1036),
.B1(n_1032),
.B2(n_1033),
.C1(n_1012),
.C2(n_1037),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1063),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1065),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_1075),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1062),
.A2(n_898),
.B(n_891),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1081),
.A2(n_1039),
.B1(n_1041),
.B2(n_1014),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1104),
.A2(n_1039),
.B1(n_1029),
.B2(n_1034),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1089),
.A2(n_1029),
.B1(n_1034),
.B2(n_1018),
.Y(n_1131)
);

BUFx4f_ASAP7_75t_SL g1132 ( 
.A(n_1077),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1092),
.A2(n_1002),
.B1(n_1029),
.B2(n_1018),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1103),
.A2(n_1034),
.B1(n_1033),
.B2(n_1032),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1099),
.A2(n_1034),
.B1(n_1036),
.B2(n_1016),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_1075),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1053),
.B(n_891),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1098),
.A2(n_1002),
.B1(n_993),
.B2(n_995),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1093),
.A2(n_1101),
.B1(n_1110),
.B2(n_1016),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1051),
.A2(n_1026),
.B1(n_1013),
.B2(n_1007),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1064),
.A2(n_1007),
.B1(n_1009),
.B2(n_1001),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1082),
.A2(n_993),
.B1(n_995),
.B2(n_877),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_1082),
.A2(n_1007),
.B1(n_1009),
.B2(n_1001),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1069),
.B(n_1043),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1057),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_1055),
.A2(n_1001),
.B1(n_1007),
.B2(n_1009),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1052),
.A2(n_993),
.B1(n_995),
.B2(n_877),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1094),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1052),
.A2(n_877),
.B1(n_851),
.B2(n_862),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1055),
.A2(n_1011),
.B1(n_1009),
.B2(n_1019),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1070),
.A2(n_1026),
.B1(n_1013),
.B2(n_1011),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1050),
.A2(n_889),
.B1(n_850),
.B2(n_857),
.Y(n_1152)
);

OAI222xp33_ASAP7_75t_L g1153 ( 
.A1(n_1054),
.A2(n_889),
.B1(n_976),
.B2(n_966),
.C1(n_991),
.C2(n_902),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1069),
.B(n_983),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1054),
.A2(n_1011),
.B1(n_1028),
.B2(n_991),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_SL g1156 ( 
.A(n_1077),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1085),
.A2(n_1011),
.B1(n_965),
.B2(n_991),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1050),
.A2(n_874),
.B1(n_890),
.B2(n_857),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1107),
.A2(n_874),
.B1(n_890),
.B2(n_857),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1058),
.A2(n_901),
.B1(n_982),
.B2(n_987),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1059),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1086),
.A2(n_874),
.B1(n_890),
.B2(n_853),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1072),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1091),
.A2(n_987),
.B1(n_982),
.B2(n_902),
.Y(n_1164)
);

AOI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1086),
.A2(n_868),
.B1(n_854),
.B2(n_880),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_1094),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1071),
.A2(n_868),
.B1(n_854),
.B2(n_880),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1084),
.A2(n_868),
.B1(n_854),
.B2(n_880),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1068),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_1047),
.B(n_1076),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1067),
.A2(n_1106),
.B(n_822),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1072),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1085),
.A2(n_868),
.B1(n_854),
.B2(n_880),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1076),
.Y(n_1174)
);

OAI21xp33_ASAP7_75t_L g1175 ( 
.A1(n_1095),
.A2(n_897),
.B(n_904),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1079),
.Y(n_1176)
);

INVxp67_ASAP7_75t_SL g1177 ( 
.A(n_1079),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_1048),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1065),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1128),
.B(n_1088),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1113),
.B(n_1090),
.Y(n_1181)
);

AOI222xp33_ASAP7_75t_L g1182 ( 
.A1(n_1137),
.A2(n_897),
.B1(n_904),
.B2(n_1109),
.C1(n_819),
.C2(n_822),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1136),
.A2(n_892),
.B(n_58),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1116),
.A2(n_1111),
.B1(n_1056),
.B2(n_875),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1113),
.A2(n_854),
.B1(n_868),
.B2(n_880),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_1139),
.A2(n_854),
.B1(n_868),
.B2(n_880),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1138),
.A2(n_892),
.B1(n_875),
.B2(n_1100),
.Y(n_1187)
);

AOI222xp33_ASAP7_75t_L g1188 ( 
.A1(n_1124),
.A2(n_819),
.B1(n_1100),
.B2(n_1095),
.C1(n_814),
.C2(n_812),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1149),
.A2(n_1152),
.B1(n_1117),
.B2(n_1119),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1112),
.A2(n_892),
.B1(n_875),
.B2(n_814),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1122),
.A2(n_875),
.B1(n_812),
.B2(n_965),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1123),
.B(n_1090),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1122),
.A2(n_965),
.B1(n_1087),
.B2(n_1083),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1125),
.Y(n_1194)
);

OAI222xp33_ASAP7_75t_L g1195 ( 
.A1(n_1130),
.A2(n_1105),
.B1(n_1102),
.B2(n_1097),
.C1(n_1065),
.C2(n_1083),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1123),
.B(n_1097),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1171),
.A2(n_1087),
.B1(n_1102),
.B2(n_1105),
.C(n_1096),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_SL g1198 ( 
.A1(n_1127),
.A2(n_1065),
.B1(n_965),
.B2(n_1096),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_L g1199 ( 
.A(n_1158),
.B(n_604),
.C(n_596),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1127),
.A2(n_1096),
.B1(n_900),
.B2(n_987),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1154),
.B(n_982),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1131),
.A2(n_1065),
.B1(n_987),
.B2(n_982),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1147),
.A2(n_956),
.B1(n_953),
.B2(n_918),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1133),
.A2(n_900),
.B1(n_828),
.B2(n_841),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1154),
.B(n_1115),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1175),
.A2(n_900),
.B1(n_828),
.B2(n_841),
.Y(n_1206)
);

NAND3xp33_ASAP7_75t_SL g1207 ( 
.A(n_1169),
.B(n_894),
.C(n_884),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1120),
.A2(n_900),
.B1(n_841),
.B2(n_838),
.Y(n_1208)
);

OAI221xp5_ASAP7_75t_L g1209 ( 
.A1(n_1114),
.A2(n_838),
.B1(n_604),
.B2(n_611),
.C(n_620),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1129),
.A2(n_1169),
.B1(n_1151),
.B2(n_1134),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1153),
.A2(n_1162),
.B(n_1135),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1136),
.A2(n_1142),
.B1(n_1170),
.B2(n_1150),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1115),
.B(n_956),
.Y(n_1213)
);

OAI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1145),
.A2(n_620),
.B(n_611),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1120),
.A2(n_631),
.B1(n_611),
.B2(n_620),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1132),
.A2(n_630),
.B1(n_631),
.B2(n_955),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1146),
.A2(n_953),
.B1(n_951),
.B2(n_952),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1156),
.A2(n_631),
.B1(n_630),
.B2(n_951),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1140),
.A2(n_630),
.B1(n_859),
.B2(n_577),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1148),
.A2(n_577),
.B1(n_59),
.B2(n_60),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1166),
.A2(n_577),
.B1(n_60),
.B2(n_61),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1121),
.A2(n_577),
.B1(n_61),
.B2(n_62),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1118),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_L g1224 ( 
.A1(n_1121),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1173),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1178),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1141),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1178),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1167),
.A2(n_101),
.B1(n_103),
.B2(n_112),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1143),
.A2(n_113),
.B1(n_115),
.B2(n_118),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1144),
.B(n_120),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1164),
.A2(n_121),
.B1(n_122),
.B2(n_128),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1168),
.A2(n_129),
.B1(n_130),
.B2(n_133),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1160),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1144),
.B(n_140),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1161),
.B(n_141),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1155),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1177),
.A2(n_148),
.B(n_149),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1157),
.A2(n_152),
.B1(n_155),
.B2(n_157),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1174),
.B(n_158),
.Y(n_1240)
);

OAI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1174),
.A2(n_159),
.B1(n_163),
.B2(n_165),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1165),
.A2(n_167),
.B1(n_169),
.B2(n_179),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1159),
.A2(n_182),
.B1(n_187),
.B2(n_189),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1176),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1125),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1205),
.B(n_1163),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1205),
.B(n_1192),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1181),
.B(n_1163),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1192),
.B(n_1172),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1212),
.A2(n_1179),
.B1(n_1126),
.B2(n_1172),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1182),
.B(n_1126),
.Y(n_1251)
);

OAI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1226),
.A2(n_1126),
.B1(n_1179),
.B2(n_199),
.C(n_200),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1181),
.B(n_1126),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1240),
.B(n_1179),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1210),
.B(n_1179),
.Y(n_1255)
);

OAI221xp5_ASAP7_75t_SL g1256 ( 
.A1(n_1224),
.A2(n_193),
.B1(n_198),
.B2(n_203),
.C(n_205),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1244),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1196),
.B(n_207),
.Y(n_1258)
);

NAND3xp33_ASAP7_75t_L g1259 ( 
.A(n_1228),
.B(n_209),
.C(n_211),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1196),
.B(n_212),
.Y(n_1260)
);

AND2x2_ASAP7_75t_SL g1261 ( 
.A(n_1186),
.B(n_215),
.Y(n_1261)
);

NOR3xp33_ASAP7_75t_L g1262 ( 
.A(n_1207),
.B(n_218),
.C(n_219),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1201),
.B(n_220),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1201),
.B(n_221),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1189),
.A2(n_222),
.B1(n_223),
.B2(n_225),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1244),
.B(n_226),
.Y(n_1266)
);

AND2x2_ASAP7_75t_SL g1267 ( 
.A(n_1184),
.B(n_227),
.Y(n_1267)
);

OAI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1220),
.A2(n_229),
.B(n_230),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1213),
.B(n_233),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_L g1270 ( 
.A(n_1223),
.B(n_235),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1213),
.B(n_236),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1194),
.B(n_238),
.Y(n_1272)
);

NAND4xp25_ASAP7_75t_L g1273 ( 
.A(n_1215),
.B(n_242),
.C(n_244),
.D(n_245),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1194),
.B(n_251),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1212),
.B(n_253),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1180),
.B(n_1184),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1180),
.B(n_254),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1231),
.B(n_255),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1185),
.B(n_257),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1214),
.A2(n_262),
.B(n_263),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1222),
.A2(n_264),
.B1(n_266),
.B2(n_268),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1188),
.B(n_272),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1235),
.B(n_1236),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1193),
.B(n_1202),
.Y(n_1284)
);

NOR3xp33_ASAP7_75t_L g1285 ( 
.A(n_1183),
.B(n_274),
.C(n_275),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1211),
.B(n_277),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1191),
.B(n_278),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1197),
.A2(n_280),
.B1(n_281),
.B2(n_283),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1221),
.A2(n_284),
.B(n_285),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1217),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1227),
.A2(n_287),
.B1(n_290),
.B2(n_295),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1198),
.B(n_296),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1187),
.B(n_297),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1190),
.B(n_298),
.Y(n_1294)
);

NAND3xp33_ASAP7_75t_L g1295 ( 
.A(n_1262),
.B(n_1225),
.C(n_1238),
.Y(n_1295)
);

AOI221xp5_ASAP7_75t_L g1296 ( 
.A1(n_1275),
.A2(n_1241),
.B1(n_1230),
.B2(n_1209),
.C(n_1218),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1247),
.B(n_1257),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_1285),
.B(n_1234),
.C(n_1245),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1286),
.B(n_1237),
.C(n_1216),
.Y(n_1299)
);

NAND4xp75_ASAP7_75t_L g1300 ( 
.A(n_1267),
.B(n_1239),
.C(n_1195),
.D(n_1232),
.Y(n_1300)
);

AOI221xp5_ASAP7_75t_L g1301 ( 
.A1(n_1268),
.A2(n_1208),
.B1(n_1200),
.B2(n_1203),
.C(n_1229),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1276),
.B(n_1219),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1257),
.B(n_1199),
.Y(n_1303)
);

NAND3xp33_ASAP7_75t_L g1304 ( 
.A(n_1286),
.B(n_1233),
.C(n_1243),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1253),
.B(n_1242),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1248),
.B(n_1204),
.Y(n_1306)
);

AO21x2_ASAP7_75t_L g1307 ( 
.A1(n_1266),
.A2(n_1206),
.B(n_300),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1253),
.B(n_299),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1276),
.B(n_303),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1246),
.B(n_1248),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1259),
.A2(n_328),
.B(n_306),
.Y(n_1311)
);

NOR2x1_ASAP7_75t_L g1312 ( 
.A(n_1280),
.B(n_305),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_1270),
.A2(n_307),
.B1(n_309),
.B2(n_311),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1246),
.B(n_312),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1256),
.B(n_1277),
.C(n_1265),
.Y(n_1315)
);

NAND4xp75_ASAP7_75t_L g1316 ( 
.A(n_1267),
.B(n_313),
.C(n_317),
.D(n_318),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1249),
.B(n_321),
.Y(n_1317)
);

NAND3xp33_ASAP7_75t_L g1318 ( 
.A(n_1277),
.B(n_322),
.C(n_323),
.Y(n_1318)
);

NOR3xp33_ASAP7_75t_L g1319 ( 
.A(n_1268),
.B(n_324),
.C(n_325),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1261),
.A2(n_326),
.B1(n_327),
.B2(n_1270),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1254),
.B(n_1264),
.Y(n_1321)
);

NAND4xp25_ASAP7_75t_L g1322 ( 
.A(n_1283),
.B(n_1255),
.C(n_1251),
.D(n_1291),
.Y(n_1322)
);

AND2x4_ASAP7_75t_SL g1323 ( 
.A(n_1303),
.B(n_1321),
.Y(n_1323)
);

BUFx2_ASAP7_75t_SL g1324 ( 
.A(n_1303),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1297),
.Y(n_1325)
);

HB1xp67_ASAP7_75t_L g1326 ( 
.A(n_1310),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1314),
.Y(n_1327)
);

NAND4xp75_ASAP7_75t_SL g1328 ( 
.A(n_1316),
.B(n_1280),
.C(n_1292),
.D(n_1284),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1312),
.B(n_1284),
.Y(n_1329)
);

BUFx12f_ASAP7_75t_L g1330 ( 
.A(n_1317),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1312),
.B(n_1280),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1314),
.B(n_1290),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1308),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1306),
.Y(n_1334)
);

INVx2_ASAP7_75t_SL g1335 ( 
.A(n_1306),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1305),
.B(n_1280),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1307),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1302),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1322),
.B(n_1290),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1307),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1309),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1318),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1295),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1334),
.Y(n_1344)
);

INVxp67_ASAP7_75t_L g1345 ( 
.A(n_1343),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1334),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1325),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1325),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1338),
.B(n_1250),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1335),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1335),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1335),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1323),
.B(n_1263),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1323),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1342),
.A2(n_1319),
.B1(n_1315),
.B2(n_1320),
.Y(n_1355)
);

INVx2_ASAP7_75t_SL g1356 ( 
.A(n_1323),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1326),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1344),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1354),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1352),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1346),
.Y(n_1361)
);

OA22x2_ASAP7_75t_L g1362 ( 
.A1(n_1355),
.A2(n_1343),
.B1(n_1324),
.B2(n_1329),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1355),
.A2(n_1342),
.B1(n_1329),
.B2(n_1338),
.Y(n_1363)
);

XOR2x2_ASAP7_75t_L g1364 ( 
.A(n_1353),
.B(n_1328),
.Y(n_1364)
);

OA22x2_ASAP7_75t_L g1365 ( 
.A1(n_1345),
.A2(n_1324),
.B1(n_1329),
.B2(n_1336),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1347),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1348),
.Y(n_1367)
);

AO22x2_ASAP7_75t_L g1368 ( 
.A1(n_1345),
.A2(n_1340),
.B1(n_1337),
.B2(n_1331),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1350),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1357),
.Y(n_1370)
);

AOI22x1_ASAP7_75t_L g1371 ( 
.A1(n_1354),
.A2(n_1340),
.B1(n_1337),
.B2(n_1339),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1356),
.A2(n_1300),
.B1(n_1331),
.B2(n_1340),
.Y(n_1372)
);

OA22x2_ASAP7_75t_L g1373 ( 
.A1(n_1351),
.A2(n_1336),
.B1(n_1331),
.B2(n_1326),
.Y(n_1373)
);

OA22x2_ASAP7_75t_L g1374 ( 
.A1(n_1353),
.A2(n_1336),
.B1(n_1341),
.B2(n_1313),
.Y(n_1374)
);

OA22x2_ASAP7_75t_L g1375 ( 
.A1(n_1349),
.A2(n_1341),
.B1(n_1340),
.B2(n_1332),
.Y(n_1375)
);

CKINVDCx16_ASAP7_75t_R g1376 ( 
.A(n_1372),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1364),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1367),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1368),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1367),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1366),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1358),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1361),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1368),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1360),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1370),
.Y(n_1386)
);

NAND4xp25_ASAP7_75t_L g1387 ( 
.A(n_1386),
.B(n_1363),
.C(n_1340),
.D(n_1296),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1376),
.A2(n_1362),
.B1(n_1377),
.B2(n_1374),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1382),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1382),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1378),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1385),
.A2(n_1365),
.B1(n_1359),
.B2(n_1375),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1380),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1381),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1383),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1379),
.A2(n_1373),
.B1(n_1371),
.B2(n_1384),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1389),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1390),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1391),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1393),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1394),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1388),
.A2(n_1371),
.B1(n_1384),
.B2(n_1379),
.C(n_1311),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1395),
.Y(n_1403)
);

AO22x2_ASAP7_75t_L g1404 ( 
.A1(n_1398),
.A2(n_1385),
.B1(n_1396),
.B2(n_1387),
.Y(n_1404)
);

AOI31xp33_ASAP7_75t_L g1405 ( 
.A1(n_1397),
.A2(n_1392),
.A3(n_1339),
.B(n_1299),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1399),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1401),
.B(n_1369),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1403),
.B(n_1339),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1400),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_1402),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1402),
.B(n_1341),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1408),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1407),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1410),
.A2(n_1337),
.B1(n_1330),
.B2(n_1298),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1411),
.B(n_1333),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1406),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1404),
.A2(n_1330),
.B1(n_1327),
.B2(n_1304),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1409),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1413),
.Y(n_1419)
);

NAND4xp25_ASAP7_75t_L g1420 ( 
.A(n_1417),
.B(n_1404),
.C(n_1405),
.D(n_1252),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1414),
.A2(n_1415),
.B1(n_1412),
.B2(n_1418),
.Y(n_1421)
);

NAND4xp25_ASAP7_75t_L g1422 ( 
.A(n_1416),
.B(n_1273),
.C(n_1281),
.D(n_1292),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1417),
.A2(n_1330),
.B1(n_1327),
.B2(n_1282),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1419),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1420),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1421),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1422),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1423),
.Y(n_1428)
);

AO22x2_ASAP7_75t_L g1429 ( 
.A1(n_1421),
.A2(n_1328),
.B1(n_1289),
.B2(n_1288),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1426),
.A2(n_1327),
.B1(n_1333),
.B2(n_1263),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1429),
.A2(n_1333),
.B1(n_1264),
.B2(n_1291),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1429),
.A2(n_1261),
.B1(n_1332),
.B2(n_1271),
.Y(n_1432)
);

AOI211xp5_ASAP7_75t_L g1433 ( 
.A1(n_1424),
.A2(n_1278),
.B(n_1287),
.C(n_1269),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1430),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1433),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1432),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1431),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1434),
.A2(n_1428),
.B1(n_1425),
.B2(n_1427),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1437),
.A2(n_1332),
.B1(n_1260),
.B2(n_1258),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1436),
.A2(n_1435),
.B1(n_1332),
.B2(n_1287),
.Y(n_1440)
);

INVxp67_ASAP7_75t_L g1441 ( 
.A(n_1438),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1440),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1441),
.A2(n_1439),
.B1(n_1332),
.B2(n_1279),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1443),
.Y(n_1444)
);

AOI221x1_ASAP7_75t_L g1445 ( 
.A1(n_1444),
.A2(n_1442),
.B1(n_1272),
.B2(n_1274),
.C(n_1293),
.Y(n_1445)
);

AOI211xp5_ASAP7_75t_L g1446 ( 
.A1(n_1445),
.A2(n_1279),
.B(n_1294),
.C(n_1301),
.Y(n_1446)
);


endmodule