module fake_jpeg_24098_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_31),
.B(n_20),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2x1_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_20),
.B1(n_18),
.B2(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_15),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_23),
.B1(n_30),
.B2(n_25),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_20),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_17),
.B1(n_30),
.B2(n_18),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_32),
.B(n_29),
.C(n_30),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_32),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_21),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_68),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_67),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_38),
.B1(n_34),
.B2(n_41),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_65),
.A2(n_66),
.B1(n_48),
.B2(n_42),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_70),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_32),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_75),
.B(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_19),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_54),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_32),
.B(n_29),
.C(n_40),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_52),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_90),
.B(n_97),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_47),
.B1(n_42),
.B2(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_88),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_76),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_91),
.B(n_94),
.Y(n_120)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_93),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_98),
.A2(n_72),
.B1(n_28),
.B2(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_58),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_77),
.B(n_80),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_106),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_107),
.B(n_76),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_73),
.C(n_74),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_112),
.C(n_115),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_72),
.B1(n_87),
.B2(n_98),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_83),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_100),
.B1(n_88),
.B2(n_82),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_44),
.C(n_78),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_44),
.C(n_80),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_66),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_118),
.B(n_64),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_76),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_87),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_75),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_124),
.B1(n_137),
.B2(n_102),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_101),
.B1(n_100),
.B2(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_126),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_133),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_129),
.B1(n_106),
.B2(n_112),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_81),
.B1(n_89),
.B2(n_45),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_132),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_89),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_81),
.B(n_70),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_140),
.B(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_47),
.B1(n_55),
.B2(n_99),
.Y(n_137)
);

AOI22x1_ASAP7_75t_SL g139 ( 
.A1(n_122),
.A2(n_70),
.B1(n_58),
.B2(n_43),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_36),
.B1(n_61),
.B2(n_48),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_91),
.B(n_84),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_92),
.A3(n_43),
.B1(n_83),
.B2(n_40),
.C1(n_36),
.C2(n_55),
.Y(n_141)
);

OAI322xp33_ASAP7_75t_L g152 ( 
.A1(n_141),
.A2(n_130),
.A3(n_139),
.B1(n_136),
.B2(n_121),
.C1(n_140),
.C2(n_127),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_157),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_119),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_138),
.C(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_151),
.B1(n_136),
.B2(n_123),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_155),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_129),
.A2(n_117),
.B1(n_120),
.B2(n_102),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_154),
.B1(n_158),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_109),
.B1(n_103),
.B2(n_113),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_155),
.A3(n_156),
.B1(n_144),
.B2(n_160),
.C1(n_145),
.C2(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_153),
.Y(n_170)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_158),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_61),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_168),
.B1(n_169),
.B2(n_174),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_166),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_138),
.Y(n_163)
);

OA21x2_ASAP7_75t_SL g177 ( 
.A1(n_163),
.A2(n_165),
.B(n_27),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_43),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_40),
.C(n_21),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_24),
.C(n_19),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_29),
.B1(n_21),
.B2(n_14),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_1),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_27),
.B1(n_24),
.B2(n_19),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_162),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_177),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_27),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_179),
.C(n_187),
.Y(n_193)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_175),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_188),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_1),
.B(n_2),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_186),
.B1(n_7),
.B2(n_8),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_168),
.A2(n_170),
.B1(n_167),
.B2(n_169),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_27),
.Y(n_187)
);

NOR3xp33_ASAP7_75t_SL g188 ( 
.A(n_172),
.B(n_3),
.C(n_5),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_174),
.B(n_6),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_193),
.B(n_11),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_186),
.B(n_3),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_197),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_27),
.C(n_24),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_19),
.C(n_24),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_196),
.Y(n_204)
);

OAI221xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_188),
.B1(n_176),
.B2(n_180),
.C(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_199),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

OAI221xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_203),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_194),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_205),
.B(n_11),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_9),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_202),
.A2(n_189),
.B1(n_200),
.B2(n_196),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_12),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_12),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_12),
.C(n_13),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_213),
.A2(n_215),
.B(n_208),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_214),
.A2(n_216),
.B(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_19),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_214),
.A2(n_212),
.B(n_13),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_221),
.A2(n_24),
.B(n_27),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_220),
.Y(n_223)
);


endmodule