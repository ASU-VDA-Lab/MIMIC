module fake_jpeg_2553_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_8),
.B(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_44),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_30),
.B1(n_40),
.B2(n_36),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_55),
.B1(n_45),
.B2(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_37),
.B1(n_31),
.B2(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

AOI222xp33_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_44),
.B1(n_47),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_66),
.B1(n_54),
.B2(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_0),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_1),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_65),
.C(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_46),
.B1(n_3),
.B2(n_6),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_57),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_21),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_75),
.Y(n_83)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_47),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_56),
.B1(n_7),
.B2(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_1),
.B1(n_7),
.B2(n_9),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_86),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_88),
.B(n_10),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_15),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_22),
.B1(n_11),
.B2(n_14),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_90),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_SL g90 ( 
.A1(n_88),
.A2(n_76),
.A3(n_68),
.B1(n_10),
.B2(n_77),
.C1(n_24),
.C2(n_25),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_81),
.B1(n_85),
.B2(n_27),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_97),
.C(n_91),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_92),
.C(n_96),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_98),
.Y(n_101)
);

OAI21x1_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_93),
.B(n_85),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_17),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_19),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_28),
.CI(n_29),
.CON(n_106),
.SN(n_106)
);


endmodule