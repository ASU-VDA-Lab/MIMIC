module fake_jpeg_573_n_205 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_205);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_7),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_49),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_51),
.Y(n_87)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_71),
.B1(n_58),
.B2(n_73),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_94),
.B1(n_71),
.B2(n_67),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_72),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_72),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_68),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_70),
.B1(n_73),
.B2(n_57),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_98),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_95),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_112),
.Y(n_127)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_78),
.B1(n_66),
.B2(n_71),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_106),
.B1(n_56),
.B2(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_52),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_107),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_95),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_111),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_23),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_92),
.B(n_65),
.Y(n_111)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_62),
.Y(n_123)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_121),
.A2(n_53),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_132),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_106),
.A2(n_61),
.B1(n_55),
.B2(n_56),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_130),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_103),
.B1(n_98),
.B2(n_114),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_60),
.B1(n_63),
.B2(n_53),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_74),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_0),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_0),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_136),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_143),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_63),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_151),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_126),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_146),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_152),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_1),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_11),
.B(n_13),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_1),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_150),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_53),
.C(n_26),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_153),
.B(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_157),
.Y(n_160)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_28),
.C(n_45),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_122),
.C(n_34),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_13),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_162),
.B(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_169),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_36),
.C(n_43),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_173),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_14),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_30),
.B(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_171),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_172),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_24),
.C(n_40),
.Y(n_173)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_147),
.B(n_159),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_168),
.B(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_150),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_174),
.A2(n_151),
.B1(n_158),
.B2(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_163),
.B1(n_167),
.B2(n_161),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_193),
.B(n_183),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g188 ( 
.A(n_177),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_190),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_170),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_175),
.C(n_168),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_191),
.B(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_195),
.A2(n_196),
.B1(n_189),
.B2(n_181),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_192),
.C(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_199),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_179),
.B(n_194),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_180),
.C(n_186),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_22),
.A3(n_39),
.B1(n_17),
.B2(n_19),
.C1(n_21),
.C2(n_41),
.Y(n_203)
);

AOI211xp5_ASAP7_75t_SL g204 ( 
.A1(n_203),
.A2(n_37),
.B(n_38),
.C(n_14),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_204),
.B(n_16),
.Y(n_205)
);


endmodule