module real_jpeg_316_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_1),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_1),
.A2(n_36),
.B1(n_59),
.B2(n_61),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_46),
.B1(n_59),
.B2(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_2),
.A2(n_29),
.B1(n_35),
.B2(n_46),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_2),
.A2(n_46),
.B1(n_73),
.B2(n_74),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_29),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_5),
.A2(n_73),
.B1(n_74),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_5),
.A2(n_59),
.B1(n_61),
.B2(n_81),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_81),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_5),
.A2(n_29),
.B1(n_35),
.B2(n_81),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_6),
.A2(n_73),
.B1(n_74),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_59),
.B1(n_61),
.B2(n_83),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_83),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_83),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_73),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_7),
.B(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_7),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_73),
.B(n_136),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_7),
.B(n_63),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g205 ( 
.A1(n_7),
.A2(n_61),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_7),
.B(n_29),
.C(n_49),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_7),
.B(n_32),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_7),
.B(n_54),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_12),
.A2(n_53),
.B1(n_59),
.B2(n_61),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_12),
.A2(n_29),
.B1(n_35),
.B2(n_53),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_13),
.A2(n_73),
.B1(n_74),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_13),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_13),
.A2(n_59),
.B1(n_61),
.B2(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_13),
.A2(n_43),
.B1(n_44),
.B2(n_126),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_13),
.A2(n_29),
.B1(n_35),
.B2(n_126),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_73),
.B1(n_74),
.B2(n_146),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_14),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_59),
.B1(n_61),
.B2(n_146),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_146),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_14),
.A2(n_29),
.B1(n_35),
.B2(n_146),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_15),
.A2(n_43),
.B1(n_44),
.B2(n_58),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_15),
.A2(n_29),
.B1(n_35),
.B2(n_58),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_264),
.B1(n_286),
.B2(n_287),
.Y(n_19)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_20),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_128),
.B(n_263),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_110),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_22),
.B(n_110),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_84),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_23),
.B(n_94),
.C(n_109),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_55),
.C(n_69),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_24),
.A2(n_25),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_39),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_26),
.A2(n_27),
.B1(n_39),
.B2(n_40),
.Y(n_148)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_28),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_28),
.A2(n_32),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_28),
.A2(n_32),
.B1(n_139),
.B2(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_28),
.A2(n_32),
.B1(n_176),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_28),
.A2(n_32),
.B1(n_172),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_28),
.A2(n_32),
.B1(n_226),
.B2(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_29),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_29),
.B(n_224),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_31),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_31),
.A2(n_34),
.B1(n_98),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_31),
.A2(n_98),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_31),
.A2(n_98),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_42),
.A2(n_51),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_44),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_43),
.B(n_65),
.Y(n_173)
);

INVx5_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_44),
.A2(n_61),
.A3(n_64),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_44),
.B(n_214),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_54),
.B1(n_91),
.B2(n_92),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_91),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_47),
.A2(n_54),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_47),
.A2(n_54),
.B1(n_168),
.B2(n_188),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_47),
.A2(n_54),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_47),
.A2(n_54),
.B1(n_196),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_47),
.A2(n_54),
.B(n_92),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_51),
.A2(n_119),
.B1(n_167),
.B2(n_208),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_69),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_67),
.B2(n_68),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_57),
.A2(n_63),
.B1(n_88),
.B2(n_123),
.Y(n_122)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_65),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_61),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_59),
.B(n_76),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_59),
.B(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g135 ( 
.A1(n_61),
.A2(n_74),
.A3(n_77),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_62),
.A2(n_68),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_62),
.A2(n_68),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_62),
.A2(n_68),
.B1(n_142),
.B2(n_158),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_62),
.A2(n_68),
.B1(n_157),
.B2(n_205),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_63),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_63),
.A2(n_88),
.B1(n_89),
.B2(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_78),
.B1(n_79),
.B2(n_82),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_78),
.B1(n_82),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_70),
.A2(n_78),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_70),
.A2(n_78),
.B1(n_145),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_70),
.A2(n_78),
.B1(n_107),
.B2(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_80),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_78),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_94),
.B1(n_95),
.B2(n_109),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B(n_93),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_90),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_93),
.A2(n_270),
.B1(n_282),
.B2(n_283),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_93),
.Y(n_282)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_102),
.B1(n_103),
.B2(n_108),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_114)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_104),
.A2(n_106),
.B(n_108),
.Y(n_268)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.C(n_115),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.C(n_124),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_117),
.B(n_120),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_118),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_124),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_123),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_151),
.B(n_262),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_149),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_130),
.B(n_149),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_148),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_131),
.B(n_148),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_133),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_141),
.C(n_144),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_134),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_138),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_141),
.B(n_144),
.Y(n_252)
);

AOI31xp33_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_246),
.A3(n_255),
.B(n_259),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_191),
.B(n_245),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_178),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_154),
.B(n_178),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_165),
.C(n_169),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_155),
.B(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_160),
.C(n_164),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_164),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_162),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_165),
.B(n_169),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_174),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_171),
.Y(n_206)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_183),
.B(n_186),
.C(n_190),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_187),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_240),
.B(n_244),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_209),
.B(n_239),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_201),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_198),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_200),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_204),
.C(n_207),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_220),
.B(n_238),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_218),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_215),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_232),
.B(n_237),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_231),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_243),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_250),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_254),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_285),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_284),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_284),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_281),
.Y(n_275)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);


endmodule