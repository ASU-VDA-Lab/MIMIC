module real_jpeg_25972_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_1),
.A2(n_21),
.B1(n_26),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_1),
.A2(n_23),
.B1(n_30),
.B2(n_51),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_128)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_75),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_23),
.B1(n_27),
.B2(n_30),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_2),
.B(n_35),
.C(n_57),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_2),
.B(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_2),
.A2(n_32),
.B1(n_121),
.B2(n_128),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_3),
.A2(n_34),
.B1(n_35),
.B2(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_3),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_6),
.A2(n_23),
.B1(n_30),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_6),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_63),
.Y(n_111)
);

INVx8_ASAP7_75t_SL g78 ( 
.A(n_7),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_8),
.A2(n_23),
.B1(n_30),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_8),
.A2(n_21),
.B1(n_26),
.B2(n_54),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_9),
.A2(n_34),
.B1(n_35),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_23),
.B1(n_30),
.B2(n_40),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_94),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_64),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_18),
.B(n_64),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_46),
.C(n_52),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_19),
.B(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_20),
.B(n_31),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.A3(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_20)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_21),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_21),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_21),
.A2(n_26),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

AO22x1_ASAP7_75t_L g49 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g56 ( 
.A1(n_23),
.A2(n_30),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_23),
.B(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_27),
.CON(n_25),
.SN(n_25)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_27),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_27),
.B(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_38),
.B(n_41),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_32),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_32),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_33),
.B(n_42),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_33),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_34),
.A2(n_35),
.B1(n_57),
.B2(n_59),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_34),
.B(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_37),
.Y(n_130)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_39),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g113 ( 
.A(n_45),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_46),
.B(n_52),
.Y(n_141)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_55),
.B1(n_61),
.B2(n_101),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_62),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_61),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_85),
.B2(n_86),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_87),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_138),
.B(n_142),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_114),
.B(n_137),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_102),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_110),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_109),
.C(n_110),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_124),
.B(n_136),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_123),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_123),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_131),
.B(n_135),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_126),
.B(n_127),
.Y(n_135)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_139),
.B(n_140),
.Y(n_142)
);


endmodule