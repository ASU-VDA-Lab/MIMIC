module fake_jpeg_3025_n_80 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx4_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_2),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_28),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_10),
.B(n_9),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx24_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

CKINVDCx12_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_27),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_48),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_44),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_23),
.B(n_29),
.C(n_24),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_15),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_14),
.B1(n_20),
.B2(n_21),
.Y(n_50)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_9),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_54),
.A2(n_46),
.B1(n_42),
.B2(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_20),
.B1(n_25),
.B2(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_55),
.B1(n_60),
.B2(n_53),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_66),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_51),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_66),
.C(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_67),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_1),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_74),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_55),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_33),
.Y(n_80)
);


endmodule