module fake_netlist_1_7853_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2xp33_ASAP7_75t_L g11 ( .A(n_2), .B(n_9), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_6), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_10), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
AOI21x1_ASAP7_75t_L g16 ( .A1(n_1), .A2(n_7), .B(n_0), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_4), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_16), .B(n_1), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_15), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_12), .B(n_2), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_13), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_22), .B(n_14), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_18), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_21), .Y(n_27) );
OAI21xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_25), .B(n_21), .Y(n_28) );
AOI211x1_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_19), .B(n_3), .C(n_27), .Y(n_29) );
CKINVDCx5p33_ASAP7_75t_R g30 ( .A(n_29), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
OAI22x1_ASAP7_75t_SL g32 ( .A1(n_30), .A2(n_3), .B1(n_11), .B2(n_8), .Y(n_32) );
AOI22xp5_ASAP7_75t_SL g33 ( .A1(n_32), .A2(n_31), .B1(n_5), .B2(n_25), .Y(n_33) );
endmodule