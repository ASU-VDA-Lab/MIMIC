module fake_jpeg_28776_n_180 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_55),
.B(n_50),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_81),
.B(n_55),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_51),
.B1(n_48),
.B2(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_80),
.B1(n_50),
.B2(n_48),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_95),
.B(n_88),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_56),
.B1(n_51),
.B2(n_62),
.Y(n_95)
);

NAND2x1p5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_49),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_116),
.Y(n_119)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_57),
.B1(n_70),
.B2(n_69),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_101),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

BUFx2_ASAP7_75t_SL g108 ( 
.A(n_85),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_108),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_85),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_85),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_2),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_109),
.A2(n_59),
.B1(n_66),
.B2(n_68),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_123),
.B1(n_133),
.B2(n_139),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_67),
.B1(n_65),
.B2(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_60),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_136),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_58),
.B(n_49),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_8),
.B(n_9),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_6),
.B(n_7),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_1),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_98),
.B1(n_110),
.B2(n_4),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_2),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_134),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_23),
.A3(n_45),
.B1(n_43),
.B2(n_42),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_138),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_3),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_155),
.B1(n_157),
.B2(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_148),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_25),
.C(n_40),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_156),
.C(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_10),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_150),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_152),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_16),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_17),
.B1(n_19),
.B2(n_21),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_158),
.B(n_159),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_130),
.C(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_160),
.A2(n_143),
.B1(n_156),
.B2(n_154),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_164),
.C(n_166),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_161),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_167),
.B1(n_141),
.B2(n_165),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_165),
.C(n_168),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_140),
.B(n_154),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_153),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_122),
.C(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_24),
.C(n_26),
.Y(n_180)
);


endmodule