module fake_ariane_3176_n_1905 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1905);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1905;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_189),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_57),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_63),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_30),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_8),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_50),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_7),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_42),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_182),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_77),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_33),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_42),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_27),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_178),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_117),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_3),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_35),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_66),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_64),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_144),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_175),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_62),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_170),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_106),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_114),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_97),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_58),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_40),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_181),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_103),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_123),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_132),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_16),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_120),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_12),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_136),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_19),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_78),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_177),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_143),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_20),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_67),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_179),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_184),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_171),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_160),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_89),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_79),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_57),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_118),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_161),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_74),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_1),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_72),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_167),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_44),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_83),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_17),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_180),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_109),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_107),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_166),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_38),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_32),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_75),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_157),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_141),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_5),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_146),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_48),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_125),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_59),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_88),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_127),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_59),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_99),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_31),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_90),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_137),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_23),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_14),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_50),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_54),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_29),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_190),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_93),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_95),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_55),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_149),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_41),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_194),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_12),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_11),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_108),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_85),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_94),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_8),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_145),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_40),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_119),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_68),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_48),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_140),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_27),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_150),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_26),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_3),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_168),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_173),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_4),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_165),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_5),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_82),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_115),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_49),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_159),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_53),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_188),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_193),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_29),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_101),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_37),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_34),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_26),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_152),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_148),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_153),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_71),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_135),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_164),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_169),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_110),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_76),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_102),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_21),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_61),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_13),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_4),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_172),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_37),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_126),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_38),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_163),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_121),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_6),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_113),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_56),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_61),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_18),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_55),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_34),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_116),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_65),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_19),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_186),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_21),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_6),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_41),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_56),
.Y(n_379)
);

BUFx10_ASAP7_75t_L g380 ( 
.A(n_0),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_22),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_69),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_28),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_28),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_11),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_33),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_7),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_47),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_124),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_122),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_73),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_133),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_52),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_206),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_384),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_206),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_347),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_220),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_312),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_244),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_225),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_280),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_280),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_300),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_237),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_300),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_360),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_369),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_387),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_209),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_387),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_238),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_266),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_215),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_215),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_246),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_246),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_248),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_297),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_297),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_317),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_317),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVxp67_ASAP7_75t_SL g426 ( 
.A(n_281),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_363),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_268),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_287),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_294),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_295),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_303),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_241),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_265),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_307),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_292),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_316),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_266),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_318),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_266),
.Y(n_440)
);

INVxp33_ASAP7_75t_SL g441 ( 
.A(n_224),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g442 ( 
.A(n_376),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_202),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_199),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_279),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_202),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_329),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_234),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_201),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_199),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_340),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_234),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_358),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_201),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_200),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_204),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_207),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_200),
.Y(n_460)
);

INVxp33_ASAP7_75t_SL g461 ( 
.A(n_207),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_383),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_201),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_299),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_352),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_205),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_228),
.Y(n_467)
);

CKINVDCx14_ASAP7_75t_R g468 ( 
.A(n_304),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_299),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_299),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_365),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

INVx2_ASAP7_75t_SL g475 ( 
.A(n_380),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_308),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_232),
.Y(n_477)
);

INVxp33_ASAP7_75t_SL g478 ( 
.A(n_210),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_233),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_243),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_345),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_245),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_210),
.Y(n_483)
);

INVxp33_ASAP7_75t_SL g484 ( 
.A(n_212),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_372),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_203),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_247),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_249),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_250),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_255),
.Y(n_490)
);

INVxp33_ASAP7_75t_SL g491 ( 
.A(n_212),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_259),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_412),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_416),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_416),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_485),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_372),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_485),
.B(n_346),
.Y(n_498)
);

NOR2x1_ASAP7_75t_L g499 ( 
.A(n_448),
.B(n_291),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_441),
.A2(n_355),
.B1(n_357),
.B2(n_367),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_442),
.A2(n_377),
.B1(n_325),
.B2(n_302),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_448),
.B(n_372),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_417),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_452),
.B(n_261),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_417),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_346),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_414),
.A2(n_337),
.B1(n_388),
.B2(n_386),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_418),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_419),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_419),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_394),
.B(n_213),
.Y(n_513)
);

OA21x2_ASAP7_75t_L g514 ( 
.A1(n_421),
.A2(n_264),
.B(n_262),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_452),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_433),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_422),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_434),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_269),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_466),
.B(n_270),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_457),
.Y(n_527)
);

BUFx2_ASAP7_75t_L g528 ( 
.A(n_395),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_405),
.A2(n_393),
.B1(n_273),
.B2(n_211),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_425),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_479),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_425),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_468),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_445),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_277),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_476),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_457),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_480),
.B(n_278),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_482),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_481),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_467),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_467),
.B(n_282),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_487),
.B(n_306),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_488),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_401),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_488),
.B(n_322),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_492),
.B(n_336),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_399),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_489),
.B(n_490),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_490),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_429),
.A2(n_349),
.B(n_348),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_396),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_403),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_403),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_404),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

INVxp33_ASAP7_75t_L g562 ( 
.A(n_446),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_402),
.B(n_350),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_406),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_406),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_395),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_407),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_464),
.B(n_353),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_407),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_408),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_408),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_519),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_529),
.A2(n_405),
.B1(n_221),
.B2(n_235),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_502),
.B(n_506),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_519),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_552),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_R g578 ( 
.A(n_534),
.B(n_465),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_562),
.B(n_397),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_519),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_502),
.B(n_415),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_507),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_566),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_507),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_519),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_519),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_519),
.Y(n_588)
);

NAND2xp33_ASAP7_75t_L g589 ( 
.A(n_497),
.B(n_444),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_506),
.B(n_415),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_496),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_496),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_520),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_520),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_506),
.B(n_438),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_520),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g597 ( 
.A(n_500),
.B(n_438),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_547),
.B(n_450),
.C(n_444),
.Y(n_598)
);

NOR3xp33_ASAP7_75t_L g599 ( 
.A(n_508),
.B(n_370),
.C(n_450),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_520),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_549),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_520),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_520),
.Y(n_603)
);

AND2x6_ASAP7_75t_L g604 ( 
.A(n_499),
.B(n_375),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_520),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_566),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_566),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_497),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_566),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_515),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_513),
.B(n_397),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_506),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_513),
.B(n_455),
.Y(n_615)
);

OAI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_529),
.A2(n_461),
.B1(n_478),
.B2(n_443),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_569),
.B(n_475),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_496),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_541),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_547),
.B(n_440),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_566),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_547),
.B(n_440),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_515),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_503),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_503),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_541),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_541),
.Y(n_628)
);

NAND3xp33_ASAP7_75t_L g629 ( 
.A(n_547),
.B(n_486),
.C(n_460),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_564),
.B(n_460),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_503),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

INVx5_ASAP7_75t_L g633 ( 
.A(n_497),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_543),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_515),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_554),
.B(n_498),
.Y(n_636)
);

OAI22x1_ASAP7_75t_L g637 ( 
.A1(n_500),
.A2(n_428),
.B1(n_436),
.B2(n_454),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_543),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_554),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_505),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_554),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_505),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_497),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_554),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_505),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_511),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_564),
.B(n_486),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_511),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_511),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_498),
.B(n_475),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_569),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_497),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_524),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_497),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_498),
.B(n_469),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_524),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_524),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_561),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_525),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_525),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_525),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_563),
.A2(n_491),
.B1(n_484),
.B2(n_335),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_532),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_497),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_497),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_532),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_531),
.B(n_449),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_526),
.A2(n_459),
.B1(n_439),
.B2(n_453),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_499),
.B(n_470),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_532),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_533),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_498),
.B(n_472),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_544),
.B(n_411),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_533),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_497),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_531),
.B(n_471),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_526),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_533),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_535),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_531),
.B(n_473),
.Y(n_680)
);

BUFx2_ASAP7_75t_L g681 ( 
.A(n_528),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_535),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_535),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_557),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_526),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_544),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_548),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_536),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_548),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_557),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_555),
.Y(n_691)
);

AO21x2_ASAP7_75t_L g692 ( 
.A1(n_556),
.A2(n_474),
.B(n_426),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_558),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_555),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_526),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_558),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_558),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_569),
.B(n_420),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_R g699 ( 
.A(n_567),
.B(n_398),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_494),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_495),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_569),
.B(n_429),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_560),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_560),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_560),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_545),
.B(n_203),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_495),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_568),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_509),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_508),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_509),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_568),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_545),
.B(n_208),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_510),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_510),
.Y(n_715)
);

NAND2xp33_ASAP7_75t_L g716 ( 
.A(n_553),
.B(n_208),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_512),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_545),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_545),
.B(n_430),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_568),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_514),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_639),
.Y(n_722)
);

AND2x6_ASAP7_75t_SL g723 ( 
.A(n_580),
.B(n_537),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_635),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_610),
.B(n_546),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_639),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_630),
.A2(n_546),
.B1(n_550),
.B2(n_537),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_647),
.B(n_546),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_614),
.B(n_677),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_641),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_615),
.B(n_557),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_635),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_635),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_612),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_624),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_710),
.A2(n_514),
.B1(n_546),
.B2(n_550),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_598),
.B(n_550),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_614),
.B(n_550),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_644),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_681),
.B(n_501),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_721),
.A2(n_514),
.B1(n_539),
.B2(n_512),
.Y(n_741)
);

OAI22xp33_ASAP7_75t_L g742 ( 
.A1(n_574),
.A2(n_501),
.B1(n_553),
.B2(n_523),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_681),
.Y(n_743)
);

OAI22x1_ASAP7_75t_SL g744 ( 
.A1(n_688),
.A2(n_493),
.B1(n_516),
.B2(n_521),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_677),
.B(n_527),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_612),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_610),
.Y(n_747)
);

A2O1A1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_698),
.A2(n_556),
.B(n_523),
.C(n_540),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_721),
.A2(n_514),
.B1(n_539),
.B2(n_518),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_652),
.B(n_517),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_685),
.B(n_527),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_685),
.B(n_695),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_610),
.B(n_556),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_610),
.Y(n_754)
);

CKINVDCx11_ASAP7_75t_R g755 ( 
.A(n_577),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_718),
.B(n_527),
.Y(n_756)
);

AO22x2_ASAP7_75t_L g757 ( 
.A1(n_599),
.A2(n_540),
.B1(n_551),
.B2(n_522),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_583),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_683),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_683),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_718),
.B(n_551),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_575),
.B(n_561),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_652),
.B(n_214),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_702),
.B(n_582),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_644),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_702),
.B(n_561),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_683),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_598),
.B(n_504),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_652),
.B(n_214),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_636),
.A2(n_572),
.B(n_571),
.C(n_561),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_684),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_664),
.B(n_216),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_686),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_L g774 ( 
.A(n_658),
.B(n_620),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_702),
.B(n_565),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_664),
.B(n_216),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_624),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_613),
.B(n_236),
.C(n_219),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_702),
.B(n_673),
.Y(n_779)
);

BUFx4f_ASAP7_75t_L g780 ( 
.A(n_669),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_601),
.B(n_565),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_664),
.B(n_217),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_673),
.B(n_565),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_623),
.B(n_565),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_667),
.B(n_571),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_629),
.B(n_504),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_624),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_676),
.B(n_571),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_688),
.Y(n_789)
);

AO22x1_ASAP7_75t_L g790 ( 
.A1(n_617),
.A2(n_662),
.B1(n_583),
.B2(n_585),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_617),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_719),
.B(n_571),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_680),
.B(n_572),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_687),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_665),
.B(n_217),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_574),
.B(n_538),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_665),
.B(n_218),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_629),
.A2(n_517),
.B1(n_530),
.B2(n_522),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_590),
.B(n_572),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_624),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_665),
.B(n_218),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_595),
.B(n_572),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_617),
.A2(n_518),
.B1(n_530),
.B2(n_227),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_577),
.Y(n_804)
);

NAND2x1_ASAP7_75t_L g805 ( 
.A(n_675),
.B(n_514),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_617),
.A2(n_223),
.B1(n_240),
.B2(n_392),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_689),
.B(n_559),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_658),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_591),
.A2(n_559),
.B(n_570),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_675),
.B(n_222),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_689),
.B(n_691),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_675),
.B(n_222),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_694),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_694),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_668),
.B(n_542),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_669),
.B(n_570),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_651),
.B(n_223),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_625),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_578),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_SL g820 ( 
.A(n_699),
.B(n_219),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_626),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_669),
.B(n_310),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_651),
.B(n_226),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_631),
.Y(n_824)
);

OAI22xp33_ASAP7_75t_L g825 ( 
.A1(n_655),
.A2(n_344),
.B1(n_242),
.B2(n_236),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_669),
.B(n_314),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_650),
.A2(n_344),
.B1(n_242),
.B2(n_335),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_706),
.B(n_253),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_597),
.Y(n_829)
);

BUFx8_ASAP7_75t_L g830 ( 
.A(n_669),
.Y(n_830)
);

NOR3xp33_ASAP7_75t_L g831 ( 
.A(n_616),
.B(n_343),
.C(n_342),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_591),
.B(n_339),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_669),
.B(n_226),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_713),
.B(n_263),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_672),
.A2(n_388),
.B1(n_342),
.B2(n_343),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_651),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_597),
.B(n_400),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_700),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_701),
.B(n_229),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_684),
.B(n_271),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_701),
.B(n_229),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_707),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_707),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_684),
.B(n_274),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_709),
.B(n_230),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_709),
.B(n_230),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_711),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_651),
.B(n_643),
.Y(n_848)
);

NAND2x1p5_ASAP7_75t_L g849 ( 
.A(n_690),
.B(n_409),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_711),
.B(n_231),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_640),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_640),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_714),
.B(n_231),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_714),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_715),
.A2(n_432),
.B(n_430),
.C(n_431),
.Y(n_855)
);

INVx8_ASAP7_75t_L g856 ( 
.A(n_633),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_643),
.B(n_239),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_721),
.A2(n_462),
.B1(n_458),
.B2(n_456),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_690),
.B(n_285),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_642),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_715),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_717),
.Y(n_862)
);

AO22x2_ASAP7_75t_L g863 ( 
.A1(n_616),
.A2(n_431),
.B1(n_432),
.B2(n_447),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_637),
.B(n_435),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_648),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_648),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_717),
.A2(n_362),
.B1(n_385),
.B2(n_386),
.Y(n_867)
);

BUFx5_ASAP7_75t_L g868 ( 
.A(n_592),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_604),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_589),
.A2(n_240),
.B1(n_392),
.B2(n_391),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_690),
.B(n_289),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_592),
.B(n_239),
.Y(n_872)
);

NAND2xp33_ASAP7_75t_L g873 ( 
.A(n_658),
.B(n_334),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_637),
.B(n_437),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_607),
.B(n_298),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_658),
.B(n_451),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_607),
.B(n_618),
.Y(n_877)
);

INVx1_ASAP7_75t_SL g878 ( 
.A(n_804),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_768),
.B(n_618),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_SL g880 ( 
.A(n_778),
.B(n_385),
.C(n_362),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_789),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_742),
.A2(n_837),
.B1(n_796),
.B2(n_820),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_856),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_818),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_735),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_742),
.A2(n_604),
.B1(n_721),
.B2(n_696),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_768),
.B(n_645),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_773),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_727),
.A2(n_658),
.B1(n_645),
.B2(n_646),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_791),
.B(n_633),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_764),
.B(n_633),
.Y(n_891)
);

AND2x4_ASAP7_75t_SL g892 ( 
.A(n_819),
.B(n_646),
.Y(n_892)
);

AO22x1_ASAP7_75t_L g893 ( 
.A1(n_829),
.A2(n_604),
.B1(n_331),
.B2(n_309),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_811),
.A2(n_593),
.B(n_587),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_755),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_737),
.A2(n_716),
.B1(n_604),
.B2(n_653),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_794),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_737),
.A2(n_604),
.B1(n_653),
.B2(n_670),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_786),
.B(n_656),
.Y(n_899)
);

INVx5_ASAP7_75t_L g900 ( 
.A(n_856),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_736),
.A2(n_604),
.B1(n_712),
.B2(n_708),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_736),
.A2(n_604),
.B1(n_712),
.B2(n_708),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_815),
.A2(n_720),
.B1(n_705),
.B2(n_704),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_813),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_814),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_SL g906 ( 
.A1(n_743),
.A2(n_326),
.B1(n_301),
.B2(n_311),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_784),
.A2(n_593),
.B(n_587),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_744),
.Y(n_908)
);

NAND2xp33_ASAP7_75t_SL g909 ( 
.A(n_728),
.B(n_587),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_779),
.B(n_656),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_758),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_786),
.B(n_659),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_838),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_781),
.B(n_633),
.Y(n_914)
);

INVx1_ASAP7_75t_SL g915 ( 
.A(n_740),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_842),
.B(n_659),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_832),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_843),
.B(n_660),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_832),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_SL g920 ( 
.A(n_831),
.B(n_323),
.C(n_321),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_723),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_847),
.Y(n_922)
);

INVxp67_ASAP7_75t_SL g923 ( 
.A(n_771),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_821),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_854),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_824),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_864),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_861),
.B(n_660),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_SL g929 ( 
.A(n_831),
.B(n_356),
.C(n_332),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_862),
.B(n_661),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_722),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_863),
.A2(n_720),
.B1(n_705),
.B2(n_704),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_726),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_874),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_761),
.B(n_661),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_R g936 ( 
.A(n_830),
.B(n_593),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_730),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_790),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_762),
.B(n_670),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_757),
.A2(n_679),
.B1(n_678),
.B2(n_682),
.Y(n_940)
);

INVxp67_ASAP7_75t_SL g941 ( 
.A(n_771),
.Y(n_941)
);

BUFx12f_ASAP7_75t_L g942 ( 
.A(n_830),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_739),
.Y(n_943)
);

INVxp67_ASAP7_75t_SL g944 ( 
.A(n_752),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_856),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_731),
.B(n_678),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_836),
.B(n_633),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_851),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_869),
.B(n_633),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_765),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_799),
.B(n_679),
.Y(n_951)
);

INVx2_ASAP7_75t_SL g952 ( 
.A(n_876),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_725),
.B(n_654),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_729),
.B(n_654),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_832),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_799),
.B(n_682),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_807),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_757),
.A2(n_703),
.B1(n_697),
.B2(n_696),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_735),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_766),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_852),
.Y(n_961)
);

BUFx8_ASAP7_75t_L g962 ( 
.A(n_832),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_802),
.B(n_649),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_731),
.B(n_649),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_802),
.B(n_657),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_783),
.B(n_657),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_775),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_725),
.B(n_654),
.Y(n_968)
);

AND2x6_ASAP7_75t_SL g969 ( 
.A(n_828),
.B(n_410),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_SL g970 ( 
.A1(n_863),
.A2(n_368),
.B1(n_379),
.B2(n_378),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_748),
.B(n_663),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_785),
.B(n_663),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_832),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_757),
.Y(n_974)
);

NOR2x1p5_ASAP7_75t_L g975 ( 
.A(n_839),
.B(n_371),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_L g976 ( 
.A(n_806),
.B(n_666),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_828),
.B(n_619),
.Y(n_977)
);

INVx4_ASAP7_75t_L g978 ( 
.A(n_750),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_735),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_788),
.B(n_666),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_747),
.B(n_654),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_840),
.A2(n_703),
.B1(n_697),
.B2(n_693),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_858),
.A2(n_693),
.B1(n_674),
.B2(n_671),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_747),
.B(n_654),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_808),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_792),
.B(n_671),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_745),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_746),
.B(n_654),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_734),
.Y(n_989)
);

INVx5_ASAP7_75t_L g990 ( 
.A(n_750),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_858),
.A2(n_674),
.B1(n_619),
.B2(n_638),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_877),
.B(n_627),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_751),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_863),
.A2(n_638),
.B1(n_634),
.B2(n_632),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_877),
.B(n_627),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_860),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_827),
.B(n_410),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_750),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_865),
.Y(n_999)
);

INVx2_ASAP7_75t_SL g1000 ( 
.A(n_840),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_750),
.B(n_628),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_750),
.B(n_628),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_866),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_793),
.B(n_632),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_759),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_868),
.B(n_634),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_844),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_760),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_735),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_746),
.B(n_413),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_867),
.B(n_413),
.Y(n_1011)
);

NOR2x1p5_ASAP7_75t_L g1012 ( 
.A(n_841),
.B(n_334),
.Y(n_1012)
);

AND2x6_ASAP7_75t_SL g1013 ( 
.A(n_834),
.B(n_0),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_868),
.B(n_573),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_767),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_808),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_868),
.B(n_573),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_844),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_868),
.B(n_576),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_868),
.B(n_576),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_SL g1021 ( 
.A(n_825),
.B(n_338),
.C(n_391),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_774),
.A2(n_594),
.B(n_622),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_754),
.B(n_579),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_868),
.B(n_579),
.Y(n_1024)
);

INVx4_ASAP7_75t_L g1025 ( 
.A(n_808),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_724),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_780),
.B(n_584),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_834),
.A2(n_822),
.B1(n_826),
.B2(n_817),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_817),
.A2(n_692),
.B1(n_622),
.B2(n_621),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_756),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_823),
.A2(n_692),
.B1(n_621),
.B2(n_611),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_859),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_738),
.B(n_581),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_780),
.B(n_584),
.Y(n_1034)
);

NOR2xp67_ASAP7_75t_L g1035 ( 
.A(n_845),
.B(n_581),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_859),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_808),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_754),
.B(n_584),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_798),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_871),
.B(n_584),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_848),
.B(n_586),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_871),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_741),
.B(n_586),
.Y(n_1043)
);

OR2x6_ASAP7_75t_L g1044 ( 
.A(n_849),
.B(n_588),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_849),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_803),
.B(n_584),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_833),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_823),
.A2(n_692),
.B1(n_611),
.B2(n_609),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_732),
.Y(n_1049)
);

BUFx8_ASAP7_75t_L g1050 ( 
.A(n_733),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_741),
.B(n_588),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_855),
.Y(n_1052)
);

AND2x2_ASAP7_75t_L g1053 ( 
.A(n_875),
.B(n_594),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_749),
.B(n_596),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_875),
.A2(n_596),
.B1(n_608),
.B2(n_606),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_749),
.B(n_600),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_977),
.A2(n_770),
.B(n_850),
.C(n_846),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1007),
.B(n_825),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_900),
.B(n_945),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_887),
.A2(n_753),
.B(n_848),
.Y(n_1060)
);

INVx1_ASAP7_75t_SL g1061 ( 
.A(n_878),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_915),
.B(n_882),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_887),
.A2(n_912),
.B(n_899),
.Y(n_1063)
);

BUFx8_ASAP7_75t_L g1064 ( 
.A(n_895),
.Y(n_1064)
);

INVx5_ASAP7_75t_L g1065 ( 
.A(n_942),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_888),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_911),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1032),
.A2(n_835),
.B(n_853),
.C(n_872),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_900),
.B(n_777),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1042),
.B(n_870),
.Y(n_1070)
);

BUFx4f_ASAP7_75t_L g1071 ( 
.A(n_881),
.Y(n_1071)
);

O2A1O1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1036),
.A2(n_835),
.B(n_873),
.C(n_776),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_1039),
.A2(n_857),
.B1(n_816),
.B2(n_812),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_884),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1000),
.B(n_1018),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_899),
.A2(n_753),
.B(n_812),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_969),
.B(n_857),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_920),
.A2(n_929),
.B(n_957),
.C(n_1021),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_908),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_974),
.A2(n_772),
.B1(n_763),
.B2(n_769),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_912),
.A2(n_772),
.B(n_763),
.Y(n_1081)
);

OAI22x1_ASAP7_75t_L g1082 ( 
.A1(n_938),
.A2(n_795),
.B1(n_801),
.B2(n_776),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_990),
.B(n_787),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_946),
.A2(n_809),
.B(n_810),
.C(n_801),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_1016),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_951),
.A2(n_797),
.B(n_795),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_990),
.B(n_800),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_SL g1088 ( 
.A(n_921),
.B(n_338),
.C(n_390),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_960),
.B(n_769),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_927),
.B(n_600),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_989),
.B(n_906),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_951),
.A2(n_810),
.B(n_797),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_967),
.B(n_782),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1052),
.A2(n_782),
.B(n_606),
.C(n_609),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_952),
.B(n_602),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_SL g1096 ( 
.A1(n_978),
.A2(n_608),
.B(n_605),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_879),
.A2(n_605),
.B(n_603),
.C(n_602),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_924),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_934),
.B(n_603),
.Y(n_1099)
);

CKINVDCx6p67_ASAP7_75t_R g1100 ( 
.A(n_900),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_1011),
.B(n_805),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_896),
.A2(n_390),
.B(n_389),
.C(n_341),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_879),
.A2(n_1),
.B(n_2),
.C(n_9),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_997),
.B(n_341),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_L g1105 ( 
.A1(n_971),
.A2(n_361),
.B(n_351),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_897),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_956),
.A2(n_296),
.B(n_382),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_956),
.A2(n_965),
.B(n_963),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1028),
.A2(n_351),
.B(n_354),
.C(n_359),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_904),
.B(n_354),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_992),
.A2(n_389),
.B1(n_359),
.B2(n_366),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_905),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_926),
.Y(n_1113)
);

INVx6_ASAP7_75t_L g1114 ( 
.A(n_1050),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_963),
.A2(n_373),
.B(n_364),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_935),
.B(n_361),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_883),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_971),
.A2(n_361),
.B(n_139),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_990),
.B(n_1045),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_992),
.A2(n_333),
.B1(n_254),
.B2(n_252),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_900),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1016),
.Y(n_1122)
);

INVx4_ASAP7_75t_L g1123 ( 
.A(n_945),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_936),
.Y(n_1124)
);

INVx4_ASAP7_75t_L g1125 ( 
.A(n_945),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_913),
.B(n_2),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_1016),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_922),
.B(n_251),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_925),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1037),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_883),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_944),
.B(n_9),
.Y(n_1132)
);

BUFx12f_ASAP7_75t_L g1133 ( 
.A(n_962),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_1010),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_965),
.A2(n_256),
.B(n_330),
.Y(n_1135)
);

CKINVDCx16_ASAP7_75t_R g1136 ( 
.A(n_1010),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_990),
.B(n_257),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_995),
.A2(n_258),
.B(n_328),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_995),
.A2(n_260),
.B(n_327),
.Y(n_1139)
);

INVx4_ASAP7_75t_L g1140 ( 
.A(n_945),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1004),
.A2(n_267),
.B(n_324),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_976),
.A2(n_290),
.B(n_320),
.C(n_319),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_898),
.A2(n_286),
.B(n_315),
.C(n_313),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_935),
.B(n_10),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1037),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1053),
.A2(n_284),
.B(n_305),
.C(n_293),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1004),
.A2(n_272),
.B(n_288),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_892),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_987),
.B(n_275),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_978),
.B(n_13),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1045),
.B(n_283),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_931),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_1047),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_998),
.B(n_276),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_998),
.B(n_361),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_948),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_R g1157 ( 
.A(n_1025),
.B(n_14),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1006),
.A2(n_80),
.B(n_198),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1037),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_917),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_962),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1006),
.A2(n_70),
.B(n_197),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_933),
.B(n_15),
.C(n_16),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_975),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_993),
.B(n_15),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_937),
.A2(n_18),
.B(n_22),
.C(n_23),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_949),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_939),
.A2(n_87),
.B(n_195),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_1030),
.A2(n_361),
.B(n_25),
.C(n_30),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_939),
.A2(n_86),
.B(n_191),
.Y(n_1170)
);

NOR3xp33_ASAP7_75t_SL g1171 ( 
.A(n_943),
.B(n_24),
.C(n_25),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_970),
.B(n_953),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_950),
.B(n_31),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_916),
.A2(n_32),
.B(n_35),
.C(n_36),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1014),
.A2(n_96),
.B(n_187),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_961),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_910),
.B(n_36),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1014),
.A2(n_92),
.B(n_185),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_889),
.A2(n_361),
.B(n_43),
.C(n_46),
.Y(n_1179)
);

AOI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1040),
.A2(n_361),
.B(n_91),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_907),
.A2(n_39),
.B(n_43),
.C(n_46),
.Y(n_1181)
);

INVx4_ASAP7_75t_SL g1182 ( 
.A(n_919),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_916),
.B(n_39),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_918),
.A2(n_47),
.B(n_49),
.C(n_51),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_949),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_953),
.B(n_361),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_996),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1017),
.A2(n_128),
.B(n_158),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_893),
.B(n_51),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_918),
.B(n_52),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_928),
.B(n_54),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_999),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1017),
.A2(n_130),
.B(n_84),
.Y(n_1193)
);

O2A1O1Ixp5_ASAP7_75t_L g1194 ( 
.A1(n_909),
.A2(n_60),
.B(n_100),
.C(n_104),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_889),
.A2(n_60),
.B(n_131),
.C(n_147),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_880),
.B(n_155),
.Y(n_1196)
);

O2A1O1Ixp33_ASAP7_75t_L g1197 ( 
.A1(n_928),
.A2(n_162),
.B(n_930),
.C(n_1012),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1049),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_SL g1199 ( 
.A1(n_1046),
.A2(n_983),
.B(n_991),
.C(n_985),
.Y(n_1199)
);

AOI32xp33_ASAP7_75t_L g1200 ( 
.A1(n_1013),
.A2(n_886),
.A3(n_973),
.B1(n_955),
.B2(n_901),
.Y(n_1200)
);

INVx8_ASAP7_75t_L g1201 ( 
.A(n_1044),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_930),
.A2(n_972),
.B(n_980),
.C(n_1033),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1019),
.A2(n_1020),
.B(n_1024),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1022),
.A2(n_1056),
.B(n_1043),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_972),
.A2(n_980),
.B(n_1033),
.C(n_986),
.Y(n_1205)
);

OAI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_940),
.A2(n_902),
.B1(n_986),
.B2(n_966),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1063),
.A2(n_1024),
.B(n_1020),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1204),
.A2(n_1019),
.B(n_894),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_1114),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1118),
.A2(n_1056),
.B(n_1043),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1058),
.A2(n_966),
.B1(n_941),
.B2(n_923),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1062),
.B(n_1005),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1061),
.B(n_1008),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1199),
.A2(n_1051),
.B(n_1054),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1108),
.A2(n_1001),
.B(n_1002),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1061),
.B(n_1015),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1203),
.A2(n_1001),
.B(n_1002),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1114),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1180),
.A2(n_1054),
.B(n_1051),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1105),
.A2(n_964),
.B(n_1035),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1136),
.B(n_903),
.Y(n_1221)
);

OA21x2_ASAP7_75t_L g1222 ( 
.A1(n_1076),
.A2(n_1029),
.B(n_1031),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1144),
.A2(n_982),
.B1(n_958),
.B2(n_994),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1060),
.A2(n_1048),
.B(n_1055),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1081),
.A2(n_991),
.B(n_983),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1134),
.B(n_1026),
.Y(n_1226)
);

OAI22x1_ASAP7_75t_L g1227 ( 
.A1(n_1077),
.A2(n_1041),
.B1(n_1003),
.B2(n_985),
.Y(n_1227)
);

INVx5_ASAP7_75t_L g1228 ( 
.A(n_1201),
.Y(n_1228)
);

NOR4xp25_ASAP7_75t_L g1229 ( 
.A(n_1103),
.B(n_932),
.C(n_891),
.D(n_954),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1104),
.B(n_1153),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1071),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1057),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1153),
.B(n_885),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_1067),
.Y(n_1234)
);

OR2x2_ASAP7_75t_L g1235 ( 
.A(n_1075),
.B(n_1044),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_1179),
.B(n_1041),
.C(n_1044),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1068),
.A2(n_968),
.B(n_914),
.C(n_1023),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1097),
.A2(n_1034),
.B(n_1027),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1084),
.A2(n_1038),
.B(n_1025),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1086),
.A2(n_947),
.B(n_890),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1082),
.A2(n_1023),
.A3(n_1034),
.B(n_1027),
.Y(n_1241)
);

AO31x2_ASAP7_75t_L g1242 ( 
.A1(n_1206),
.A2(n_885),
.A3(n_979),
.B(n_959),
.Y(n_1242)
);

AOI211x1_ASAP7_75t_L g1243 ( 
.A1(n_1070),
.A2(n_981),
.B(n_984),
.C(n_1009),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1096),
.A2(n_959),
.B(n_979),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1206),
.B(n_1101),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1090),
.B(n_959),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1189),
.A2(n_968),
.B1(n_914),
.B2(n_988),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1092),
.A2(n_1009),
.B(n_979),
.Y(n_1248)
);

INVx4_ASAP7_75t_L g1249 ( 
.A(n_1071),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1158),
.A2(n_1009),
.B(n_988),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1116),
.A2(n_1195),
.A3(n_1143),
.B(n_1102),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1106),
.B(n_1112),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1116),
.A2(n_1194),
.B(n_1073),
.Y(n_1253)
);

O2A1O1Ixp33_ASAP7_75t_SL g1254 ( 
.A1(n_1183),
.A2(n_1190),
.B(n_1191),
.C(n_1177),
.Y(n_1254)
);

NOR2x1_ASAP7_75t_SL g1255 ( 
.A(n_1119),
.B(n_1121),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1094),
.A2(n_1162),
.B(n_1188),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1059),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1167),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1089),
.B(n_1093),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1064),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1073),
.A2(n_1072),
.B(n_1165),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1167),
.B(n_1185),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1185),
.B(n_1182),
.Y(n_1264)
);

NOR2xp67_ASAP7_75t_L g1265 ( 
.A(n_1091),
.B(n_1065),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1175),
.A2(n_1178),
.B(n_1193),
.Y(n_1266)
);

NOR4xp25_ASAP7_75t_L g1267 ( 
.A(n_1174),
.B(n_1184),
.C(n_1166),
.D(n_1169),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1168),
.A2(n_1170),
.B(n_1087),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1197),
.A2(n_1150),
.B(n_1155),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1150),
.A2(n_1132),
.B(n_1154),
.Y(n_1270)
);

OAI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1080),
.A2(n_1078),
.B(n_1109),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1099),
.B(n_1152),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1148),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1083),
.A2(n_1186),
.B(n_1080),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1172),
.A2(n_1111),
.B1(n_1149),
.B2(n_1148),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1137),
.A2(n_1095),
.B(n_1173),
.Y(n_1276)
);

INVx3_ASAP7_75t_SL g1277 ( 
.A(n_1065),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1115),
.A2(n_1135),
.B(n_1107),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1111),
.A2(n_1128),
.B1(n_1120),
.B2(n_1124),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1160),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1126),
.A2(n_1117),
.B(n_1131),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1138),
.A2(n_1139),
.B(n_1141),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1200),
.B(n_1187),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1147),
.A2(n_1069),
.B(n_1110),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_1151),
.B(n_1164),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1098),
.B(n_1176),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1117),
.A2(n_1131),
.B(n_1156),
.Y(n_1287)
);

OAI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1146),
.A2(n_1142),
.B(n_1120),
.Y(n_1288)
);

NAND2x1p5_ASAP7_75t_L g1289 ( 
.A(n_1059),
.B(n_1140),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1113),
.B(n_1192),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1157),
.A2(n_1181),
.B(n_1201),
.Y(n_1291)
);

AOI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1201),
.A2(n_1160),
.B1(n_1196),
.B2(n_1161),
.Y(n_1292)
);

OAI21xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1123),
.A2(n_1140),
.B(n_1125),
.Y(n_1293)
);

NAND2xp33_ASAP7_75t_R g1294 ( 
.A(n_1088),
.B(n_1079),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1198),
.Y(n_1295)
);

OAI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1163),
.A2(n_1171),
.B(n_1069),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1157),
.A2(n_1130),
.B(n_1145),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1085),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1085),
.B(n_1127),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1122),
.A2(n_1130),
.B(n_1145),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1122),
.A2(n_1127),
.B(n_1145),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1159),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1065),
.B(n_1100),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1133),
.B(n_1064),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1060),
.Y(n_1305)
);

INVx5_ASAP7_75t_L g1306 ( 
.A(n_1201),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1204),
.A2(n_1118),
.B(n_971),
.Y(n_1307)
);

NAND2x1p5_ASAP7_75t_L g1308 ( 
.A(n_1119),
.B(n_1167),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1203),
.A2(n_1108),
.B(n_1063),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1066),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1082),
.A2(n_1206),
.A3(n_1108),
.B(n_1203),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1136),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1204),
.A2(n_1118),
.B(n_971),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1204),
.A2(n_1118),
.B(n_971),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1066),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1066),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1150),
.B(n_1042),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1060),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1136),
.B(n_740),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1060),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1062),
.B(n_1042),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1063),
.B(n_957),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1203),
.A2(n_1108),
.B(n_1063),
.Y(n_1323)
);

AOI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1105),
.A2(n_1204),
.B(n_1108),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1060),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1136),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1059),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_R g1328 ( 
.A(n_1136),
.B(n_688),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1070),
.B(n_1042),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_1075),
.B(n_819),
.Y(n_1330)
);

CKINVDCx5p33_ASAP7_75t_R g1331 ( 
.A(n_1064),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1074),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1167),
.B(n_1185),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1063),
.A2(n_1076),
.B(n_1060),
.Y(n_1334)
);

INVxp67_ASAP7_75t_SL g1335 ( 
.A(n_1134),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1136),
.B(n_740),
.Y(n_1336)
);

AOI221xp5_ASAP7_75t_L g1337 ( 
.A1(n_1058),
.A2(n_616),
.B1(n_742),
.B2(n_710),
.C(n_882),
.Y(n_1337)
);

OA22x2_ASAP7_75t_L g1338 ( 
.A1(n_1172),
.A2(n_574),
.B1(n_500),
.B2(n_501),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1063),
.A2(n_1108),
.B(n_1203),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1063),
.B(n_957),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1064),
.Y(n_1341)
);

AOI211x1_ASAP7_75t_L g1342 ( 
.A1(n_1058),
.A2(n_790),
.B(n_929),
.C(n_920),
.Y(n_1342)
);

AO21x1_ASAP7_75t_L g1343 ( 
.A1(n_1063),
.A2(n_1206),
.B(n_1101),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1066),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1062),
.B(n_1042),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1063),
.A2(n_1108),
.B(n_1203),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1074),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_SL g1348 ( 
.A1(n_1197),
.A2(n_1063),
.B(n_1202),
.Y(n_1348)
);

AND2x6_ASAP7_75t_L g1349 ( 
.A(n_1150),
.B(n_1059),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1057),
.A2(n_1032),
.B(n_1007),
.C(n_1018),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1058),
.A2(n_1042),
.B1(n_727),
.B2(n_1032),
.Y(n_1351)
);

AND2x2_ASAP7_75t_SL g1352 ( 
.A(n_1150),
.B(n_882),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1066),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1167),
.B(n_1185),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_L g1355 ( 
.A(n_1057),
.B(n_1042),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1338),
.A2(n_1337),
.B1(n_1352),
.B2(n_1351),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1277),
.Y(n_1357)
);

AO21x2_ASAP7_75t_L g1358 ( 
.A1(n_1262),
.A2(n_1324),
.B(n_1348),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1272),
.B(n_1321),
.Y(n_1359)
);

BUFx8_ASAP7_75t_L g1360 ( 
.A(n_1312),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1261),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1326),
.Y(n_1362)
);

AO32x2_ASAP7_75t_L g1363 ( 
.A1(n_1211),
.A2(n_1351),
.A3(n_1223),
.B1(n_1343),
.B2(n_1242),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1242),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1339),
.A2(n_1346),
.B(n_1256),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1307),
.A2(n_1314),
.B(n_1313),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1214),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1208),
.A2(n_1268),
.B(n_1266),
.Y(n_1369)
);

OA21x2_ASAP7_75t_L g1370 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1279),
.A2(n_1275),
.B1(n_1329),
.B2(n_1245),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1338),
.A2(n_1345),
.B1(n_1355),
.B2(n_1317),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1325),
.A2(n_1334),
.B(n_1220),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1264),
.B(n_1228),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1245),
.B(n_1235),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1210),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1271),
.B(n_1342),
.C(n_1262),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1271),
.A2(n_1288),
.B1(n_1232),
.B2(n_1234),
.Y(n_1378)
);

AND2x4_ASAP7_75t_L g1379 ( 
.A(n_1264),
.B(n_1228),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1350),
.A2(n_1254),
.B(n_1288),
.C(n_1267),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1242),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1311),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1249),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1224),
.A2(n_1207),
.B(n_1225),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1311),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1349),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1311),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1211),
.A2(n_1270),
.B(n_1225),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1230),
.B(n_1319),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1325),
.A2(n_1334),
.B(n_1219),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1215),
.A2(n_1217),
.B(n_1248),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1281),
.A2(n_1224),
.B(n_1239),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1309),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1280),
.B(n_1283),
.Y(n_1394)
);

BUFx4f_ASAP7_75t_SL g1395 ( 
.A(n_1249),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1322),
.A2(n_1340),
.B(n_1323),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1309),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1238),
.A2(n_1287),
.B(n_1244),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1283),
.A2(n_1296),
.B1(n_1236),
.B2(n_1292),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1260),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1274),
.A2(n_1250),
.B(n_1278),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1223),
.A2(n_1227),
.A3(n_1237),
.B(n_1247),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1336),
.B(n_1246),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1236),
.A2(n_1269),
.B(n_1259),
.C(n_1296),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1267),
.A2(n_1282),
.B(n_1259),
.C(n_1229),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1276),
.A2(n_1284),
.B(n_1222),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1331),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1222),
.A2(n_1253),
.B(n_1291),
.Y(n_1408)
);

NAND2xp33_ASAP7_75t_L g1409 ( 
.A(n_1349),
.B(n_1282),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_SL g1410 ( 
.A1(n_1297),
.A2(n_1255),
.B(n_1301),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1335),
.B(n_1310),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1253),
.A2(n_1240),
.B(n_1300),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1229),
.A2(n_1240),
.B(n_1293),
.Y(n_1413)
);

AO31x2_ASAP7_75t_L g1414 ( 
.A1(n_1315),
.A2(n_1316),
.A3(n_1344),
.B(n_1353),
.Y(n_1414)
);

AOI222xp33_ASAP7_75t_L g1415 ( 
.A1(n_1221),
.A2(n_1212),
.B1(n_1226),
.B2(n_1213),
.C1(n_1216),
.C2(n_1273),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1265),
.A2(n_1231),
.B1(n_1243),
.B2(n_1285),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1258),
.A2(n_1303),
.B(n_1233),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1308),
.A2(n_1289),
.B(n_1299),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1341),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1286),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1330),
.A2(n_1298),
.B(n_1302),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_1308),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1241),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_SL g1424 ( 
.A1(n_1209),
.A2(n_1304),
.B(n_1218),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1228),
.B(n_1306),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1303),
.A2(n_1295),
.B(n_1354),
.C(n_1333),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1286),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1263),
.A2(n_1354),
.B(n_1333),
.C(n_1327),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1209),
.A2(n_1263),
.B1(n_1290),
.B2(n_1347),
.C(n_1332),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1290),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1257),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1294),
.A2(n_1251),
.B1(n_1306),
.B2(n_1349),
.C(n_1279),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1251),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1251),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1324),
.A2(n_1313),
.B(n_1307),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1230),
.B(n_1321),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1349),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1242),
.Y(n_1438)
);

BUFx8_ASAP7_75t_L g1439 ( 
.A(n_1312),
.Y(n_1439)
);

CKINVDCx16_ASAP7_75t_R g1440 ( 
.A(n_1328),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1231),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1338),
.A2(n_1337),
.B1(n_882),
.B2(n_1352),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1349),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1337),
.A2(n_616),
.B1(n_742),
.B2(n_710),
.C(n_831),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1230),
.B(n_1321),
.Y(n_1446)
);

BUFx8_ASAP7_75t_SL g1447 ( 
.A(n_1261),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1351),
.A2(n_1032),
.B(n_1007),
.Y(n_1448)
);

AO21x2_ASAP7_75t_L g1449 ( 
.A1(n_1262),
.A2(n_1324),
.B(n_1348),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_L g1450 ( 
.A(n_1351),
.B(n_710),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1324),
.A2(n_1313),
.B(n_1307),
.Y(n_1451)
);

INVx4_ASAP7_75t_L g1452 ( 
.A(n_1249),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1214),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1252),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_SL g1455 ( 
.A1(n_1338),
.A2(n_1352),
.B1(n_412),
.B2(n_433),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1324),
.A2(n_1313),
.B(n_1307),
.Y(n_1456)
);

BUFx8_ASAP7_75t_L g1457 ( 
.A(n_1312),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1214),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1349),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1279),
.A2(n_1042),
.B1(n_1007),
.B2(n_1032),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1252),
.Y(n_1461)
);

AOI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1220),
.A2(n_1324),
.B(n_1105),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1231),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1324),
.A2(n_1313),
.B(n_1307),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1324),
.A2(n_1339),
.B(n_1346),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1214),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1351),
.B(n_710),
.Y(n_1467)
);

NAND2x1_ASAP7_75t_L g1468 ( 
.A(n_1348),
.B(n_1349),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1339),
.A2(n_1346),
.B(n_1063),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1470)
);

BUFx2_ASAP7_75t_SL g1471 ( 
.A(n_1265),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1355),
.A2(n_1351),
.B(n_1032),
.C(n_1007),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1214),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1351),
.A2(n_1032),
.B(n_1007),
.Y(n_1475)
);

OR2x6_ASAP7_75t_L g1476 ( 
.A(n_1243),
.B(n_1201),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1249),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1349),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1324),
.A2(n_1339),
.B(n_1346),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1324),
.A2(n_1339),
.B(n_1346),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1324),
.A2(n_1339),
.B(n_1346),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1324),
.A2(n_1339),
.B(n_1346),
.Y(n_1482)
);

AOI21xp5_ASAP7_75t_L g1483 ( 
.A1(n_1339),
.A2(n_1346),
.B(n_1063),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1355),
.A2(n_1351),
.B(n_1032),
.C(n_1007),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1305),
.A2(n_1320),
.B(n_1318),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1338),
.A2(n_1352),
.B1(n_412),
.B2(n_433),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1324),
.A2(n_1313),
.B(n_1307),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_SL g1489 ( 
.A1(n_1448),
.A2(n_1475),
.B(n_1466),
.C(n_1458),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1409),
.A2(n_1483),
.B(n_1469),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1375),
.B(n_1378),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1472),
.A2(n_1485),
.B(n_1467),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1384),
.A2(n_1380),
.B(n_1404),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1403),
.B(n_1436),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1450),
.A2(n_1467),
.B(n_1445),
.C(n_1356),
.Y(n_1495)
);

O2A1O1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1371),
.A2(n_1450),
.B(n_1460),
.C(n_1399),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1408),
.A2(n_1369),
.B(n_1465),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1356),
.A2(n_1442),
.B(n_1377),
.C(n_1372),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1375),
.B(n_1394),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1447),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1442),
.A2(n_1405),
.B(n_1394),
.C(n_1487),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_L g1502 ( 
.A1(n_1455),
.A2(n_1432),
.B(n_1413),
.C(n_1426),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1414),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1478),
.A2(n_1425),
.B(n_1416),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1446),
.B(n_1389),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1359),
.B(n_1411),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1360),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_SL g1508 ( 
.A1(n_1440),
.A2(n_1407),
.B1(n_1419),
.B2(n_1361),
.Y(n_1508)
);

O2A1O1Ixp33_ASAP7_75t_L g1509 ( 
.A1(n_1424),
.A2(n_1362),
.B(n_1421),
.C(n_1468),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1454),
.B(n_1461),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1478),
.A2(n_1428),
.B(n_1379),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1408),
.A2(n_1482),
.B(n_1481),
.Y(n_1512)
);

AND2x6_ASAP7_75t_L g1513 ( 
.A(n_1386),
.B(n_1437),
.Y(n_1513)
);

AND2x4_ASAP7_75t_L g1514 ( 
.A(n_1374),
.B(n_1379),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_1383),
.B(n_1452),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1364),
.A2(n_1484),
.B1(n_1486),
.B2(n_1443),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1400),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1437),
.B(n_1444),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1357),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1431),
.A2(n_1358),
.B(n_1449),
.C(n_1463),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1465),
.A2(n_1479),
.B(n_1482),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1370),
.A2(n_1474),
.B1(n_1470),
.B2(n_1443),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1479),
.A2(n_1481),
.B(n_1480),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1420),
.B(n_1427),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1430),
.B(n_1370),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1480),
.A2(n_1401),
.B(n_1406),
.Y(n_1526)
);

A2O1A1Ixp33_ASAP7_75t_L g1527 ( 
.A1(n_1429),
.A2(n_1433),
.B(n_1459),
.C(n_1444),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1441),
.B(n_1463),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1443),
.A2(n_1470),
.B1(n_1474),
.B2(n_1484),
.Y(n_1529)
);

OAI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1486),
.A2(n_1441),
.B1(n_1459),
.B2(n_1395),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1415),
.B(n_1402),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1417),
.B(n_1476),
.Y(n_1532)
);

INVxp33_ASAP7_75t_SL g1533 ( 
.A(n_1361),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1477),
.A2(n_1476),
.B1(n_1471),
.B2(n_1422),
.Y(n_1534)
);

NOR2xp67_ASAP7_75t_L g1535 ( 
.A(n_1477),
.B(n_1438),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1358),
.A2(n_1449),
.B(n_1466),
.C(n_1453),
.Y(n_1536)
);

OA21x2_ASAP7_75t_L g1537 ( 
.A1(n_1401),
.A2(n_1406),
.B(n_1366),
.Y(n_1537)
);

OA21x2_ASAP7_75t_L g1538 ( 
.A1(n_1366),
.A2(n_1373),
.B(n_1367),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1360),
.Y(n_1539)
);

INVx1_ASAP7_75t_SL g1540 ( 
.A(n_1365),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1418),
.B(n_1363),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1447),
.Y(n_1542)
);

A2O1A1Ixp33_ASAP7_75t_L g1543 ( 
.A1(n_1434),
.A2(n_1392),
.B(n_1363),
.C(n_1382),
.Y(n_1543)
);

AOI31xp33_ASAP7_75t_L g1544 ( 
.A1(n_1365),
.A2(n_1438),
.A3(n_1381),
.B(n_1363),
.Y(n_1544)
);

AOI21xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1390),
.A2(n_1434),
.B(n_1385),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1360),
.B(n_1457),
.Y(n_1546)
);

O2A1O1Ixp33_ASAP7_75t_L g1547 ( 
.A1(n_1368),
.A2(n_1473),
.B(n_1410),
.C(n_1376),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1367),
.A2(n_1488),
.B(n_1451),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1363),
.B(n_1402),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1435),
.A2(n_1464),
.B(n_1456),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1439),
.Y(n_1551)
);

O2A1O1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1376),
.A2(n_1387),
.B(n_1393),
.C(n_1397),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1392),
.A2(n_1396),
.B(n_1423),
.C(n_1402),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_SL g1554 ( 
.A1(n_1390),
.A2(n_1393),
.B(n_1397),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1412),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1398),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1407),
.A2(n_1419),
.B1(n_1439),
.B2(n_1457),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_SL g1558 ( 
.A1(n_1439),
.A2(n_1457),
.B1(n_1391),
.B2(n_1398),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1391),
.B(n_1462),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1357),
.Y(n_1560)
);

OA21x2_ASAP7_75t_L g1561 ( 
.A1(n_1408),
.A2(n_1369),
.B(n_1465),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1378),
.A2(n_1485),
.B(n_1472),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1375),
.B(n_1245),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1409),
.A2(n_1483),
.B(n_1469),
.Y(n_1564)
);

OA21x2_ASAP7_75t_L g1565 ( 
.A1(n_1408),
.A2(n_1369),
.B(n_1465),
.Y(n_1565)
);

A2O1A1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1450),
.A2(n_1467),
.B(n_1445),
.C(n_1275),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1378),
.A2(n_1485),
.B(n_1472),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1414),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1408),
.A2(n_1369),
.B(n_1465),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1403),
.B(n_1436),
.Y(n_1570)
);

AND2x2_ASAP7_75t_SL g1571 ( 
.A(n_1356),
.B(n_1450),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1403),
.B(n_1436),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1447),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1478),
.B(n_1374),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_SL g1575 ( 
.A1(n_1378),
.A2(n_1485),
.B(n_1472),
.Y(n_1575)
);

O2A1O1Ixp5_ASAP7_75t_L g1576 ( 
.A1(n_1378),
.A2(n_1388),
.B(n_1371),
.C(n_1262),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1408),
.A2(n_1369),
.B(n_1465),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1450),
.A2(n_1467),
.B(n_1445),
.C(n_1275),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1403),
.B(n_1436),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1375),
.B(n_1245),
.Y(n_1580)
);

CKINVDCx20_ASAP7_75t_R g1581 ( 
.A(n_1447),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1414),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1409),
.A2(n_1483),
.B(n_1469),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1403),
.B(n_1436),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1371),
.A2(n_1355),
.B(n_1485),
.C(n_1472),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1375),
.B(n_1245),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1411),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_1478),
.B(n_1374),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1375),
.B(n_1245),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1490),
.A2(n_1583),
.B(n_1564),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1587),
.B(n_1525),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1525),
.B(n_1491),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1503),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1491),
.B(n_1517),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1506),
.Y(n_1595)
);

AO21x2_ASAP7_75t_L g1596 ( 
.A1(n_1493),
.A2(n_1553),
.B(n_1543),
.Y(n_1596)
);

OAI211xp5_ASAP7_75t_L g1597 ( 
.A1(n_1496),
.A2(n_1562),
.B(n_1575),
.C(n_1567),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1541),
.B(n_1549),
.Y(n_1598)
);

AO21x2_ASAP7_75t_L g1599 ( 
.A1(n_1554),
.A2(n_1531),
.B(n_1544),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1558),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_SL g1601 ( 
.A(n_1532),
.B(n_1534),
.Y(n_1601)
);

OAI222xp33_ASAP7_75t_L g1602 ( 
.A1(n_1531),
.A2(n_1585),
.B1(n_1571),
.B2(n_1563),
.C1(n_1586),
.C2(n_1580),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1499),
.B(n_1516),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_R g1604 ( 
.A(n_1500),
.B(n_1542),
.Y(n_1604)
);

OA21x2_ASAP7_75t_L g1605 ( 
.A1(n_1576),
.A2(n_1544),
.B(n_1582),
.Y(n_1605)
);

INVx2_ASAP7_75t_SL g1606 ( 
.A(n_1528),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1568),
.A2(n_1545),
.B(n_1489),
.Y(n_1607)
);

INVx4_ASAP7_75t_L g1608 ( 
.A(n_1513),
.Y(n_1608)
);

INVxp67_ASAP7_75t_SL g1609 ( 
.A(n_1520),
.Y(n_1609)
);

AO21x2_ASAP7_75t_L g1610 ( 
.A1(n_1516),
.A2(n_1522),
.B(n_1529),
.Y(n_1610)
);

AO21x1_ASAP7_75t_SL g1611 ( 
.A1(n_1555),
.A2(n_1589),
.B(n_1586),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1499),
.B(n_1522),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1529),
.B(n_1563),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1494),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1572),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1579),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1584),
.B(n_1505),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1510),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1540),
.B(n_1524),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1559),
.Y(n_1620)
);

OA21x2_ASAP7_75t_L g1621 ( 
.A1(n_1556),
.A2(n_1527),
.B(n_1524),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1530),
.Y(n_1622)
);

OAI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1492),
.A2(n_1578),
.B(n_1566),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1530),
.B(n_1514),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1552),
.Y(n_1625)
);

NAND3xp33_ASAP7_75t_L g1626 ( 
.A(n_1501),
.B(n_1495),
.C(n_1498),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1535),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1547),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1502),
.A2(n_1509),
.B(n_1515),
.Y(n_1629)
);

AO21x2_ASAP7_75t_L g1630 ( 
.A1(n_1536),
.A2(n_1534),
.B(n_1504),
.Y(n_1630)
);

AOI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1550),
.A2(n_1548),
.B(n_1497),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1550),
.Y(n_1632)
);

AOI21x1_ASAP7_75t_L g1633 ( 
.A1(n_1548),
.A2(n_1561),
.B(n_1497),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1532),
.B(n_1551),
.Y(n_1634)
);

OR2x2_ASAP7_75t_L g1635 ( 
.A(n_1532),
.B(n_1507),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_L g1636 ( 
.A(n_1533),
.B(n_1508),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1513),
.B(n_1518),
.Y(n_1637)
);

BUFx6f_ASAP7_75t_L g1638 ( 
.A(n_1513),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1538),
.B(n_1512),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1513),
.B(n_1588),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1565),
.A2(n_1577),
.B(n_1569),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1569),
.B(n_1526),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1593),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1592),
.B(n_1537),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1613),
.B(n_1537),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1598),
.B(n_1611),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1603),
.B(n_1523),
.Y(n_1647)
);

AOI22xp33_ASAP7_75t_L g1648 ( 
.A1(n_1626),
.A2(n_1560),
.B1(n_1519),
.B2(n_1574),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1608),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1632),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1521),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1521),
.Y(n_1652)
);

BUFx2_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

OR2x6_ASAP7_75t_L g1654 ( 
.A(n_1638),
.B(n_1511),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1610),
.B(n_1620),
.Y(n_1655)
);

INVx3_ASAP7_75t_L g1656 ( 
.A(n_1633),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1610),
.B(n_1519),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1638),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1603),
.B(n_1612),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1610),
.B(n_1560),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1594),
.B(n_1557),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1642),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1642),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_SL g1664 ( 
.A(n_1623),
.B(n_1557),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1591),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1590),
.A2(n_1597),
.B(n_1596),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1590),
.B(n_1539),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1591),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1619),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1614),
.A2(n_1546),
.B1(n_1573),
.B2(n_1581),
.Y(n_1671)
);

AO21x2_ASAP7_75t_L g1672 ( 
.A1(n_1666),
.A2(n_1609),
.B(n_1631),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1646),
.B(n_1657),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1650),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1657),
.A2(n_1599),
.B1(n_1596),
.B2(n_1622),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1664),
.A2(n_1602),
.B(n_1600),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1671),
.Y(n_1677)
);

OA21x2_ASAP7_75t_L g1678 ( 
.A1(n_1666),
.A2(n_1633),
.B(n_1641),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1665),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1646),
.B(n_1606),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1657),
.B(n_1622),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_SL g1682 ( 
.A1(n_1660),
.A2(n_1600),
.B1(n_1608),
.B2(n_1638),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1664),
.A2(n_1629),
.B1(n_1635),
.B2(n_1634),
.Y(n_1683)
);

AOI211x1_ASAP7_75t_L g1684 ( 
.A1(n_1671),
.A2(n_1660),
.B(n_1659),
.C(n_1655),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1659),
.B(n_1618),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1660),
.B(n_1605),
.C(n_1628),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1665),
.B(n_1595),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1658),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1653),
.B(n_1624),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1643),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1655),
.A2(n_1599),
.B1(n_1596),
.B2(n_1625),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1669),
.B(n_1615),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1669),
.B(n_1616),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1667),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1653),
.B(n_1601),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1643),
.Y(n_1697)
);

INVxp67_ASAP7_75t_SL g1698 ( 
.A(n_1645),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1601),
.Y(n_1699)
);

BUFx12f_ASAP7_75t_L g1700 ( 
.A(n_1649),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1658),
.A2(n_1638),
.B1(n_1605),
.B2(n_1640),
.Y(n_1701)
);

INVx4_ASAP7_75t_L g1702 ( 
.A(n_1649),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1670),
.B(n_1617),
.Y(n_1703)
);

OAI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1654),
.A2(n_1605),
.B1(n_1637),
.B2(n_1621),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1679),
.Y(n_1705)
);

OA21x2_ASAP7_75t_L g1706 ( 
.A1(n_1686),
.A2(n_1675),
.B(n_1691),
.Y(n_1706)
);

NAND3xp33_ASAP7_75t_L g1707 ( 
.A(n_1676),
.B(n_1651),
.C(n_1668),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1692),
.B(n_1662),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1692),
.B(n_1662),
.Y(n_1709)
);

AND2x6_ASAP7_75t_L g1710 ( 
.A(n_1699),
.B(n_1640),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1686),
.A2(n_1656),
.B(n_1645),
.Y(n_1711)
);

AND4x1_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1648),
.C(n_1636),
.D(n_1668),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1678),
.Y(n_1713)
);

INVxp67_ASAP7_75t_L g1714 ( 
.A(n_1672),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1678),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1699),
.B(n_1696),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1678),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1661),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1690),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1674),
.A2(n_1652),
.B(n_1639),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1690),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1673),
.B(n_1663),
.Y(n_1723)
);

OAI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1683),
.A2(n_1668),
.B(n_1628),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1697),
.Y(n_1725)
);

BUFx6f_ASAP7_75t_L g1726 ( 
.A(n_1672),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1697),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1718),
.B(n_1684),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1719),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1716),
.B(n_1689),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1707),
.B(n_1694),
.Y(n_1731)
);

NOR2x1_ASAP7_75t_L g1732 ( 
.A(n_1707),
.B(n_1688),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_R g1733 ( 
.A(n_1718),
.B(n_1700),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1707),
.B(n_1696),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1684),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1705),
.B(n_1698),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1724),
.B(n_1681),
.Y(n_1737)
);

INVx5_ASAP7_75t_L g1738 ( 
.A(n_1726),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1724),
.B(n_1694),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1724),
.B(n_1644),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1716),
.B(n_1696),
.Y(n_1741)
);

NAND2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1712),
.B(n_1702),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1719),
.B(n_1644),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1712),
.B(n_1681),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1723),
.B(n_1680),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1712),
.A2(n_1701),
.B(n_1704),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1719),
.B(n_1687),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_SL g1748 ( 
.A(n_1710),
.B(n_1604),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1723),
.B(n_1680),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1706),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1706),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1727),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1706),
.A2(n_1672),
.B1(n_1630),
.B2(n_1607),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1708),
.B(n_1685),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1727),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1722),
.B(n_1725),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1708),
.B(n_1693),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.B(n_1688),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1706),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1727),
.B(n_1703),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1722),
.B(n_1647),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1720),
.B(n_1688),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1756),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1756),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1729),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1752),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1755),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1736),
.Y(n_1768)
);

NAND2x1p5_ASAP7_75t_L g1769 ( 
.A(n_1732),
.B(n_1682),
.Y(n_1769)
);

OAI221xp5_ASAP7_75t_L g1770 ( 
.A1(n_1746),
.A2(n_1706),
.B1(n_1714),
.B2(n_1726),
.C(n_1720),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1738),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1747),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1759),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1760),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1750),
.B(n_1722),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1738),
.Y(n_1776)
);

OAI21xp33_ASAP7_75t_L g1777 ( 
.A1(n_1728),
.A2(n_1711),
.B(n_1714),
.Y(n_1777)
);

NOR2xp67_ASAP7_75t_L g1778 ( 
.A(n_1734),
.B(n_1695),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1742),
.B(n_1720),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1751),
.B(n_1731),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1761),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1726),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1743),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1740),
.B(n_1709),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1743),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1740),
.B(n_1709),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1754),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1735),
.B(n_1709),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1744),
.A2(n_1706),
.B(n_1711),
.Y(n_1789)
);

INVx2_ASAP7_75t_SL g1790 ( 
.A(n_1741),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1757),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1731),
.Y(n_1792)
);

OAI322xp33_ASAP7_75t_L g1793 ( 
.A1(n_1739),
.A2(n_1737),
.A3(n_1726),
.B1(n_1715),
.B2(n_1721),
.C1(n_1713),
.C2(n_1717),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1733),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1738),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1745),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1745),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1749),
.B(n_1706),
.Y(n_1798)
);

INVx3_ASAP7_75t_L g1799 ( 
.A(n_1769),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1769),
.B(n_1734),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1769),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1773),
.B(n_1726),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1780),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1778),
.B(n_1738),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1794),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1773),
.B(n_1774),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1780),
.Y(n_1807)
);

OAI21x1_ASAP7_75t_L g1808 ( 
.A1(n_1789),
.A2(n_1753),
.B(n_1711),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1774),
.B(n_1763),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1779),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1779),
.B(n_1734),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1792),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1766),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1764),
.B(n_1726),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1790),
.B(n_1730),
.Y(n_1816)
);

AND3x1_ASAP7_75t_L g1817 ( 
.A(n_1777),
.B(n_1748),
.C(n_1758),
.Y(n_1817)
);

BUFx3_ASAP7_75t_L g1818 ( 
.A(n_1775),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1767),
.Y(n_1819)
);

BUFx2_ASAP7_75t_SL g1820 ( 
.A(n_1790),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1770),
.A2(n_1726),
.B1(n_1672),
.B2(n_1721),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1775),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1768),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1796),
.B(n_1730),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1771),
.Y(n_1825)
);

NOR2xp33_ASAP7_75t_L g1826 ( 
.A(n_1805),
.B(n_1772),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1805),
.B(n_1787),
.Y(n_1827)
);

NAND2x1_ASAP7_75t_L g1828 ( 
.A(n_1800),
.B(n_1799),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1818),
.Y(n_1829)
);

OAI222xp33_ASAP7_75t_L g1830 ( 
.A1(n_1807),
.A2(n_1798),
.B1(n_1788),
.B2(n_1758),
.C1(n_1762),
.C2(n_1738),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1800),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1818),
.Y(n_1832)
);

OAI211xp5_ASAP7_75t_SL g1833 ( 
.A1(n_1823),
.A2(n_1795),
.B(n_1776),
.C(n_1771),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1823),
.B(n_1791),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1818),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1818),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1817),
.A2(n_1793),
.B(n_1782),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1807),
.B(n_1783),
.Y(n_1838)
);

OAI31xp33_ASAP7_75t_SL g1839 ( 
.A1(n_1800),
.A2(n_1782),
.A3(n_1711),
.B(n_1762),
.Y(n_1839)
);

INVxp67_ASAP7_75t_L g1840 ( 
.A(n_1820),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1813),
.B(n_1797),
.Y(n_1841)
);

AOI322xp5_ASAP7_75t_L g1842 ( 
.A1(n_1803),
.A2(n_1784),
.A3(n_1786),
.B1(n_1715),
.B2(n_1713),
.C1(n_1717),
.C2(n_1721),
.Y(n_1842)
);

OAI21xp5_ASAP7_75t_L g1843 ( 
.A1(n_1808),
.A2(n_1785),
.B(n_1715),
.Y(n_1843)
);

NAND2x1p5_ASAP7_75t_L g1844 ( 
.A(n_1799),
.B(n_1682),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1816),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1822),
.B(n_1781),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1803),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1843),
.A2(n_1803),
.B1(n_1808),
.B2(n_1801),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1831),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1845),
.B(n_1816),
.Y(n_1850)
);

NAND2xp33_ASAP7_75t_L g1851 ( 
.A(n_1838),
.B(n_1733),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1826),
.B(n_1813),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1827),
.B(n_1822),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1829),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1832),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1835),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1834),
.B(n_1803),
.Y(n_1857)
);

NOR2x1_ASAP7_75t_R g1858 ( 
.A(n_1836),
.B(n_1820),
.Y(n_1858)
);

O2A1O1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1857),
.A2(n_1833),
.B(n_1847),
.C(n_1799),
.Y(n_1859)
);

NOR3xp33_ASAP7_75t_L g1860 ( 
.A(n_1853),
.B(n_1840),
.C(n_1799),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1850),
.B(n_1816),
.Y(n_1861)
);

AOI221xp5_ASAP7_75t_L g1862 ( 
.A1(n_1848),
.A2(n_1837),
.B1(n_1817),
.B2(n_1843),
.C(n_1821),
.Y(n_1862)
);

OAI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1848),
.A2(n_1839),
.B1(n_1821),
.B2(n_1799),
.C(n_1801),
.Y(n_1863)
);

NOR3xp33_ASAP7_75t_L g1864 ( 
.A(n_1852),
.B(n_1828),
.C(n_1846),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1849),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_R g1866 ( 
.A(n_1851),
.B(n_1841),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1849),
.B(n_1824),
.Y(n_1867)
);

AOI322xp5_ASAP7_75t_L g1868 ( 
.A1(n_1854),
.A2(n_1801),
.A3(n_1812),
.B1(n_1810),
.B2(n_1806),
.C1(n_1839),
.C2(n_1809),
.Y(n_1868)
);

XOR2xp5_ASAP7_75t_L g1869 ( 
.A(n_1867),
.B(n_1855),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1861),
.Y(n_1870)
);

AOI22xp5_ASAP7_75t_L g1871 ( 
.A1(n_1862),
.A2(n_1801),
.B1(n_1808),
.B2(n_1810),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1865),
.Y(n_1872)
);

AOI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1863),
.A2(n_1810),
.B1(n_1812),
.B2(n_1726),
.Y(n_1873)
);

OAI21xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1868),
.A2(n_1842),
.B(n_1812),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1874),
.B(n_1866),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1869),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1870),
.B(n_1864),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1872),
.Y(n_1878)
);

NOR2x1_ASAP7_75t_L g1879 ( 
.A(n_1873),
.B(n_1856),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1871),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1869),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1876),
.Y(n_1882)
);

NAND4xp75_ASAP7_75t_L g1883 ( 
.A(n_1875),
.B(n_1880),
.C(n_1881),
.D(n_1877),
.Y(n_1883)
);

INVx3_ASAP7_75t_SL g1884 ( 
.A(n_1878),
.Y(n_1884)
);

OAI22xp5_ASAP7_75t_SL g1885 ( 
.A1(n_1879),
.A2(n_1806),
.B1(n_1809),
.B2(n_1825),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1876),
.Y(n_1886)
);

CKINVDCx20_ASAP7_75t_R g1887 ( 
.A(n_1876),
.Y(n_1887)
);

XNOR2xp5_ASAP7_75t_L g1888 ( 
.A(n_1883),
.B(n_1860),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1884),
.B(n_1858),
.Y(n_1889)
);

INVx3_ASAP7_75t_SL g1890 ( 
.A(n_1887),
.Y(n_1890)
);

NOR4xp25_ASAP7_75t_SL g1891 ( 
.A(n_1885),
.B(n_1859),
.C(n_1814),
.D(n_1811),
.Y(n_1891)
);

OAI31xp33_ASAP7_75t_L g1892 ( 
.A1(n_1888),
.A2(n_1886),
.A3(n_1882),
.B(n_1830),
.Y(n_1892)
);

AOI32xp33_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1889),
.A3(n_1890),
.B1(n_1891),
.B2(n_1810),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1893),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1893),
.Y(n_1895)
);

OAI22x1_ASAP7_75t_L g1896 ( 
.A1(n_1895),
.A2(n_1844),
.B1(n_1825),
.B2(n_1819),
.Y(n_1896)
);

XNOR2x1_ASAP7_75t_L g1897 ( 
.A(n_1894),
.B(n_1844),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1810),
.B1(n_1819),
.B2(n_1811),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1896),
.A2(n_1802),
.B(n_1814),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1898),
.Y(n_1900)
);

XOR2xp5_ASAP7_75t_L g1901 ( 
.A(n_1900),
.B(n_1899),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1901),
.B(n_1776),
.Y(n_1902)
);

OAI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1802),
.B1(n_1815),
.B2(n_1795),
.Y(n_1903)
);

AOI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1804),
.B1(n_1815),
.B2(n_1824),
.Y(n_1904)
);

AOI211xp5_ASAP7_75t_L g1905 ( 
.A1(n_1904),
.A2(n_1804),
.B(n_1824),
.C(n_1726),
.Y(n_1905)
);


endmodule