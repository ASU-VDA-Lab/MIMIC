module fake_jpeg_8683_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_4),
.B(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

AND2x2_ASAP7_75t_SL g12 ( 
.A(n_5),
.B(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_22),
.Y(n_27)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.Y(n_25)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

FAx1_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_12),
.CI(n_17),
.CON(n_29),
.SN(n_29)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_14),
.B1(n_11),
.B2(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_1),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_14),
.B1(n_17),
.B2(n_11),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_30),
.B1(n_31),
.B2(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_21),
.B1(n_9),
.B2(n_16),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_18),
.A2(n_9),
.B1(n_15),
.B2(n_2),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_29),
.B(n_25),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_4),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_29),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_40),
.B1(n_37),
.B2(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_50),
.C(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_43),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_45),
.B(n_46),
.C(n_51),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_32),
.B(n_44),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_32),
.Y(n_58)
);


endmodule