module fake_jpeg_27977_n_273 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_273);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_9),
.B(n_3),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_38),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_3),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_29),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_33),
.B2(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_45),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_29),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_47),
.B1(n_56),
.B2(n_58),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_53),
.B(n_45),
.C(n_49),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_83),
.B(n_21),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_67),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_37),
.C(n_34),
.Y(n_68)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_38),
.C(n_24),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_41),
.A2(n_27),
.B1(n_31),
.B2(n_19),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_77),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_43),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_80),
.Y(n_95)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_75),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_59),
.A2(n_34),
.B1(n_31),
.B2(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_76),
.A2(n_78),
.B1(n_44),
.B2(n_47),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_34),
.B1(n_18),
.B2(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_32),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_20),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_20),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_44),
.A2(n_19),
.B1(n_30),
.B2(n_28),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_101),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_15),
.C(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_87),
.B(n_93),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_44),
.B1(n_56),
.B2(n_54),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_92),
.B1(n_97),
.B2(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_101),
.B1(n_108),
.B2(n_83),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_17),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_91),
.B(n_3),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_58),
.B1(n_51),
.B2(n_38),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_99),
.B(n_84),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_38),
.B1(n_22),
.B2(n_28),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_80),
.C(n_74),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_24),
.B(n_26),
.C(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_21),
.B1(n_32),
.B2(n_20),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_20),
.B1(n_26),
.B2(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_105),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_20),
.B1(n_26),
.B2(n_24),
.Y(n_108)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_116),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_67),
.B1(n_63),
.B2(n_79),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_131),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_64),
.B1(n_78),
.B2(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_123),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g150 ( 
.A1(n_118),
.A2(n_119),
.B(n_137),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_95),
.B(n_109),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_100),
.B(n_105),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_136),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_129),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_103),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_86),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_133),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_91),
.B(n_15),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_75),
.Y(n_136)
);

OAI21xp33_ASAP7_75t_SL g137 ( 
.A1(n_99),
.A2(n_4),
.B(n_5),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_153),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_114),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_127),
.B1(n_71),
.B2(n_126),
.Y(n_171)
);

NOR2x1_ASAP7_75t_R g152 ( 
.A(n_119),
.B(n_97),
.Y(n_152)
);

XOR2x2_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_157),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_159),
.Y(n_174)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_75),
.B(n_107),
.C(n_71),
.D(n_82),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_122),
.C(n_134),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_82),
.B(n_5),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_118),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_162),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_113),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_71),
.B1(n_85),
.B2(n_72),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_111),
.B(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_85),
.Y(n_165)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_181),
.C(n_182),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_130),
.B1(n_127),
.B2(n_135),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_169),
.A2(n_183),
.B1(n_160),
.B2(n_143),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_171),
.B(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_173),
.B(n_175),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_155),
.B1(n_163),
.B2(n_140),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_72),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_72),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_149),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_188),
.C(n_164),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_8),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_180),
.A2(n_142),
.B1(n_159),
.B2(n_153),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_191),
.A2(n_195),
.B1(n_200),
.B2(n_204),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_193),
.A2(n_203),
.B(n_210),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_197),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_152),
.B1(n_146),
.B2(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_201),
.B(n_208),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_157),
.C(n_150),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_146),
.B1(n_141),
.B2(n_151),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_202),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

HAxp5_ASAP7_75t_SL g211 ( 
.A(n_184),
.B(n_141),
.CON(n_211),
.SN(n_211)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_183),
.B1(n_168),
.B2(n_188),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_216),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_187),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_167),
.C(n_181),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_182),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_184),
.C(n_169),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_191),
.C(n_204),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_227),
.C(n_201),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_10),
.B(n_11),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_151),
.B1(n_154),
.B2(n_12),
.Y(n_225)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_226),
.B(n_199),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_154),
.Y(n_227)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_231),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_215),
.A2(n_196),
.B(n_222),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_235),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_198),
.B1(n_200),
.B2(n_210),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_238),
.B1(n_227),
.B2(n_217),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_198),
.B(n_197),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_216),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_228),
.C(n_236),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_213),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_249),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_239),
.B(n_224),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_246),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_218),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_247),
.A2(n_240),
.B1(n_243),
.B2(n_235),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_10),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g251 ( 
.A(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_251),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_254),
.C(n_241),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_234),
.B(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_255),
.Y(n_260)
);

OAI21xp33_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_238),
.B(n_11),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_256),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_10),
.C(n_11),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_252),
.C(n_12),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_12),
.B(n_13),
.C(n_251),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_260),
.Y(n_269)
);

NAND2xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_262),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_268),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_264),
.Y(n_273)
);


endmodule