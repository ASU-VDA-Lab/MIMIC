module fake_netlist_5_194_n_1885 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1885);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1885;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_368;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g189 ( 
.A(n_61),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_107),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_158),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_63),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_37),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_51),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_60),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_29),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_75),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_154),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_134),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_0),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_71),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_56),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_8),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_155),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_3),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_0),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_76),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_42),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_43),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_58),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_141),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_4),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_135),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_36),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_167),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_81),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_166),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_92),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_39),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_78),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_103),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_80),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_24),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_146),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_157),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_28),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_28),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_46),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_77),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_25),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_85),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_65),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_149),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_102),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_176),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_45),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_51),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_138),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_116),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_21),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_114),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_21),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_79),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_41),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_131),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_37),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_97),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_12),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_175),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_34),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_12),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_87),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_66),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_31),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_82),
.Y(n_276)
);

BUFx8_ASAP7_75t_SL g277 ( 
.A(n_162),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_115),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_35),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_29),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_132),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_111),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_109),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_86),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_17),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_46),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_20),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_23),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_129),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_130),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_127),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_16),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_1),
.Y(n_293)
);

INVxp33_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_124),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_160),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_161),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_70),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_137),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_106),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_178),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_39),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_2),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_147),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_153),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_22),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_93),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_91),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_74),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_32),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_52),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_27),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_38),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_9),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_119),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_35),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_22),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_26),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_45),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_83),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_24),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_73),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_159),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_14),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_11),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_89),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_42),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_16),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_4),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_180),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_55),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_95),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_19),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_185),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_183),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_59),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_40),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_14),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_33),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_19),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_52),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_99),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_174),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_105),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_118),
.Y(n_345)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_148),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_44),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_184),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g349 ( 
.A(n_2),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_49),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_113),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_139),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_64),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_88),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_84),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_121),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_164),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_177),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_90),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_152),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_20),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_123),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_96),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_27),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_43),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_94),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_67),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_30),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_125),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_69),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_17),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_101),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_3),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_18),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_49),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_133),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_349),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_349),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_224),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_349),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_277),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_205),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_363),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_271),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_359),
.B(n_5),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_191),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_192),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_193),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_196),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_224),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_242),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_349),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_264),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_228),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_230),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_223),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_303),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_223),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_195),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g404 ( 
.A(n_223),
.B(n_5),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_303),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_231),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_232),
.Y(n_407)
);

BUFx6f_ASAP7_75t_SL g408 ( 
.A(n_366),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_303),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_246),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_359),
.B(n_6),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_280),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_303),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_242),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_238),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_244),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_253),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_254),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_316),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_276),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_311),
.B(n_6),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_233),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_316),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_316),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_316),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_276),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_278),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_211),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_350),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_251),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_278),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_350),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_248),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_298),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_248),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_321),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_255),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_298),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_233),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_259),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_261),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_285),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_285),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_287),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_301),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_345),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_265),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_267),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_367),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_287),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_293),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_293),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_301),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_345),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_256),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_338),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_269),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_331),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_338),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_274),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_194),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_364),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_367),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g467 ( 
.A(n_369),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_281),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_331),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_237),
.B(n_7),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_203),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_379),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_393),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_401),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_404),
.B(n_369),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_388),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_389),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_400),
.B(n_237),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_409),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_206),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_409),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_394),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_414),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_392),
.B(n_397),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_399),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_406),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_413),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_407),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_415),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_416),
.B(n_417),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_418),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_R g496 ( 
.A(n_382),
.B(n_439),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_402),
.B(n_419),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_396),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_419),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_441),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_423),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_441),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_448),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_442),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_443),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_430),
.B(n_309),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_423),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g509 ( 
.A(n_387),
.B(n_346),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_449),
.B(n_272),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_451),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_425),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_450),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_272),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_429),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_459),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_377),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_462),
.B(n_330),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_422),
.B(n_311),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_431),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_468),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_386),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_433),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_420),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_471),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_426),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_427),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_434),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_432),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_378),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_436),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_378),
.B(n_330),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_440),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_381),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_381),
.B(n_189),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_447),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_383),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_428),
.B(n_366),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_455),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_460),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_383),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_390),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_476),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_536),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_509),
.B(n_481),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_477),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_SL g555 ( 
.A1(n_510),
.A2(n_385),
.B1(n_384),
.B2(n_411),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_501),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_481),
.B(n_273),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_536),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_509),
.B(n_428),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_542),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_509),
.A2(n_351),
.B1(n_467),
.B2(n_456),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_501),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_520),
.B(n_408),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_498),
.B(n_503),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_512),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_542),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_550),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_481),
.B(n_273),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_546),
.B(n_351),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_504),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_499),
.B(n_410),
.Y(n_575)
);

AND3x2_ASAP7_75t_L g576 ( 
.A(n_530),
.B(n_470),
.C(n_457),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_511),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_390),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_545),
.Y(n_580)
);

INVx2_ASAP7_75t_SL g581 ( 
.A(n_504),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_539),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_514),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_498),
.B(n_408),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_498),
.B(n_408),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_483),
.B(n_463),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_487),
.A2(n_494),
.B1(n_507),
.B2(n_478),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_514),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_481),
.B(n_395),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_545),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_550),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_521),
.B(n_412),
.C(n_403),
.Y(n_592)
);

INVx5_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_545),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_539),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_549),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_540),
.A2(n_421),
.B1(n_197),
.B2(n_266),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_521),
.B(n_380),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_543),
.B(n_273),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_475),
.B(n_435),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_549),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_512),
.Y(n_602)
);

OR2x2_ASAP7_75t_L g603 ( 
.A(n_475),
.B(n_380),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_549),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_475),
.B(n_438),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_543),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_475),
.B(n_435),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_512),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_488),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_480),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_543),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_543),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_488),
.B(n_519),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_540),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_512),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_540),
.A2(n_347),
.B1(n_240),
.B2(n_236),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_529),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_488),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_488),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_519),
.B(n_395),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_535),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_535),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_540),
.B(n_273),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_531),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_474),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_519),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_489),
.B(n_438),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_519),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_474),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_516),
.B(n_291),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_472),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_SL g632 ( 
.A(n_490),
.B(n_279),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_538),
.B(n_398),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_516),
.A2(n_341),
.B1(n_260),
.B2(n_241),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_532),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_492),
.B(n_291),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_474),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_473),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_516),
.B(n_291),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_493),
.B(n_291),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_495),
.B(n_190),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_505),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_474),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_538),
.B(n_474),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_538),
.B(n_398),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_506),
.B(n_198),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_479),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_508),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_508),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_538),
.B(n_464),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_508),
.B(n_218),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_508),
.Y(n_652)
);

AND2x6_ASAP7_75t_L g653 ( 
.A(n_516),
.B(n_199),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_508),
.B(n_243),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_515),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_479),
.B(n_464),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_482),
.Y(n_657)
);

OR2x6_ASAP7_75t_L g658 ( 
.A(n_485),
.B(n_465),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_482),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_518),
.B(n_200),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_491),
.B(n_249),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_491),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_497),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_497),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_486),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_537),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_500),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_500),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_526),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_502),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_502),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_513),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_513),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_204),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_517),
.B(n_215),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_522),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_522),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_541),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_523),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_523),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_524),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_527),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_544),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_496),
.B(n_465),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_525),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_525),
.B(n_295),
.Y(n_686)
);

INVx3_ASAP7_75t_L g687 ( 
.A(n_528),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_528),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_533),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_533),
.B(n_367),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_547),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_548),
.B(n_437),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_534),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_536),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_472),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_481),
.B(n_221),
.Y(n_696)
);

BUFx10_ASAP7_75t_L g697 ( 
.A(n_527),
.Y(n_697)
);

AO22x2_ASAP7_75t_L g698 ( 
.A1(n_546),
.A2(n_339),
.B1(n_317),
.B2(n_312),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_545),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_498),
.B(n_296),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_510),
.B(n_201),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_476),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_614),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_553),
.A2(n_263),
.B1(n_225),
.B2(n_376),
.Y(n_704)
);

INVx6_ASAP7_75t_L g705 ( 
.A(n_689),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_682),
.B(n_279),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_586),
.B(n_201),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_614),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_579),
.B(n_589),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_606),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_586),
.B(n_202),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_650),
.B(n_466),
.Y(n_712)
);

OAI221xp5_ASAP7_75t_L g713 ( 
.A1(n_616),
.A2(n_220),
.B1(n_319),
.B2(n_219),
.C(n_262),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_650),
.B(n_466),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_551),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_553),
.A2(n_283),
.B1(n_372),
.B2(n_360),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_606),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_568),
.B(n_367),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_568),
.B(n_367),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_701),
.B(n_469),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_567),
.B(n_367),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_611),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_701),
.B(n_294),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_603),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_564),
.A2(n_258),
.B1(n_307),
.B2(n_252),
.Y(n_725)
);

AO22x1_ASAP7_75t_L g726 ( 
.A1(n_605),
.A2(n_340),
.B1(n_337),
.B2(n_333),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_611),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_560),
.B(n_202),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_552),
.B(n_227),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_561),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_560),
.B(n_207),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_684),
.B(n_207),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_559),
.B(n_229),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_612),
.Y(n_734)
);

O2A1O1Ixp5_ASAP7_75t_L g735 ( 
.A1(n_571),
.A2(n_284),
.B(n_358),
.C(n_355),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_598),
.B(n_210),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_610),
.B(n_208),
.Y(n_737)
);

INVx8_ASAP7_75t_L g738 ( 
.A(n_658),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_563),
.B(n_235),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_575),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_692),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_598),
.B(n_210),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_627),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_641),
.B(n_212),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_569),
.B(n_239),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_SL g746 ( 
.A(n_682),
.B(n_292),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_605),
.B(n_256),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_641),
.B(n_212),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_570),
.B(n_367),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_612),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_554),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_565),
.Y(n_752)
);

O2A1O1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_555),
.A2(n_286),
.B(n_375),
.C(n_374),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_608),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_592),
.B(n_203),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_600),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_591),
.B(n_289),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_696),
.A2(n_334),
.B1(n_336),
.B2(n_342),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_694),
.B(n_662),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_697),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_558),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_587),
.B(n_216),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_658),
.B(n_213),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_646),
.B(n_216),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_696),
.A2(n_290),
.B1(n_353),
.B2(n_371),
.Y(n_765)
);

AOI221xp5_ASAP7_75t_L g766 ( 
.A1(n_698),
.A2(n_310),
.B1(n_325),
.B2(n_292),
.C(n_288),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_646),
.B(n_217),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_617),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_558),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_566),
.B(n_217),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_662),
.B(n_668),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_668),
.B(n_297),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_658),
.B(n_631),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_572),
.B(n_250),
.C(n_373),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_638),
.B(n_213),
.Y(n_775)
);

BUFx5_ASAP7_75t_L g776 ( 
.A(n_628),
.Y(n_776)
);

O2A1O1Ixp5_ASAP7_75t_L g777 ( 
.A1(n_571),
.A2(n_461),
.B(n_458),
.C(n_454),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_562),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_633),
.B(n_299),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_645),
.B(n_300),
.Y(n_780)
);

BUFx5_ASAP7_75t_L g781 ( 
.A(n_628),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_562),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_620),
.B(n_304),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_596),
.B(n_305),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_642),
.B(n_256),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_601),
.B(n_308),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_669),
.B(n_461),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_604),
.B(n_315),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_696),
.B(n_653),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_660),
.B(n_222),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_574),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_L g792 ( 
.A(n_696),
.B(n_320),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_609),
.B(n_322),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_618),
.B(n_323),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_619),
.B(n_626),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_660),
.B(n_222),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_600),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_693),
.B(n_209),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_671),
.B(n_326),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_636),
.B(n_282),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_671),
.B(n_356),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_584),
.A2(n_357),
.B1(n_370),
.B2(n_362),
.Y(n_802)
);

OAI22xp5_ASAP7_75t_L g803 ( 
.A1(n_700),
.A2(n_282),
.B1(n_332),
.B2(n_335),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_680),
.B(n_332),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_680),
.B(n_335),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_644),
.A2(n_343),
.B(n_344),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_584),
.A2(n_365),
.B(n_313),
.C(n_302),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_566),
.B(n_343),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_696),
.A2(n_268),
.B1(n_368),
.B2(n_328),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_600),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_655),
.B(n_344),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_607),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_617),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_585),
.A2(n_361),
.B(n_354),
.C(n_352),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_607),
.Y(n_815)
);

NAND2xp33_ASAP7_75t_L g816 ( 
.A(n_653),
.B(n_348),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_608),
.A2(n_607),
.B1(n_602),
.B2(n_615),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_636),
.B(n_348),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_687),
.B(n_352),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_676),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_574),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_565),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_585),
.A2(n_354),
.B1(n_325),
.B2(n_310),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_676),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_687),
.B(n_226),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_677),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_640),
.B(n_573),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_677),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_632),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_556),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_689),
.B(n_234),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_681),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_640),
.B(n_366),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_572),
.A2(n_327),
.B1(n_245),
.B2(n_247),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_683),
.B(n_62),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_681),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_581),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_672),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_647),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_602),
.B(n_257),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_577),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_577),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_615),
.B(n_314),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_608),
.A2(n_270),
.B1(n_275),
.B2(n_306),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_630),
.B(n_329),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_578),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_630),
.A2(n_214),
.B1(n_288),
.B2(n_333),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_582),
.B(n_318),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_578),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_613),
.B(n_324),
.Y(n_850)
);

OAI221xp5_ASAP7_75t_L g851 ( 
.A1(n_616),
.A2(n_634),
.B1(n_597),
.B2(n_656),
.C(n_661),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_657),
.B(n_663),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_664),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_667),
.B(n_458),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_653),
.A2(n_214),
.B1(n_337),
.B2(n_340),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_670),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_595),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_624),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_576),
.Y(n_859)
);

OAI21xp33_ASAP7_75t_L g860 ( 
.A1(n_597),
.A2(n_698),
.B(n_634),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_686),
.B(n_454),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_679),
.B(n_453),
.Y(n_862)
);

NAND3xp33_ASAP7_75t_L g863 ( 
.A(n_656),
.B(n_453),
.C(n_452),
.Y(n_863)
);

AND2x6_ASAP7_75t_SL g864 ( 
.A(n_665),
.B(n_452),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_688),
.B(n_446),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_L g866 ( 
.A(n_691),
.B(n_98),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_688),
.B(n_446),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_693),
.B(n_445),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_688),
.B(n_445),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_688),
.B(n_444),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_583),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_740),
.B(n_624),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_838),
.B(n_651),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_709),
.A2(n_594),
.B(n_580),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_709),
.A2(n_594),
.B(n_580),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_832),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_817),
.A2(n_698),
.B1(n_691),
.B2(n_654),
.Y(n_877)
);

AO32x1_ASAP7_75t_L g878 ( 
.A1(n_704),
.A2(n_702),
.A3(n_583),
.B1(n_588),
.B2(n_621),
.Y(n_878)
);

AND2x6_ASAP7_75t_L g879 ( 
.A(n_827),
.B(n_625),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_787),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_850),
.B(n_685),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_865),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_789),
.A2(n_594),
.B(n_649),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_860),
.A2(n_623),
.B(n_690),
.C(n_588),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_723),
.A2(n_653),
.B1(n_674),
.B2(n_675),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_728),
.A2(n_731),
.B1(n_748),
.B2(n_744),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_712),
.A2(n_623),
.B(n_690),
.Y(n_887)
);

OR2x2_ASAP7_75t_L g888 ( 
.A(n_775),
.B(n_695),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_718),
.A2(n_625),
.B(n_629),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_715),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_832),
.B(n_697),
.Y(n_891)
);

BUFx12f_ASAP7_75t_L g892 ( 
.A(n_859),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_771),
.A2(n_590),
.B(n_561),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_712),
.A2(n_590),
.B(n_561),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_714),
.A2(n_590),
.B(n_561),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_754),
.B(n_590),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_720),
.B(n_635),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_741),
.B(n_635),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_706),
.B(n_666),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_764),
.B(n_678),
.C(n_437),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_865),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_850),
.B(n_557),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_867),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_832),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_743),
.B(n_678),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_852),
.B(n_557),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_852),
.B(n_557),
.Y(n_907)
);

A2O1A1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_767),
.A2(n_702),
.B(n_621),
.C(n_622),
.Y(n_908)
);

A2O1A1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_790),
.A2(n_622),
.B(n_629),
.C(n_648),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_714),
.A2(n_648),
.B(n_652),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_839),
.B(n_557),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_853),
.B(n_557),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_721),
.A2(n_652),
.B(n_653),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_856),
.B(n_675),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_796),
.A2(n_675),
.B1(n_674),
.B2(n_599),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_800),
.A2(n_444),
.B(n_659),
.C(n_673),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_721),
.A2(n_699),
.B(n_593),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_851),
.A2(n_674),
.B(n_675),
.C(n_659),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_718),
.A2(n_719),
.B(n_754),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_773),
.Y(n_920)
);

OAI21x1_ASAP7_75t_L g921 ( 
.A1(n_795),
.A2(n_599),
.B(n_675),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_705),
.A2(n_659),
.B1(n_673),
.B2(n_643),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_719),
.A2(n_593),
.B(n_699),
.Y(n_923)
);

OAI21x1_ASAP7_75t_L g924 ( 
.A1(n_795),
.A2(n_599),
.B(n_674),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_759),
.B(n_825),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_730),
.A2(n_593),
.B(n_699),
.Y(n_926)
);

AO21x1_ASAP7_75t_L g927 ( 
.A1(n_716),
.A2(n_674),
.B(n_599),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_783),
.A2(n_699),
.B(n_593),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_847),
.A2(n_697),
.B(n_643),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_836),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_707),
.B(n_643),
.Y(n_931)
);

AOI21xp33_ASAP7_75t_L g932 ( 
.A1(n_725),
.A2(n_7),
.B(n_8),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_825),
.B(n_659),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_836),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_762),
.A2(n_673),
.B(n_599),
.C(n_639),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_867),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_711),
.B(n_829),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_783),
.A2(n_780),
.B(n_779),
.Y(n_938)
);

AOI21x1_ASAP7_75t_L g939 ( 
.A1(n_779),
.A2(n_643),
.B(n_637),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_768),
.B(n_673),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_760),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_780),
.A2(n_799),
.B(n_772),
.Y(n_942)
);

NAND2xp33_ASAP7_75t_L g943 ( 
.A(n_776),
.B(n_639),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_801),
.A2(n_637),
.B(n_639),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_724),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_747),
.B(n_637),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_836),
.B(n_637),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_840),
.A2(n_639),
.B(n_68),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_843),
.A2(n_639),
.B(n_188),
.Y(n_949)
);

OAI321xp33_ASAP7_75t_L g950 ( 
.A1(n_766),
.A2(n_10),
.A3(n_11),
.B1(n_13),
.B2(n_15),
.C(n_18),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_820),
.B(n_10),
.Y(n_951)
);

OR2x2_ASAP7_75t_L g952 ( 
.A(n_868),
.B(n_13),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_756),
.A2(n_104),
.B1(n_179),
.B2(n_172),
.Y(n_953)
);

INVx1_ASAP7_75t_SL g954 ( 
.A(n_813),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_793),
.A2(n_181),
.B(n_169),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_793),
.A2(n_168),
.B(n_163),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_785),
.B(n_830),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_823),
.A2(n_15),
.B1(n_26),
.B2(n_30),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_746),
.B(n_156),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_705),
.A2(n_144),
.B1(n_143),
.B2(n_140),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_794),
.A2(n_136),
.B(n_128),
.Y(n_961)
);

OAI22xp5_ASAP7_75t_L g962 ( 
.A1(n_705),
.A2(n_122),
.B1(n_117),
.B2(n_110),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_868),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_794),
.A2(n_108),
.B(n_32),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_710),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_868),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_824),
.B(n_38),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_736),
.B(n_40),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_753),
.A2(n_54),
.B(n_44),
.C(n_47),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_792),
.A2(n_41),
.B(n_47),
.Y(n_970)
);

CKINVDCx10_ASAP7_75t_R g971 ( 
.A(n_737),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_784),
.A2(n_48),
.B(n_50),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_858),
.B(n_48),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_784),
.A2(n_50),
.B(n_53),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_777),
.A2(n_53),
.B(n_54),
.Y(n_975)
);

NOR2x1_ASAP7_75t_L g976 ( 
.A(n_835),
.B(n_811),
.Y(n_976)
);

BUFx12f_ASAP7_75t_L g977 ( 
.A(n_859),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_786),
.A2(n_788),
.B(n_815),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_703),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_752),
.B(n_822),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_786),
.A2(n_788),
.B(n_812),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_763),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_814),
.A2(n_749),
.B(n_845),
.Y(n_983)
);

NAND3xp33_ASAP7_75t_L g984 ( 
.A(n_717),
.B(n_734),
.C(n_750),
.Y(n_984)
);

AOI22x1_ASAP7_75t_L g985 ( 
.A1(n_722),
.A2(n_727),
.B1(n_708),
.B2(n_826),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_R g986 ( 
.A(n_837),
.B(n_857),
.Y(n_986)
);

AOI22x1_ASAP7_75t_L g987 ( 
.A1(n_828),
.A2(n_871),
.B1(n_821),
.B2(n_751),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_797),
.A2(n_810),
.B(n_819),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_761),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_769),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_778),
.A2(n_782),
.B(n_791),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_831),
.B(n_805),
.Y(n_992)
);

CKINVDCx6p67_ASAP7_75t_R g993 ( 
.A(n_738),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_798),
.Y(n_994)
);

BUFx6f_ASAP7_75t_L g995 ( 
.A(n_798),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_869),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_869),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_804),
.A2(n_844),
.B(n_757),
.C(n_729),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_861),
.A2(n_749),
.B(n_739),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_841),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_798),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_870),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_870),
.A2(n_846),
.B(n_842),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_733),
.B(n_745),
.Y(n_1004)
);

AOI21x1_ASAP7_75t_L g1005 ( 
.A1(n_849),
.A2(n_862),
.B(n_854),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_737),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_802),
.B(n_774),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_SL g1008 ( 
.A(n_834),
.B(n_855),
.C(n_755),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_803),
.B(n_732),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_742),
.B(n_808),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_776),
.B(n_781),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_770),
.A2(n_818),
.B1(n_833),
.B2(n_816),
.Y(n_1012)
);

AND2x6_ASAP7_75t_SL g1013 ( 
.A(n_737),
.B(n_862),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_776),
.B(n_781),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_L g1015 ( 
.A(n_726),
.B(n_848),
.C(n_713),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_765),
.A2(n_809),
.B1(n_758),
.B2(n_866),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_807),
.B(n_854),
.C(n_806),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_738),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_735),
.A2(n_863),
.B(n_776),
.C(n_781),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_776),
.B(n_781),
.Y(n_1020)
);

AO32x2_ASAP7_75t_L g1021 ( 
.A1(n_776),
.A2(n_716),
.A3(n_704),
.B1(n_587),
.B2(n_803),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_738),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_781),
.B(n_864),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_781),
.A2(n_860),
.B1(n_509),
.B2(n_851),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_740),
.B(n_379),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_832),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_704),
.B(n_553),
.C(n_850),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_715),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_858),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_741),
.B(n_598),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_741),
.B(n_598),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_762),
.A2(n_553),
.B(n_814),
.C(n_709),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_817),
.A2(n_709),
.B1(n_827),
.B2(n_771),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_838),
.B(n_709),
.Y(n_1039)
);

AND2x6_ASAP7_75t_L g1040 ( 
.A(n_709),
.B(n_827),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_865),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_787),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_865),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_744),
.A2(n_764),
.B(n_767),
.C(n_748),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_754),
.B(n_832),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_740),
.B(n_379),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_715),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_838),
.B(n_709),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_860),
.A2(n_553),
.B(n_851),
.C(n_762),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_838),
.B(n_709),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_860),
.A2(n_553),
.B(n_851),
.C(n_762),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_838),
.B(n_709),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_709),
.A2(n_714),
.B(n_712),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1056)
);

A2O1A1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_744),
.A2(n_764),
.B(n_767),
.C(n_748),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_744),
.A2(n_764),
.B(n_767),
.C(n_748),
.Y(n_1058)
);

NOR2x1_ASAP7_75t_L g1059 ( 
.A(n_835),
.B(n_682),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_709),
.A2(n_568),
.B(n_608),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_817),
.A2(n_709),
.B1(n_827),
.B2(n_771),
.Y(n_1061)
);

AOI221xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1044),
.A2(n_1058),
.B1(n_1057),
.B2(n_958),
.C(n_968),
.Y(n_1062)
);

NAND2xp33_ASAP7_75t_SL g1063 ( 
.A(n_1022),
.B(n_1023),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_886),
.B(n_1039),
.Y(n_1064)
);

AOI21x1_ASAP7_75t_SL g1065 ( 
.A1(n_902),
.A2(n_914),
.B(n_992),
.Y(n_1065)
);

AOI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_897),
.A2(n_1010),
.B(n_1049),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_904),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_892),
.Y(n_1069)
);

AND3x4_ASAP7_75t_L g1070 ( 
.A(n_872),
.B(n_900),
.C(n_1031),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_977),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_941),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_1035),
.A2(n_1052),
.B(n_1036),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1048),
.B(n_1050),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1053),
.A2(n_1060),
.B(n_1056),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_938),
.A2(n_983),
.B(n_1055),
.C(n_1061),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_993),
.Y(n_1077)
);

INVx6_ASAP7_75t_L g1078 ( 
.A(n_904),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1054),
.B(n_881),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_921),
.A2(n_919),
.B(n_939),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1055),
.A2(n_1038),
.B(n_946),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_890),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_896),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_894),
.A2(n_895),
.B(n_987),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_925),
.A2(n_887),
.B(n_978),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1008),
.A2(n_958),
.B(n_982),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_893),
.A2(n_1003),
.B(n_883),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_910),
.A2(n_1005),
.B(n_917),
.Y(n_1088)
);

AND2x4_ASAP7_75t_L g1089 ( 
.A(n_963),
.B(n_1022),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1032),
.B(n_1034),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_887),
.A2(n_981),
.B(n_913),
.Y(n_1091)
);

AOI21x1_ASAP7_75t_L g1092 ( 
.A1(n_942),
.A2(n_933),
.B(n_1011),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_913),
.A2(n_875),
.B(n_874),
.Y(n_1093)
);

BUFx12f_ASAP7_75t_L g1094 ( 
.A(n_1022),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_910),
.A2(n_988),
.B(n_923),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_954),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1040),
.B(n_882),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_985),
.A2(n_944),
.B(n_928),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_927),
.A2(n_877),
.A3(n_909),
.B(n_908),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_896),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_SL g1101 ( 
.A1(n_906),
.A2(n_907),
.B(n_911),
.Y(n_1101)
);

NOR2x1_ASAP7_75t_L g1102 ( 
.A(n_1059),
.B(n_898),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1014),
.A2(n_1020),
.B(n_999),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1029),
.A2(n_1051),
.B(n_983),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_969),
.A2(n_998),
.A3(n_1016),
.B(n_916),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1004),
.A2(n_1037),
.B(n_918),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1040),
.B(n_901),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_884),
.A2(n_873),
.B(n_943),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1029),
.A2(n_1002),
.B(n_936),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1040),
.B(n_903),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_945),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1040),
.B(n_996),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1019),
.A2(n_926),
.B(n_935),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_997),
.A2(n_1041),
.B(n_1043),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_947),
.A2(n_948),
.B(n_949),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1024),
.A2(n_931),
.B(n_878),
.Y(n_1116)
);

AO31x2_ASAP7_75t_L g1117 ( 
.A1(n_970),
.A2(n_972),
.A3(n_974),
.B(n_878),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_922),
.A2(n_912),
.B(n_990),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_1017),
.A2(n_984),
.B(n_975),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_888),
.B(n_982),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_1009),
.A2(n_1017),
.B(n_1007),
.C(n_964),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_SL g1122 ( 
.A1(n_975),
.A2(n_961),
.B(n_955),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_880),
.B(n_1042),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_878),
.A2(n_915),
.B(n_984),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_937),
.B(n_957),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_976),
.A2(n_1012),
.B(n_934),
.Y(n_1126)
);

AOI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1025),
.A2(n_1046),
.B(n_905),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_1015),
.A2(n_929),
.B(n_885),
.C(n_932),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_956),
.A2(n_1030),
.B(n_1000),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1045),
.A2(n_1047),
.B(n_989),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_876),
.B(n_930),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_979),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_951),
.A2(n_967),
.B(n_962),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_879),
.B(n_980),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_904),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1026),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_891),
.A2(n_959),
.B(n_960),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_879),
.B(n_980),
.Y(n_1138)
);

BUFx12f_ASAP7_75t_L g1139 ( 
.A(n_994),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_L g1140 ( 
.A1(n_965),
.A2(n_1021),
.B(n_879),
.C(n_952),
.Y(n_1140)
);

AO21x1_ASAP7_75t_L g1141 ( 
.A1(n_953),
.A2(n_1021),
.B(n_950),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_940),
.A2(n_1018),
.B(n_1006),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_920),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_1021),
.A2(n_879),
.B(n_973),
.C(n_950),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_966),
.A2(n_1026),
.B(n_1001),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_954),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_899),
.B(n_994),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1026),
.A2(n_986),
.B(n_1013),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_995),
.B(n_994),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_995),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_SL g1151 ( 
.A1(n_995),
.A2(n_1057),
.B(n_1044),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_971),
.B(n_886),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_886),
.B(n_1039),
.Y(n_1154)
);

OAI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_886),
.A2(n_723),
.B(n_632),
.Y(n_1155)
);

INVx4_ASAP7_75t_L g1156 ( 
.A(n_904),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1032),
.B(n_1034),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_1031),
.Y(n_1159)
);

AOI211x1_ASAP7_75t_L g1160 ( 
.A1(n_958),
.A2(n_860),
.B(n_932),
.C(n_1039),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_886),
.A2(n_1044),
.B(n_1058),
.C(n_1057),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_890),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_886),
.B(n_1039),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_1031),
.B(n_738),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_963),
.B(n_1022),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_886),
.A2(n_1057),
.B1(n_1058),
.B2(n_1044),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_889),
.A2(n_991),
.B(n_924),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_890),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_886),
.B(n_1039),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_889),
.A2(n_991),
.B(n_924),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_904),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_886),
.B(n_1039),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_990),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_SL g1182 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_889),
.A2(n_991),
.B(n_924),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1184)
);

HB1xp67_ASAP7_75t_L g1185 ( 
.A(n_945),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_886),
.A2(n_1044),
.B(n_1058),
.C(n_1057),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_904),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_SL g1189 ( 
.A1(n_902),
.A2(n_914),
.B(n_992),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_889),
.A2(n_991),
.B(n_924),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_889),
.A2(n_991),
.B(n_924),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1031),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_890),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1194)
);

AOI21x1_ASAP7_75t_SL g1195 ( 
.A1(n_902),
.A2(n_914),
.B(n_992),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_904),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_886),
.B(n_1039),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1027),
.A2(n_1033),
.B(n_1028),
.Y(n_1198)
);

INVx4_ASAP7_75t_L g1199 ( 
.A(n_904),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_886),
.B(n_1044),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_990),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_889),
.A2(n_991),
.B(n_924),
.Y(n_1202)
);

OAI211xp5_ASAP7_75t_L g1203 ( 
.A1(n_886),
.A2(n_766),
.B(n_823),
.C(n_564),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_SL g1204 ( 
.A(n_897),
.B(n_768),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_904),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_897),
.B(n_886),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_890),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_990),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1032),
.B(n_1034),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_SL g1210 ( 
.A1(n_1049),
.A2(n_1051),
.B(n_927),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_886),
.A2(n_1057),
.B1(n_1058),
.B2(n_1044),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1044),
.A2(n_1058),
.B(n_1057),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_886),
.B(n_1039),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1089),
.B(n_1167),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1079),
.B(n_1074),
.Y(n_1215)
);

AND2x2_ASAP7_75t_SL g1216 ( 
.A(n_1206),
.B(n_1204),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1146),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1159),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1082),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1089),
.B(n_1167),
.Y(n_1220)
);

CKINVDCx6p67_ASAP7_75t_R g1221 ( 
.A(n_1094),
.Y(n_1221)
);

INVxp67_ASAP7_75t_SL g1222 ( 
.A(n_1185),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1177),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1163),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_1177),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1173),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1155),
.A2(n_1200),
.B1(n_1066),
.B2(n_1169),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1192),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1182),
.A2(n_1184),
.B(n_1085),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1158),
.B(n_1209),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1090),
.B(n_1125),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_1111),
.B(n_1120),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_L g1233 ( 
.A(n_1064),
.B(n_1154),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1203),
.A2(n_1086),
.B1(n_1211),
.B2(n_1170),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1085),
.A2(n_1091),
.B(n_1093),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1177),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1193),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_1196),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1207),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1150),
.B(n_1149),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1090),
.B(n_1147),
.Y(n_1241)
);

AO32x1_ASAP7_75t_L g1242 ( 
.A1(n_1141),
.A2(n_1062),
.A3(n_1212),
.B1(n_1161),
.B2(n_1179),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1096),
.B(n_1127),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1091),
.A2(n_1093),
.B(n_1106),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1083),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1185),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1106),
.A2(n_1108),
.B(n_1153),
.Y(n_1247)
);

OR2x6_ASAP7_75t_L g1248 ( 
.A(n_1166),
.B(n_1139),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_SL g1249 ( 
.A1(n_1203),
.A2(n_1152),
.B1(n_1180),
.B2(n_1188),
.Y(n_1249)
);

OR2x6_ASAP7_75t_L g1250 ( 
.A(n_1166),
.B(n_1151),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1181),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1143),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1162),
.A2(n_1186),
.B(n_1128),
.C(n_1197),
.Y(n_1253)
);

OAI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1165),
.A2(n_1213),
.B1(n_1174),
.B2(n_1178),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1123),
.B(n_1132),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1114),
.B(n_1160),
.Y(n_1256)
);

AO21x2_ASAP7_75t_L g1257 ( 
.A1(n_1104),
.A2(n_1122),
.B(n_1116),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1196),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1109),
.B(n_1081),
.Y(n_1259)
);

BUFx2_ASAP7_75t_L g1260 ( 
.A(n_1150),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1071),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1134),
.B(n_1138),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1148),
.B(n_1201),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1076),
.B(n_1121),
.C(n_1137),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1166),
.Y(n_1265)
);

AOI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1070),
.A2(n_1063),
.B1(n_1107),
.B2(n_1097),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1208),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1108),
.A2(n_1175),
.B(n_1153),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1135),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1068),
.A2(n_1175),
.B(n_1157),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1130),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1077),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1110),
.A2(n_1112),
.B1(n_1210),
.B2(n_1137),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1131),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1136),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1102),
.B(n_1145),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1205),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1072),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1076),
.A2(n_1164),
.B(n_1157),
.Y(n_1279)
);

OR2x6_ASAP7_75t_L g1280 ( 
.A(n_1145),
.B(n_1067),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1068),
.A2(n_1164),
.B(n_1168),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1205),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1121),
.A2(n_1144),
.B(n_1126),
.C(n_1140),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1205),
.Y(n_1284)
);

HB1xp67_ASAP7_75t_L g1285 ( 
.A(n_1078),
.Y(n_1285)
);

O2A1O1Ixp5_ASAP7_75t_SL g1286 ( 
.A1(n_1100),
.A2(n_1065),
.B(n_1195),
.C(n_1189),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1069),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_SL g1288 ( 
.A(n_1067),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1078),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1081),
.B(n_1126),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1078),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1156),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1073),
.A2(n_1171),
.B(n_1075),
.Y(n_1293)
);

BUFx2_ASAP7_75t_SL g1294 ( 
.A(n_1156),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1142),
.Y(n_1296)
);

CKINVDCx8_ASAP7_75t_R g1297 ( 
.A(n_1119),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1199),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1199),
.B(n_1100),
.Y(n_1299)
);

OR2x2_ASAP7_75t_L g1300 ( 
.A(n_1105),
.B(n_1133),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1116),
.A2(n_1124),
.B(n_1144),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_SL g1302 ( 
.A1(n_1124),
.A2(n_1129),
.B(n_1073),
.C(n_1075),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1129),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1168),
.A2(n_1198),
.B(n_1194),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1105),
.B(n_1099),
.Y(n_1305)
);

AOI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1095),
.A2(n_1088),
.B1(n_1113),
.B2(n_1118),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1115),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1103),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_L g1309 ( 
.A(n_1171),
.B(n_1194),
.C(n_1198),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1105),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1117),
.B(n_1099),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1098),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1099),
.Y(n_1313)
);

INVx1_ASAP7_75t_SL g1314 ( 
.A(n_1172),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1099),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1117),
.B(n_1092),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1087),
.A2(n_1084),
.B(n_1080),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1065),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1176),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1183),
.A2(n_1190),
.B(n_1191),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1117),
.A2(n_1189),
.B1(n_1195),
.B2(n_1101),
.Y(n_1321)
);

AND2x6_ASAP7_75t_L g1322 ( 
.A(n_1101),
.B(n_1117),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1202),
.A2(n_1085),
.B(n_938),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1158),
.B(n_1209),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1079),
.B(n_1074),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1089),
.B(n_1167),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1085),
.A2(n_938),
.B(n_1079),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1062),
.A2(n_886),
.B(n_1211),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1079),
.B(n_1074),
.Y(n_1329)
);

INVx3_ASAP7_75t_L g1330 ( 
.A(n_1083),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1089),
.B(n_1167),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1192),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1159),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1082),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1120),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1182),
.A2(n_1184),
.B(n_1085),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1146),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1085),
.A2(n_938),
.B(n_1079),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1206),
.A2(n_886),
.B1(n_1203),
.B2(n_1155),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1079),
.B(n_1074),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1177),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1206),
.A2(n_886),
.B(n_1057),
.C(n_1044),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1079),
.B(n_1074),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1159),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_1159),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1159),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1082),
.Y(n_1347)
);

BUFx2_ASAP7_75t_SL g1348 ( 
.A(n_1159),
.Y(n_1348)
);

INVx8_ASAP7_75t_L g1349 ( 
.A(n_1094),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1082),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1120),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1206),
.A2(n_1155),
.B1(n_886),
.B2(n_1200),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1089),
.B(n_1167),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1182),
.A2(n_1184),
.B(n_1085),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1089),
.B(n_1167),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1206),
.A2(n_886),
.B1(n_1203),
.B2(n_1155),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1158),
.B(n_1209),
.Y(n_1357)
);

NOR2xp67_ASAP7_75t_L g1358 ( 
.A(n_1125),
.B(n_682),
.Y(n_1358)
);

NAND2x1_ASAP7_75t_L g1359 ( 
.A(n_1083),
.B(n_1100),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1071),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1083),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1249),
.A2(n_1352),
.B1(n_1356),
.B2(n_1339),
.Y(n_1362)
);

INVx3_ASAP7_75t_L g1363 ( 
.A(n_1250),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1339),
.A2(n_1356),
.B1(n_1216),
.B2(n_1234),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1250),
.Y(n_1365)
);

INVxp33_ASAP7_75t_L g1366 ( 
.A(n_1243),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1215),
.B(n_1325),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1219),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1333),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1224),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_SL g1371 ( 
.A1(n_1231),
.A2(n_1254),
.B1(n_1241),
.B2(n_1233),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1239),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1226),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1215),
.B(n_1325),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1342),
.A2(n_1227),
.B(n_1254),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1234),
.B(n_1329),
.Y(n_1376)
);

AND2x4_ASAP7_75t_L g1377 ( 
.A(n_1250),
.B(n_1240),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1315),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1245),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1240),
.B(n_1245),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1266),
.A2(n_1256),
.B(n_1310),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1328),
.A2(n_1324),
.B1(n_1230),
.B2(n_1357),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1329),
.B(n_1340),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1237),
.Y(n_1384)
);

OAI22xp5_ASAP7_75t_L g1385 ( 
.A1(n_1340),
.A2(n_1343),
.B1(n_1266),
.B2(n_1253),
.Y(n_1385)
);

BUFx2_ASAP7_75t_SL g1386 ( 
.A(n_1238),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1328),
.A2(n_1343),
.B(n_1336),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1217),
.Y(n_1388)
);

INVx2_ASAP7_75t_SL g1389 ( 
.A(n_1238),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1229),
.A2(n_1336),
.B1(n_1354),
.B2(n_1318),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1229),
.A2(n_1354),
.B1(n_1276),
.B2(n_1335),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1246),
.Y(n_1392)
);

OAI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1335),
.A2(n_1351),
.B1(n_1232),
.B2(n_1303),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1351),
.A2(n_1222),
.B1(n_1358),
.B2(n_1273),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1262),
.B(n_1313),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1305),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1305),
.Y(n_1397)
);

AO21x1_ASAP7_75t_SL g1398 ( 
.A1(n_1256),
.A2(n_1301),
.B(n_1290),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1259),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1348),
.A2(n_1263),
.B1(n_1337),
.B2(n_1264),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1259),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1345),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1252),
.Y(n_1403)
);

BUFx2_ASAP7_75t_R g1404 ( 
.A(n_1287),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1260),
.Y(n_1405)
);

NAND2x1_ASAP7_75t_L g1406 ( 
.A(n_1280),
.B(n_1271),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1334),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1317),
.A2(n_1279),
.B(n_1304),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1274),
.B(n_1311),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1347),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1350),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1297),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1278),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1320),
.A2(n_1268),
.B(n_1304),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1301),
.B(n_1257),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1261),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1320),
.A2(n_1281),
.B(n_1270),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1242),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1257),
.A2(n_1264),
.B1(n_1214),
.B2(n_1220),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1214),
.A2(n_1220),
.B1(n_1355),
.B2(n_1353),
.Y(n_1420)
);

AOI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1279),
.A2(n_1281),
.B(n_1323),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1242),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1247),
.A2(n_1293),
.B(n_1244),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1300),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1242),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1321),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1269),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1228),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_1332),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1280),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1330),
.B(n_1361),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1321),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1309),
.A2(n_1235),
.B(n_1306),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1286),
.A2(n_1327),
.B(n_1338),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1316),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1283),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1326),
.A2(n_1355),
.B1(n_1353),
.B2(n_1331),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1255),
.B(n_1331),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1267),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1251),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1302),
.Y(n_1441)
);

BUFx12f_ASAP7_75t_L g1442 ( 
.A(n_1360),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1285),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1309),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1314),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1306),
.A2(n_1359),
.B(n_1361),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1330),
.A2(n_1275),
.B(n_1312),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1280),
.B(n_1284),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1308),
.Y(n_1449)
);

AO21x1_ASAP7_75t_SL g1450 ( 
.A1(n_1282),
.A2(n_1322),
.B(n_1296),
.Y(n_1450)
);

CKINVDCx12_ASAP7_75t_R g1451 ( 
.A(n_1248),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1291),
.B(n_1289),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1221),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1265),
.B(n_1299),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1277),
.B(n_1218),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1292),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1349),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1322),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1322),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1319),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1307),
.A2(n_1288),
.B(n_1248),
.Y(n_1462)
);

NAND2x1p5_ASAP7_75t_L g1463 ( 
.A(n_1307),
.B(n_1292),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1223),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1248),
.B(n_1223),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1298),
.A2(n_1295),
.B1(n_1288),
.B2(n_1294),
.Y(n_1466)
);

BUFx2_ASAP7_75t_R g1467 ( 
.A(n_1344),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1225),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1225),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1346),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1236),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1272),
.Y(n_1472)
);

INVx1_ASAP7_75t_SL g1473 ( 
.A(n_1349),
.Y(n_1473)
);

BUFx2_ASAP7_75t_R g1474 ( 
.A(n_1292),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1236),
.B(n_1258),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1258),
.A2(n_1341),
.B1(n_1216),
.B2(n_1206),
.Y(n_1476)
);

HB1xp67_ASAP7_75t_L g1477 ( 
.A(n_1246),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1279),
.A2(n_1247),
.B(n_1268),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1250),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1310),
.B(n_1276),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1238),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1249),
.A2(n_1206),
.B1(n_1155),
.B2(n_886),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1364),
.A2(n_1482),
.B1(n_1362),
.B2(n_1375),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1388),
.Y(n_1484)
);

OR2x6_ASAP7_75t_L g1485 ( 
.A(n_1406),
.B(n_1430),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1404),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1462),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1383),
.B(n_1367),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1480),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1388),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1409),
.B(n_1395),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1409),
.B(n_1395),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1383),
.B(n_1374),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1480),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1385),
.A2(n_1393),
.B1(n_1451),
.B2(n_1371),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1378),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1403),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1435),
.B(n_1424),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1392),
.Y(n_1499)
);

INVx4_ASAP7_75t_R g1500 ( 
.A(n_1403),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1435),
.B(n_1415),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1462),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1458),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1376),
.B(n_1438),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1408),
.A2(n_1414),
.B(n_1417),
.Y(n_1505)
);

AO21x2_ASAP7_75t_L g1506 ( 
.A1(n_1421),
.A2(n_1434),
.B(n_1387),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1369),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1366),
.B(n_1470),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1399),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1467),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1399),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1458),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1390),
.A2(n_1394),
.B(n_1391),
.Y(n_1513)
);

OR2x6_ASAP7_75t_L g1514 ( 
.A(n_1406),
.B(n_1430),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1401),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1441),
.A2(n_1381),
.B(n_1444),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1450),
.Y(n_1517)
);

BUFx3_ASAP7_75t_L g1518 ( 
.A(n_1429),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1476),
.A2(n_1400),
.B(n_1376),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1407),
.Y(n_1520)
);

INVxp67_ASAP7_75t_SL g1521 ( 
.A(n_1477),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1407),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1398),
.B(n_1396),
.Y(n_1523)
);

AND2x4_ASAP7_75t_L g1524 ( 
.A(n_1448),
.B(n_1363),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1398),
.B(n_1397),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1459),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1427),
.B(n_1405),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1410),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1397),
.B(n_1436),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1410),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1436),
.B(n_1411),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1433),
.A2(n_1426),
.B(n_1432),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1432),
.B(n_1412),
.Y(n_1533)
);

OA21x2_ASAP7_75t_L g1534 ( 
.A1(n_1418),
.A2(n_1425),
.B(n_1422),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1454),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1454),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1445),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1429),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1368),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1443),
.Y(n_1540)
);

BUFx3_ASAP7_75t_L g1541 ( 
.A(n_1413),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1447),
.A2(n_1446),
.B(n_1425),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1478),
.B(n_1418),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1446),
.A2(n_1447),
.B(n_1423),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1370),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1373),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1372),
.Y(n_1547)
);

CKINVDCx11_ASAP7_75t_R g1548 ( 
.A(n_1416),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1413),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1448),
.B(n_1384),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1419),
.B(n_1363),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1439),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1468),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1523),
.B(n_1449),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1496),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1523),
.B(n_1365),
.Y(n_1556)
);

AND2x4_ASAP7_75t_SL g1557 ( 
.A(n_1517),
.B(n_1365),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.B(n_1365),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1525),
.B(n_1479),
.Y(n_1559)
);

OR2x2_ASAP7_75t_SL g1560 ( 
.A(n_1517),
.B(n_1460),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1501),
.B(n_1382),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1532),
.B(n_1534),
.Y(n_1562)
);

AOI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1483),
.A2(n_1428),
.B1(n_1452),
.B2(n_1377),
.C(n_1455),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1495),
.B(n_1377),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1499),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1532),
.B(n_1450),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1532),
.B(n_1377),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1543),
.Y(n_1568)
);

AOI33xp33_ASAP7_75t_R g1569 ( 
.A1(n_1540),
.A2(n_1451),
.A3(n_1474),
.B1(n_1453),
.B2(n_1442),
.B3(n_1472),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1501),
.B(n_1440),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1517),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1487),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1516),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1498),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1516),
.Y(n_1576)
);

NAND2x1_ASAP7_75t_L g1577 ( 
.A(n_1485),
.B(n_1481),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1513),
.A2(n_1386),
.B(n_1380),
.C(n_1465),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1491),
.B(n_1379),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1491),
.B(n_1379),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1492),
.B(n_1463),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1492),
.B(n_1469),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1498),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1506),
.B(n_1469),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1502),
.B(n_1431),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1550),
.B(n_1529),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1550),
.B(n_1471),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1565),
.B(n_1521),
.Y(n_1588)
);

OAI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1569),
.A2(n_1519),
.B1(n_1508),
.B2(n_1504),
.C(n_1490),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1565),
.B(n_1535),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1575),
.B(n_1536),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1569),
.A2(n_1484),
.B1(n_1549),
.B2(n_1541),
.C(n_1527),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1586),
.B(n_1524),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1586),
.B(n_1524),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1556),
.B(n_1489),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1555),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1564),
.A2(n_1551),
.B1(n_1541),
.B2(n_1549),
.Y(n_1597)
);

OAI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1563),
.A2(n_1473),
.B1(n_1493),
.B2(n_1488),
.C(n_1437),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1575),
.B(n_1539),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1583),
.B(n_1545),
.Y(n_1600)
);

OAI21xp33_ASAP7_75t_L g1601 ( 
.A1(n_1563),
.A2(n_1564),
.B(n_1578),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1555),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1570),
.B(n_1547),
.Y(n_1604)
);

NAND3xp33_ASAP7_75t_L g1605 ( 
.A(n_1578),
.B(n_1551),
.C(n_1533),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1579),
.B(n_1509),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1558),
.B(n_1494),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1558),
.B(n_1494),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1580),
.B(n_1511),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1577),
.A2(n_1485),
.B(n_1514),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1533),
.C(n_1553),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1559),
.B(n_1503),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1580),
.B(n_1511),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1515),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1571),
.A2(n_1485),
.B(n_1514),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1587),
.B(n_1581),
.Y(n_1616)
);

NAND4xp25_ASAP7_75t_L g1617 ( 
.A(n_1584),
.B(n_1552),
.C(n_1518),
.D(n_1538),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1567),
.B(n_1554),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1510),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1582),
.B(n_1529),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1567),
.B(n_1512),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1585),
.B(n_1507),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1574),
.B(n_1531),
.C(n_1546),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1624)
);

OAI21xp33_ASAP7_75t_L g1625 ( 
.A1(n_1561),
.A2(n_1507),
.B(n_1531),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_SL g1626 ( 
.A(n_1577),
.B(n_1486),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1560),
.A2(n_1518),
.B1(n_1538),
.B2(n_1497),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1567),
.B(n_1512),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1576),
.B(n_1522),
.C(n_1528),
.Y(n_1630)
);

OA21x2_ASAP7_75t_L g1631 ( 
.A1(n_1573),
.A2(n_1505),
.B(n_1544),
.Y(n_1631)
);

NAND4xp25_ASAP7_75t_L g1632 ( 
.A(n_1584),
.B(n_1497),
.C(n_1530),
.D(n_1520),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1561),
.A2(n_1514),
.B1(n_1485),
.B2(n_1420),
.C(n_1465),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1554),
.B(n_1526),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1596),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1596),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1602),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1602),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1631),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1618),
.B(n_1562),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_SL g1641 ( 
.A(n_1601),
.B(n_1571),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1621),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1631),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1603),
.B(n_1562),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1600),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1630),
.B(n_1577),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1593),
.B(n_1594),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1604),
.Y(n_1649)
);

BUFx2_ASAP7_75t_L g1650 ( 
.A(n_1615),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1588),
.B(n_1568),
.Y(n_1651)
);

BUFx2_ASAP7_75t_L g1652 ( 
.A(n_1615),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1566),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1606),
.B(n_1573),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1629),
.B(n_1566),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1595),
.B(n_1566),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1591),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1609),
.B(n_1584),
.Y(n_1658)
);

NAND4xp25_ASAP7_75t_L g1659 ( 
.A(n_1601),
.B(n_1457),
.C(n_1461),
.D(n_1561),
.Y(n_1659)
);

AND2x2_ASAP7_75t_SL g1660 ( 
.A(n_1634),
.B(n_1557),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1623),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1614),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1642),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

INVxp67_ASAP7_75t_SL g1666 ( 
.A(n_1635),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_1607),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1653),
.B(n_1655),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1636),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1637),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1655),
.B(n_1608),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1635),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1654),
.B(n_1616),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1635),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1638),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1654),
.B(n_1590),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1655),
.B(n_1608),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1660),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1572),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1642),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1638),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1641),
.A2(n_1597),
.B(n_1605),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1654),
.B(n_1661),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1645),
.B(n_1612),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1640),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1643),
.B(n_1624),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1646),
.B(n_1628),
.Y(n_1691)
);

NAND4xp25_ASAP7_75t_L g1692 ( 
.A(n_1641),
.B(n_1589),
.C(n_1592),
.D(n_1598),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1638),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1638),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1651),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1651),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_L g1697 ( 
.A(n_1657),
.B(n_1486),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1639),
.Y(n_1698)
);

NAND2xp33_ASAP7_75t_R g1699 ( 
.A(n_1650),
.B(n_1548),
.Y(n_1699)
);

NOR2x1p5_ASAP7_75t_L g1700 ( 
.A(n_1659),
.B(n_1617),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1639),
.Y(n_1701)
);

AND2x4_ASAP7_75t_SL g1702 ( 
.A(n_1663),
.B(n_1571),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1665),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1665),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1674),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1686),
.B(n_1661),
.Y(n_1706)
);

INVxp67_ASAP7_75t_SL g1707 ( 
.A(n_1674),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1669),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1700),
.B(n_1661),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1685),
.A2(n_1692),
.B(n_1697),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1668),
.B(n_1650),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1661),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1681),
.B(n_1650),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1686),
.B(n_1695),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1669),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1676),
.Y(n_1716)
);

NAND2x1_ASAP7_75t_L g1717 ( 
.A(n_1682),
.B(n_1652),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1695),
.B(n_1651),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1681),
.B(n_1652),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1676),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1685),
.B(n_1681),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1676),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1682),
.B(n_1626),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1683),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1670),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1689),
.B(n_1657),
.Y(n_1727)
);

NOR3xp33_ASAP7_75t_L g1728 ( 
.A(n_1692),
.B(n_1659),
.C(n_1652),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1668),
.B(n_1656),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1682),
.B(n_1626),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1682),
.B(n_1633),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1656),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1679),
.A2(n_1625),
.B1(n_1622),
.B2(n_1632),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1684),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1648),
.Y(n_1735)
);

NAND2x1p5_ASAP7_75t_L g1736 ( 
.A(n_1696),
.B(n_1660),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1670),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1679),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1689),
.B(n_1649),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1664),
.B(n_1656),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1675),
.B(n_1658),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1690),
.B(n_1649),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1664),
.B(n_1640),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1667),
.B(n_1640),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1714),
.B(n_1675),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1710),
.A2(n_1699),
.B1(n_1660),
.B2(n_1627),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1716),
.Y(n_1747)
);

NAND2x1_ASAP7_75t_SL g1748 ( 
.A(n_1713),
.B(n_1644),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1703),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1706),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1736),
.B(n_1667),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1728),
.A2(n_1625),
.B1(n_1610),
.B2(n_1660),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1724),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1716),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1703),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1706),
.Y(n_1756)
);

INVxp67_ASAP7_75t_L g1757 ( 
.A(n_1709),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1714),
.B(n_1690),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1704),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1705),
.Y(n_1761)
);

BUFx3_ASAP7_75t_L g1762 ( 
.A(n_1717),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1672),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1736),
.B(n_1672),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1720),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1691),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1738),
.B(n_1691),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1735),
.B(n_1680),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1721),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1741),
.B(n_1671),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1715),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1741),
.B(n_1671),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1727),
.B(n_1680),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1735),
.B(n_1687),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1735),
.B(n_1687),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1715),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1726),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1711),
.B(n_1740),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1713),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1742),
.B(n_1662),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1749),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1749),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1755),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1748),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_SL g1785 ( 
.A(n_1769),
.B(n_1731),
.C(n_1717),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1750),
.B(n_1739),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1755),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1778),
.B(n_1711),
.Y(n_1788)
);

AOI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1757),
.A2(n_1707),
.B(n_1730),
.C(n_1723),
.Y(n_1789)
);

OAI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1746),
.A2(n_1733),
.B(n_1719),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1753),
.B(n_1740),
.Y(n_1791)
);

AOI221xp5_ASAP7_75t_L g1792 ( 
.A1(n_1761),
.A2(n_1756),
.B1(n_1779),
.B2(n_1766),
.C(n_1752),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1748),
.Y(n_1793)
);

AOI31xp33_ASAP7_75t_L g1794 ( 
.A1(n_1767),
.A2(n_1713),
.A3(n_1719),
.B(n_1500),
.Y(n_1794)
);

AOI22xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1761),
.A2(n_1719),
.B1(n_1702),
.B2(n_1729),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1778),
.B(n_1729),
.Y(n_1796)
);

AOI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1762),
.A2(n_1726),
.B(n_1708),
.C(n_1737),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1762),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1762),
.B(n_1732),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1759),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1768),
.B(n_1732),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1751),
.A2(n_1702),
.B(n_1611),
.C(n_1619),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1768),
.B(n_1743),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1774),
.B(n_1743),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1759),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1774),
.B(n_1744),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1781),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1788),
.B(n_1775),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1782),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1788),
.B(n_1760),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1791),
.B(n_1745),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1792),
.B(n_1775),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1798),
.B(n_1760),
.Y(n_1813)
);

AO22x1_ASAP7_75t_L g1814 ( 
.A1(n_1784),
.A2(n_1763),
.B1(n_1764),
.B2(n_1751),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1783),
.Y(n_1815)
);

NAND2x1_ASAP7_75t_SL g1816 ( 
.A(n_1799),
.B(n_1763),
.Y(n_1816)
);

OAI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1785),
.A2(n_1745),
.B1(n_1758),
.B2(n_1773),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1799),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1798),
.B(n_1787),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1800),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1799),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1805),
.B(n_1771),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1803),
.B(n_1764),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1796),
.B(n_1801),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1797),
.B(n_1771),
.Y(n_1825)
);

NAND2x1_ASAP7_75t_L g1826 ( 
.A(n_1784),
.B(n_1793),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1803),
.B(n_1744),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1817),
.A2(n_1790),
.B1(n_1789),
.B2(n_1794),
.C(n_1802),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1818),
.B(n_1804),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1825),
.A2(n_1802),
.B(n_1786),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1825),
.A2(n_1793),
.B(n_1806),
.Y(n_1831)
);

NOR4xp25_ASAP7_75t_L g1832 ( 
.A(n_1812),
.B(n_1777),
.C(n_1776),
.D(n_1754),
.Y(n_1832)
);

NAND4xp75_ASAP7_75t_L g1833 ( 
.A(n_1821),
.B(n_1804),
.C(n_1777),
.D(n_1776),
.Y(n_1833)
);

AOI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1814),
.A2(n_1795),
.B1(n_1806),
.B2(n_1754),
.C(n_1765),
.Y(n_1834)
);

AOI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1807),
.A2(n_1806),
.B1(n_1747),
.B2(n_1765),
.C(n_1754),
.Y(n_1835)
);

OAI21xp33_ASAP7_75t_L g1836 ( 
.A1(n_1816),
.A2(n_1758),
.B(n_1770),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1810),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1811),
.A2(n_1780),
.B1(n_1772),
.B2(n_1770),
.C(n_1765),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1823),
.A2(n_1780),
.B1(n_1747),
.B2(n_1772),
.Y(n_1839)
);

O2A1O1Ixp5_ASAP7_75t_L g1840 ( 
.A1(n_1826),
.A2(n_1747),
.B(n_1722),
.C(n_1734),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1830),
.B(n_1808),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1828),
.B(n_1819),
.C(n_1813),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_L g1843 ( 
.A(n_1831),
.B(n_1819),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1829),
.B(n_1827),
.Y(n_1844)
);

OAI211xp5_ASAP7_75t_SL g1845 ( 
.A1(n_1834),
.A2(n_1824),
.B(n_1813),
.C(n_1820),
.Y(n_1845)
);

NOR2x1_ASAP7_75t_L g1846 ( 
.A(n_1833),
.B(n_1809),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1832),
.B(n_1815),
.C(n_1810),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1837),
.B(n_1442),
.Y(n_1848)
);

NOR2x1_ASAP7_75t_L g1849 ( 
.A(n_1838),
.B(n_1822),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1839),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1836),
.A2(n_1840),
.B(n_1835),
.Y(n_1851)
);

NOR2x1_ASAP7_75t_L g1852 ( 
.A(n_1843),
.B(n_1822),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1846),
.Y(n_1853)
);

NOR3x1_ASAP7_75t_L g1854 ( 
.A(n_1842),
.B(n_1718),
.C(n_1725),
.Y(n_1854)
);

AOI221x1_ASAP7_75t_L g1855 ( 
.A1(n_1847),
.A2(n_1734),
.B1(n_1722),
.B2(n_1720),
.C(n_1701),
.Y(n_1855)
);

NAND4xp25_ASAP7_75t_SL g1856 ( 
.A(n_1851),
.B(n_1841),
.C(n_1849),
.D(n_1850),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1844),
.B(n_1718),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1857),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1852),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1853),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1854),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1855),
.Y(n_1862)
);

AO22x1_ASAP7_75t_L g1863 ( 
.A1(n_1856),
.A2(n_1848),
.B1(n_1845),
.B2(n_1461),
.Y(n_1863)
);

HB1xp67_ASAP7_75t_L g1864 ( 
.A(n_1853),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1864),
.Y(n_1865)
);

NAND4xp75_ASAP7_75t_L g1866 ( 
.A(n_1860),
.B(n_1389),
.C(n_1456),
.D(n_1701),
.Y(n_1866)
);

NOR2xp67_ASAP7_75t_L g1867 ( 
.A(n_1864),
.B(n_1457),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1861),
.B(n_1369),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1859),
.B(n_1725),
.Y(n_1869)
);

NAND3x2_ASAP7_75t_L g1870 ( 
.A(n_1858),
.B(n_1402),
.C(n_1646),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1868),
.B(n_1863),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1865),
.Y(n_1872)
);

NAND3x1_ASAP7_75t_L g1873 ( 
.A(n_1867),
.B(n_1862),
.C(n_1402),
.Y(n_1873)
);

HB1xp67_ASAP7_75t_L g1874 ( 
.A(n_1872),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_SL g1875 ( 
.A1(n_1874),
.A2(n_1862),
.B(n_1869),
.Y(n_1875)
);

NOR2x1p5_ASAP7_75t_L g1876 ( 
.A(n_1875),
.B(n_1871),
.Y(n_1876)
);

AO21x2_ASAP7_75t_L g1877 ( 
.A1(n_1875),
.A2(n_1873),
.B(n_1870),
.Y(n_1877)
);

AOI22xp5_ASAP7_75t_L g1878 ( 
.A1(n_1876),
.A2(n_1877),
.B1(n_1866),
.B2(n_1701),
.Y(n_1878)
);

AOI221xp5_ASAP7_75t_L g1879 ( 
.A1(n_1877),
.A2(n_1698),
.B1(n_1666),
.B2(n_1466),
.C(n_1677),
.Y(n_1879)
);

AO21x1_ASAP7_75t_L g1880 ( 
.A1(n_1878),
.A2(n_1698),
.B(n_1666),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1879),
.A2(n_1698),
.B1(n_1678),
.B2(n_1677),
.C(n_1673),
.Y(n_1881)
);

AOI222xp33_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1673),
.B1(n_1694),
.B2(n_1678),
.C1(n_1693),
.C2(n_1684),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1882),
.A2(n_1880),
.B1(n_1386),
.B2(n_1644),
.Y(n_1883)
);

AOI221xp5_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1694),
.B1(n_1693),
.B2(n_1684),
.C(n_1389),
.Y(n_1884)
);

AOI211xp5_ASAP7_75t_L g1885 ( 
.A1(n_1884),
.A2(n_1456),
.B(n_1475),
.C(n_1464),
.Y(n_1885)
);


endmodule