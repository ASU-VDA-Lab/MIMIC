module fake_jpeg_7482_n_33 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_33);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_33;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_2),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_SL g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_16),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_7),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_15)
);

AO21x2_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_13),
.B(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_18),
.B(n_15),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_11),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_28),
.C(n_13),
.Y(n_31)
);

AOI322xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_6),
.A3(n_8),
.B1(n_12),
.B2(n_14),
.C1(n_16),
.C2(n_29),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_8),
.Y(n_33)
);


endmodule