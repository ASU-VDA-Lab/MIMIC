module fake_jpeg_31189_n_414 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_414);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_414;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_56),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

AOI21xp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_9),
.B(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_23),
.B(n_9),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_65),
.Y(n_95)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_77),
.Y(n_106)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_22),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_33),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_33),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_22),
.B(n_8),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_24),
.B(n_19),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_82),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_47),
.B1(n_37),
.B2(n_21),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_38),
.B1(n_54),
.B2(n_53),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_48),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_24),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_23),
.B1(n_46),
.B2(n_45),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_110),
.A2(n_47),
.B1(n_29),
.B2(n_46),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_121),
.Y(n_135)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_33),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_29),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_29),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_87),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_147),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_144),
.Y(n_164)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_142),
.B1(n_151),
.B2(n_154),
.Y(n_176)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_152),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_100),
.A2(n_38),
.B1(n_21),
.B2(n_25),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_97),
.A2(n_82),
.B1(n_50),
.B2(n_55),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_143),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_95),
.B(n_74),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_31),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_31),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g147 ( 
.A(n_91),
.B(n_67),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_99),
.B(n_58),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_149),
.B(n_162),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_94),
.A2(n_38),
.B1(n_87),
.B2(n_41),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_157),
.B1(n_159),
.B2(n_26),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_104),
.A2(n_61),
.B1(n_57),
.B2(n_64),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_89),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_88),
.A2(n_69),
.B1(n_41),
.B2(n_81),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_96),
.A2(n_112),
.B(n_85),
.C(n_47),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_155),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_118),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_158),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_98),
.A2(n_83),
.B1(n_73),
.B2(n_72),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_189),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_106),
.B(n_26),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_168),
.B(n_178),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g171 ( 
.A(n_144),
.B(n_102),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_179),
.B1(n_171),
.B2(n_134),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_30),
.C(n_46),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_183),
.A2(n_21),
.B(n_31),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_154),
.A2(n_103),
.B1(n_92),
.B2(n_117),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_147),
.B1(n_150),
.B2(n_92),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_45),
.A3(n_30),
.B1(n_42),
.B2(n_35),
.Y(n_189)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_181),
.A2(n_157),
.B1(n_148),
.B2(n_159),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_206),
.B1(n_203),
.B2(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_165),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_208),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_105),
.B1(n_140),
.B2(n_141),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_135),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_202),
.B(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_206),
.B1(n_198),
.B2(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_147),
.C(n_131),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_173),
.C(n_183),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_155),
.B(n_152),
.C(n_147),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_205),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_151),
.B1(n_131),
.B2(n_117),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_189),
.B(n_137),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_136),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_214),
.B(n_170),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_109),
.B1(n_103),
.B2(n_155),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_173),
.B1(n_170),
.B2(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_133),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_232),
.C(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_219),
.B(n_220),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_234),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_226),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_212),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_230),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_174),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_173),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_180),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_203),
.A2(n_180),
.B1(n_133),
.B2(n_153),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_109),
.B1(n_175),
.B2(n_162),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_197),
.B1(n_194),
.B2(n_175),
.Y(n_263)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

NAND3xp33_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_201),
.C(n_198),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_256),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_208),
.B(n_199),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_223),
.B(n_217),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_242),
.Y(n_266)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_257),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_232),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_137),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_261),
.C(n_229),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_213),
.B1(n_205),
.B2(n_193),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_263),
.B1(n_216),
.B2(n_192),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_193),
.Y(n_254)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_255),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_259),
.Y(n_291)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_205),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_262),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_209),
.C(n_210),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_169),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_252),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_270),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_232),
.C(n_229),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_273),
.C(n_282),
.Y(n_293)
);

AOI22x1_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_217),
.B1(n_227),
.B2(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_209),
.C(n_216),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_264),
.B1(n_256),
.B2(n_259),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_277),
.B1(n_185),
.B2(n_177),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_276),
.A2(n_283),
.B1(n_188),
.B2(n_190),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_211),
.B1(n_192),
.B2(n_191),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_243),
.B(n_210),
.C(n_186),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_245),
.A2(n_211),
.B1(n_192),
.B2(n_188),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_263),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_238),
.A2(n_211),
.B(n_129),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_292),
.B(n_248),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_247),
.B(n_30),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_243),
.B(n_177),
.C(n_185),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_156),
.C(n_158),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_238),
.A2(n_143),
.B(n_161),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_290),
.A2(n_258),
.B1(n_241),
.B2(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_294),
.A2(n_295),
.B1(n_302),
.B2(n_303),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_276),
.A2(n_242),
.B1(n_239),
.B2(n_246),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_297),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_298),
.B(n_310),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_260),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_300),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_255),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_301),
.B(n_311),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_188),
.B1(n_182),
.B2(n_169),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_285),
.B1(n_280),
.B2(n_279),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_288),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_305),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_306),
.B(n_313),
.C(n_314),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_267),
.A2(n_182),
.B1(n_163),
.B2(n_160),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_308),
.A2(n_277),
.B1(n_278),
.B2(n_274),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_292),
.A2(n_145),
.B(n_6),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_132),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_282),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_105),
.C(n_124),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_124),
.C(n_128),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_288),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_316),
.B(n_272),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_296),
.A2(n_283),
.B1(n_265),
.B2(n_266),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_318),
.A2(n_320),
.B1(n_335),
.B2(n_336),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_299),
.Y(n_321)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_328),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_324),
.A2(n_329),
.B1(n_315),
.B2(n_305),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_326),
.B(n_331),
.Y(n_346)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_289),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_281),
.B1(n_278),
.B2(n_268),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_272),
.C(n_291),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_332),
.C(n_306),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_268),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_291),
.C(n_127),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_300),
.B(n_132),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_301),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_309),
.A2(n_108),
.B1(n_37),
.B2(n_123),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_309),
.A2(n_25),
.B1(n_35),
.B2(n_42),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_354),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_323),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_343),
.B(n_345),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_314),
.C(n_313),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_352),
.C(n_355),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_331),
.B(n_312),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_347),
.B(n_348),
.Y(n_364)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_349),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_303),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_350),
.B(n_344),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_13),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_351),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_319),
.C(n_325),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_338),
.A2(n_317),
.B1(n_337),
.B2(n_326),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_70),
.C(n_42),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_35),
.C(n_25),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_356),
.B(n_0),
.C(n_1),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_364),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_352),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_359),
.B(n_360),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_341),
.A2(n_330),
.B(n_342),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_353),
.A2(n_333),
.B1(n_335),
.B2(n_102),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_361),
.A2(n_369),
.B1(n_360),
.B2(n_370),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_356),
.B(n_10),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_363),
.B(n_367),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_10),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_355),
.A2(n_10),
.B(n_18),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_368),
.B(n_370),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_372),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_339),
.C(n_346),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_377),
.B(n_15),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_339),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_374),
.B(n_379),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_366),
.B(n_348),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_376),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_358),
.B(n_11),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_11),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_365),
.B(n_8),
.Y(n_380)
);

AOI21x1_ASAP7_75t_L g393 ( 
.A1(n_380),
.A2(n_0),
.B(n_2),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_365),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_381),
.A2(n_115),
.B1(n_49),
.B2(n_7),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_371),
.A2(n_361),
.B(n_12),
.Y(n_384)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_382),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_385),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_386),
.B(n_387),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_373),
.A2(n_18),
.B1(n_15),
.B2(n_14),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_372),
.A2(n_14),
.B(n_15),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_389),
.Y(n_394)
);

INVx11_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_393),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_385),
.A2(n_374),
.B(n_2),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_396),
.A2(n_2),
.B(n_3),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_0),
.Y(n_399)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_399),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

A2O1A1O1Ixp25_ASAP7_75t_L g402 ( 
.A1(n_395),
.A2(n_392),
.B(n_383),
.C(n_391),
.D(n_5),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_401),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_397),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_394),
.A2(n_392),
.B(n_4),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_396),
.C(n_400),
.Y(n_408)
);

AOI21x1_ASAP7_75t_L g411 ( 
.A1(n_407),
.A2(n_409),
.B(n_3),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_408),
.A2(n_404),
.B1(n_403),
.B2(n_398),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_410),
.A2(n_411),
.B(n_4),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_412),
.A2(n_5),
.B(n_298),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_413),
.B(n_5),
.Y(n_414)
);


endmodule