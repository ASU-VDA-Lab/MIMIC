module fake_jpeg_27146_n_48 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_48);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_48;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx8_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_22),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_29),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_24),
.B(n_19),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_30),
.B(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_36),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_18),
.C(n_11),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_2),
.C(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_35),
.B1(n_32),
.B2(n_4),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_38),
.C(n_39),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_44),
.B(n_42),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_38),
.C(n_43),
.Y(n_46)
);

OAI321xp33_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_2),
.A3(n_3),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_R g48 ( 
.A1(n_47),
.A2(n_6),
.B1(n_12),
.B2(n_13),
.Y(n_48)
);


endmodule