module fake_jpeg_14991_n_217 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_49),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_41),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_1),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_48),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_18),
.B(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_28),
.B1(n_24),
.B2(n_21),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_51),
.A2(n_74),
.B1(n_29),
.B2(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_24),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_69),
.Y(n_100)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_28),
.B1(n_21),
.B2(n_33),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_71),
.B1(n_34),
.B2(n_48),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_28),
.B1(n_21),
.B2(n_26),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_27),
.B(n_33),
.C(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_38),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_45),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_80),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_42),
.B1(n_44),
.B2(n_37),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_79),
.A2(n_83),
.B1(n_66),
.B2(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_57),
.B(n_49),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_29),
.B(n_2),
.C(n_3),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_44),
.B1(n_42),
.B2(n_37),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_23),
.B1(n_34),
.B2(n_31),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_25),
.B(n_3),
.Y(n_120)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_91),
.Y(n_122)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_30),
.B1(n_19),
.B2(n_47),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_92),
.B1(n_97),
.B2(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_35),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_102),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_50),
.B(n_47),
.C(n_35),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_47),
.C(n_26),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_35),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_25),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_116),
.C(n_81),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_107),
.B(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_84),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_63),
.B1(n_56),
.B2(n_53),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_113),
.B1(n_126),
.B2(n_127),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_47),
.B(n_26),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_81),
.B(n_104),
.C(n_96),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_101),
.B1(n_89),
.B2(n_8),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_2),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_76),
.B(n_95),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_4),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_100),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_87),
.A2(n_25),
.B1(n_16),
.B2(n_14),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_16),
.B1(n_13),
.B2(n_7),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_118),
.A2(n_96),
.B1(n_85),
.B2(n_88),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_131),
.B1(n_137),
.B2(n_141),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_96),
.B1(n_77),
.B2(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_132),
.B(n_140),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_134),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_143),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_105),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_111),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_117),
.B(n_120),
.Y(n_152)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_104),
.B1(n_94),
.B2(n_91),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_145),
.B(n_109),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_5),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_108),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_152),
.B(n_131),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_151),
.B(n_157),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_163),
.C(n_128),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_125),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_165),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_116),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_128),
.A2(n_140),
.A3(n_132),
.B1(n_138),
.B2(n_143),
.C1(n_146),
.C2(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_124),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_117),
.C(n_112),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_121),
.C(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_168),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_141),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_131),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_131),
.B1(n_145),
.B2(n_123),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_177),
.B1(n_179),
.B2(n_157),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_136),
.C(n_133),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_175),
.B(n_180),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_126),
.C(n_113),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_107),
.B(n_145),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_157),
.A2(n_154),
.B(n_151),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_178),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_131),
.B1(n_127),
.B2(n_123),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_169),
.A2(n_164),
.B1(n_160),
.B2(n_158),
.Y(n_182)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_155),
.C(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_190),
.C(n_191),
.Y(n_192)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_189),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_150),
.Y(n_199)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_153),
.C(n_159),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_187),
.A2(n_186),
.B(n_183),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_196),
.B(n_197),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_183),
.A2(n_167),
.B(n_180),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_190),
.A2(n_159),
.B(n_176),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_170),
.C(n_153),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_202),
.Y(n_209)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_184),
.C(n_181),
.Y(n_203)
);

AOI21x1_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_5),
.B(n_6),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_150),
.Y(n_205)
);

OAI221xp5_ASAP7_75t_L g208 ( 
.A1(n_205),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_203),
.Y(n_208)
);

AOI31xp67_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_182),
.A3(n_191),
.B(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_206),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_10),
.B(n_11),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_210),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_9),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_209),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_215),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_213),
.Y(n_217)
);


endmodule