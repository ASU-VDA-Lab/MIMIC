module real_aes_3759_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_1014;
wire n_329;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1016;
wire n_908;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_1021;
wire n_399;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_1025;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_817;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_1006;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_527;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_1031;
wire n_432;
wire n_880;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_927;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_637;
wire n_526;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_721;
wire n_446;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_967;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_0), .A2(n_168), .B1(n_439), .B2(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_1), .Y(n_309) );
AND2x4_ASAP7_75t_L g783 ( .A(n_1), .B(n_784), .Y(n_783) );
AND2x4_ASAP7_75t_L g791 ( .A(n_1), .B(n_289), .Y(n_791) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_2), .A2(n_1025), .B1(n_1026), .B2(n_1028), .Y(n_1024) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_2), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_3), .A2(n_30), .B1(n_440), .B2(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g480 ( .A(n_4), .Y(n_480) );
INVx1_ASAP7_75t_L g550 ( .A(n_5), .Y(n_550) );
AO22x1_ASAP7_75t_L g826 ( .A1(n_5), .A2(n_7), .B1(n_790), .B2(n_808), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_6), .A2(n_246), .B1(n_490), .B2(n_491), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_8), .A2(n_217), .B1(n_780), .B2(n_787), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_9), .A2(n_111), .B1(n_442), .B2(n_507), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_10), .A2(n_226), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_11), .A2(n_258), .B1(n_534), .B2(n_568), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_12), .A2(n_57), .B1(n_442), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g597 ( .A(n_13), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_14), .A2(n_92), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_15), .A2(n_278), .B1(n_484), .B2(n_486), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_16), .A2(n_33), .B1(n_467), .B2(n_469), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_17), .B(n_599), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_18), .A2(n_23), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_19), .A2(n_171), .B1(n_490), .B2(n_491), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_20), .A2(n_238), .B1(n_543), .B2(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_21), .B(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_22), .A2(n_143), .B1(n_494), .B2(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_24), .A2(n_65), .B1(n_376), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_25), .A2(n_138), .B1(n_636), .B2(n_637), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_26), .A2(n_132), .B1(n_453), .B2(n_455), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_27), .A2(n_219), .B1(n_543), .B2(n_574), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_28), .A2(n_53), .B1(n_344), .B2(n_398), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_29), .A2(n_133), .B1(n_381), .B2(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_31), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_32), .A2(n_129), .B1(n_817), .B2(n_832), .Y(n_831) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_34), .A2(n_41), .B1(n_475), .B2(n_521), .C(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_35), .A2(n_230), .B1(n_469), .B2(n_614), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_36), .A2(n_66), .B1(n_376), .B2(n_571), .Y(n_593) );
INVx1_ASAP7_75t_L g738 ( .A(n_37), .Y(n_738) );
INVx1_ASAP7_75t_L g646 ( .A(n_38), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_39), .A2(n_117), .B1(n_522), .B2(n_748), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_40), .A2(n_185), .B1(n_490), .B2(n_491), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_42), .A2(n_620), .B(n_621), .Y(n_619) );
XOR2x2_ASAP7_75t_L g316 ( .A(n_43), .B(n_317), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_44), .A2(n_155), .B1(n_487), .B2(n_620), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_45), .A2(n_239), .B1(n_524), .B2(n_525), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g1012 ( .A1(n_46), .A2(n_483), .B(n_1013), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_47), .A2(n_58), .B1(n_321), .B2(n_467), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_48), .A2(n_90), .B1(n_356), .B2(n_360), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_49), .A2(n_475), .B(n_478), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_50), .B(n_223), .Y(n_307) );
INVx1_ASAP7_75t_L g340 ( .A(n_50), .Y(n_340) );
INVxp67_ASAP7_75t_L g425 ( .A(n_50), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_51), .A2(n_173), .B1(n_507), .B2(n_532), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_52), .A2(n_95), .B1(n_376), .B2(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_54), .B(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_55), .A2(n_139), .B1(n_620), .B2(n_636), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_56), .A2(n_169), .B1(n_521), .B2(n_522), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_59), .A2(n_88), .B1(n_493), .B2(n_494), .Y(n_728) );
XNOR2x1_ASAP7_75t_L g608 ( .A(n_60), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_61), .B(n_325), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_62), .A2(n_100), .B1(n_444), .B2(n_445), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_63), .A2(n_273), .B1(n_509), .B2(n_510), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_64), .A2(n_205), .B1(n_393), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g723 ( .A(n_67), .Y(n_723) );
INVx1_ASAP7_75t_L g769 ( .A(n_68), .Y(n_769) );
INVx1_ASAP7_75t_L g699 ( .A(n_69), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_70), .A2(n_186), .B1(n_376), .B2(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_71), .A2(n_245), .B1(n_393), .B2(n_616), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_72), .A2(n_240), .B1(n_484), .B2(n_486), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_73), .A2(n_127), .B1(n_487), .B2(n_652), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_74), .A2(n_183), .B1(n_796), .B2(n_808), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_75), .A2(n_220), .B1(n_636), .B2(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g548 ( .A(n_76), .Y(n_548) );
INVx2_ASAP7_75t_L g304 ( .A(n_77), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_78), .A2(n_286), .B1(n_393), .B2(n_616), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_79), .A2(n_130), .B1(n_540), .B2(n_612), .Y(n_1000) );
INVx1_ASAP7_75t_L g365 ( .A(n_80), .Y(n_365) );
INVx1_ASAP7_75t_L g782 ( .A(n_81), .Y(n_782) );
AND2x4_ASAP7_75t_L g788 ( .A(n_81), .B(n_304), .Y(n_788) );
INVx1_ASAP7_75t_SL g830 ( .A(n_81), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_82), .A2(n_225), .B1(n_490), .B2(n_491), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_83), .A2(n_262), .B1(n_376), .B2(n_483), .Y(n_756) );
INVx1_ASAP7_75t_L g374 ( .A(n_84), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_85), .A2(n_261), .B1(n_391), .B2(n_397), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_86), .A2(n_207), .B1(n_467), .B2(n_469), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_87), .A2(n_184), .B1(n_381), .B2(n_450), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_89), .A2(n_199), .B1(n_790), .B2(n_792), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_91), .A2(n_253), .B1(n_486), .B2(n_487), .Y(n_485) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_93), .Y(n_325) );
XNOR2x2_ASAP7_75t_SL g628 ( .A(n_94), .B(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g1007 ( .A1(n_96), .A2(n_182), .B1(n_367), .B2(n_1008), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_97), .A2(n_201), .B1(n_401), .B2(n_447), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_98), .A2(n_294), .B1(n_637), .B2(n_693), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_99), .A2(n_210), .B1(n_393), .B2(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g765 ( .A(n_101), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_102), .A2(n_175), .B1(n_780), .B2(n_815), .Y(n_814) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_103), .A2(n_104), .B1(n_487), .B2(n_493), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_105), .A2(n_216), .B1(n_796), .B2(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_106), .A2(n_190), .B1(n_790), .B2(n_808), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_107), .B(n_576), .Y(n_1015) );
INVx1_ASAP7_75t_L g326 ( .A(n_108), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_108), .B(n_222), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_109), .A2(n_280), .B1(n_534), .B2(n_616), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_110), .A2(n_163), .B1(n_440), .B2(n_540), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_112), .A2(n_595), .B(n_596), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_113), .A2(n_194), .B1(n_540), .B2(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_114), .A2(n_177), .B1(n_406), .B2(n_1002), .Y(n_1001) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_115), .A2(n_181), .B1(n_780), .B2(n_785), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_116), .A2(n_166), .B1(n_376), .B2(n_571), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_118), .A2(n_264), .B1(n_650), .B2(n_651), .C(n_653), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_119), .A2(n_125), .B1(n_780), .B2(n_787), .Y(n_840) );
XNOR2x1_ASAP7_75t_L g682 ( .A(n_120), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g410 ( .A(n_121), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_122), .A2(n_142), .B1(n_509), .B2(n_510), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_123), .A2(n_251), .B1(n_381), .B2(n_576), .C(n_578), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_124), .A2(n_148), .B1(n_534), .B2(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g384 ( .A(n_126), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_128), .A2(n_224), .B1(n_778), .B2(n_785), .Y(n_777) );
XNOR2x1_ASAP7_75t_L g463 ( .A(n_129), .B(n_464), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_131), .A2(n_248), .B1(n_401), .B2(n_405), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_134), .A2(n_193), .B1(n_543), .B2(n_545), .Y(n_592) );
INVx1_ASAP7_75t_L g654 ( .A(n_135), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_136), .A2(n_279), .B1(n_780), .B2(n_787), .Y(n_823) );
INVx1_ASAP7_75t_L g473 ( .A(n_137), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_140), .A2(n_652), .B(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_141), .A2(n_269), .B1(n_693), .B2(n_697), .Y(n_763) );
INVx1_ASAP7_75t_L g690 ( .A(n_144), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_145), .A2(n_259), .B1(n_490), .B2(n_491), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_146), .A2(n_212), .B1(n_612), .B2(n_742), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_147), .A2(n_287), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_149), .A2(n_176), .B1(n_532), .B2(n_614), .Y(n_613) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_150), .B(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_151), .A2(n_154), .B1(n_543), .B2(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_152), .A2(n_381), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g641 ( .A(n_153), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_156), .A2(n_260), .B1(n_393), .B2(n_616), .Y(n_1004) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_157), .A2(n_252), .B1(n_320), .B2(n_343), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_158), .A2(n_198), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_159), .A2(n_195), .B1(n_450), .B2(n_519), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_160), .A2(n_277), .B1(n_787), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_161), .A2(n_209), .B1(n_367), .B2(n_376), .Y(n_623) );
INVx1_ASAP7_75t_L g664 ( .A(n_162), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_164), .B(n_414), .Y(n_685) );
INVx1_ASAP7_75t_L g622 ( .A(n_165), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_167), .A2(n_203), .B1(n_519), .B2(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g379 ( .A(n_170), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_172), .A2(n_187), .B1(n_636), .B2(n_637), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_174), .A2(n_270), .B1(n_493), .B2(n_494), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_178), .B(n_460), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_179), .A2(n_276), .B1(n_406), .B2(n_538), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_180), .A2(n_231), .B1(n_796), .B2(n_817), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_188), .A2(n_265), .B1(n_439), .B2(n_534), .Y(n_743) );
AO221x2_ASAP7_75t_L g825 ( .A1(n_189), .A2(n_249), .B1(n_780), .B2(n_815), .C(n_826), .Y(n_825) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_190), .B(n_1006), .Y(n_1005) );
INVxp67_ASAP7_75t_L g1017 ( .A(n_190), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_190), .A2(n_1024), .B1(n_1029), .B2(n_1031), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_191), .A2(n_250), .B1(n_620), .B2(n_707), .Y(n_706) );
OA22x2_ASAP7_75t_L g330 ( .A1(n_192), .A2(n_223), .B1(n_325), .B2(n_329), .Y(n_330) );
INVx1_ASAP7_75t_L g351 ( .A(n_192), .Y(n_351) );
INVx1_ASAP7_75t_L g579 ( .A(n_196), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_197), .A2(n_243), .B1(n_510), .B2(n_538), .Y(n_537) );
XOR2x2_ASAP7_75t_L g435 ( .A(n_199), .B(n_436), .Y(n_435) );
XNOR2x1_ASAP7_75t_L g582 ( .A(n_200), .B(n_583), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_202), .A2(n_208), .B1(n_490), .B2(n_491), .Y(n_731) );
INVx1_ASAP7_75t_SL g526 ( .A(n_204), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_204), .A2(n_283), .B1(n_792), .B2(n_796), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_206), .A2(n_244), .B1(n_417), .B2(n_545), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_211), .A2(n_275), .B1(n_693), .B2(n_697), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_213), .A2(n_282), .B1(n_507), .B2(n_512), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_214), .A2(n_241), .B1(n_484), .B2(n_486), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_215), .A2(n_221), .B1(n_493), .B2(n_494), .Y(n_760) );
INVx1_ASAP7_75t_L g770 ( .A(n_218), .Y(n_770) );
INVx1_ASAP7_75t_L g342 ( .A(n_222), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_222), .B(n_349), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_223), .A2(n_237), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_227), .B(n_705), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_228), .A2(n_254), .B1(n_398), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_229), .A2(n_272), .B1(n_532), .B2(n_614), .Y(n_1003) );
AOI221x1_ASAP7_75t_SL g735 ( .A1(n_232), .A2(n_235), .B1(n_381), .B2(n_736), .C(n_737), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_233), .A2(n_234), .B1(n_447), .B2(n_538), .Y(n_563) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_236), .A2(n_293), .B1(n_651), .B2(n_721), .C(n_722), .Y(n_720) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_237), .B(n_281), .Y(n_308) );
INVx1_ASAP7_75t_L g328 ( .A(n_237), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_242), .A2(n_256), .B1(n_417), .B2(n_426), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_247), .A2(n_477), .B(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_255), .A2(n_288), .B1(n_693), .B2(n_697), .Y(n_712) );
INVx1_ASAP7_75t_L g673 ( .A(n_257), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_263), .A2(n_285), .B1(n_510), .B2(n_538), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_266), .A2(n_268), .B1(n_356), .B2(n_442), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_267), .A2(n_290), .B1(n_344), .B2(n_439), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_271), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g1014 ( .A(n_274), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_281), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_284), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g784 ( .A(n_289), .Y(n_784) );
HB1xp67_ASAP7_75t_L g1034 ( .A(n_289), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_291), .A2(n_292), .B1(n_510), .B2(n_538), .Y(n_679) );
INVx1_ASAP7_75t_L g648 ( .A(n_295), .Y(n_648) );
AOI22x1_ASAP7_75t_L g559 ( .A1(n_296), .A2(n_560), .B1(n_561), .B2(n_580), .Y(n_559) );
INVx1_ASAP7_75t_L g580 ( .A(n_296), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_310), .B(n_773), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND3xp33_ASAP7_75t_L g301 ( .A(n_302), .B(n_305), .C(n_309), .Y(n_301) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_302), .B(n_1021), .Y(n_1020) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_302), .B(n_1022), .Y(n_1030) );
AOI21xp5_ASAP7_75t_L g1035 ( .A1(n_302), .A2(n_309), .B(n_830), .Y(n_1035) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AO21x1_ASAP7_75t_L g1032 ( .A1(n_303), .A2(n_1033), .B(n_1035), .Y(n_1032) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g781 ( .A(n_304), .B(n_782), .Y(n_781) );
AND3x4_ASAP7_75t_L g829 ( .A(n_304), .B(n_783), .C(n_830), .Y(n_829) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_305), .B(n_1022), .Y(n_1021) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AO21x2_ASAP7_75t_L g429 ( .A1(n_306), .A2(n_430), .B(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g1022 ( .A(n_309), .Y(n_1022) );
XNOR2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_659), .Y(n_310) );
XNOR2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_496), .Y(n_311) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_433), .B2(n_495), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND4xp75_ASAP7_75t_L g317 ( .A(n_318), .B(n_363), .C(n_389), .D(n_408), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_355), .Y(n_318) );
BUFx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_321), .Y(n_442) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_321), .Y(n_469) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_321), .Y(n_532) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_321), .Y(n_742) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_331), .Y(n_321) );
AND2x2_ASAP7_75t_L g357 ( .A(n_322), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g388 ( .A(n_322), .B(n_383), .Y(n_388) );
AND2x2_ASAP7_75t_L g415 ( .A(n_322), .B(n_371), .Y(n_415) );
AND2x2_ASAP7_75t_L g468 ( .A(n_322), .B(n_358), .Y(n_468) );
AND2x2_ASAP7_75t_L g477 ( .A(n_322), .B(n_371), .Y(n_477) );
AND2x4_ASAP7_75t_L g486 ( .A(n_322), .B(n_383), .Y(n_486) );
AND2x4_ASAP7_75t_L g636 ( .A(n_322), .B(n_358), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_322), .B(n_354), .Y(n_637) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_330), .Y(n_322) );
INVx1_ASAP7_75t_L g370 ( .A(n_323), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_327), .Y(n_323) );
NAND2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx2_ASAP7_75t_L g329 ( .A(n_325), .Y(n_329) );
INVx3_ASAP7_75t_L g335 ( .A(n_325), .Y(n_335) );
NAND2xp33_ASAP7_75t_L g341 ( .A(n_325), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g353 ( .A(n_325), .Y(n_353) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_325), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_326), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g424 ( .A1(n_328), .A2(n_353), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g369 ( .A(n_330), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g396 ( .A(n_330), .Y(n_396) );
AND2x2_ASAP7_75t_L g423 ( .A(n_330), .B(n_424), .Y(n_423) );
AND2x4_ASAP7_75t_L g493 ( .A(n_331), .B(n_395), .Y(n_493) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_337), .Y(n_332) );
AND2x4_ASAP7_75t_L g358 ( .A(n_333), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g372 ( .A(n_333), .Y(n_372) );
AND2x4_ASAP7_75t_L g383 ( .A(n_333), .B(n_373), .Y(n_383) );
AND2x2_ASAP7_75t_L g419 ( .A(n_333), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_335), .B(n_340), .Y(n_339) );
INVxp67_ASAP7_75t_L g349 ( .A(n_335), .Y(n_349) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_336), .B(n_348), .C(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
BUFx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g586 ( .A(n_345), .Y(n_586) );
INVx5_ASAP7_75t_L g612 ( .A(n_345), .Y(n_612) );
INVx3_ASAP7_75t_L g633 ( .A(n_345), .Y(n_633) );
INVx6_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx12f_ASAP7_75t_L g440 ( .A(n_346), .Y(n_440) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_354), .Y(n_346) );
AND2x4_ASAP7_75t_L g362 ( .A(n_347), .B(n_358), .Y(n_362) );
AND2x4_ASAP7_75t_L g377 ( .A(n_347), .B(n_371), .Y(n_377) );
AND2x4_ASAP7_75t_L g487 ( .A(n_347), .B(n_371), .Y(n_487) );
AND2x4_ASAP7_75t_L g494 ( .A(n_347), .B(n_354), .Y(n_494) );
AND2x4_ASAP7_75t_L g697 ( .A(n_347), .B(n_358), .Y(n_697) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_352), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x4_ASAP7_75t_L g399 ( .A(n_354), .B(n_395), .Y(n_399) );
BUFx8_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_357), .Y(n_507) );
AND2x4_ASAP7_75t_L g394 ( .A(n_358), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g693 ( .A(n_358), .B(n_395), .Y(n_693) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g445 ( .A(n_361), .Y(n_445) );
INVx1_ASAP7_75t_L g471 ( .A(n_361), .Y(n_471) );
INVx2_ASAP7_75t_L g512 ( .A(n_361), .Y(n_512) );
INVx4_ASAP7_75t_L g535 ( .A(n_361), .Y(n_535) );
INVx4_ASAP7_75t_L g568 ( .A(n_361), .Y(n_568) );
INVx2_ASAP7_75t_L g616 ( .A(n_361), .Y(n_616) );
INVx8_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR2x1_ASAP7_75t_L g363 ( .A(n_364), .B(n_378), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_374), .B2(n_375), .Y(n_364) );
OA21x2_ASAP7_75t_L g472 ( .A1(n_366), .A2(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g454 ( .A(n_368), .Y(n_454) );
BUFx3_ASAP7_75t_L g521 ( .A(n_368), .Y(n_521) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_368), .Y(n_571) );
BUFx8_ASAP7_75t_SL g748 ( .A(n_368), .Y(n_748) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_371), .Y(n_368) );
AND2x4_ASAP7_75t_L g382 ( .A(n_369), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g620 ( .A(n_369), .B(n_383), .Y(n_620) );
AND2x2_ASAP7_75t_L g652 ( .A(n_369), .B(n_371), .Y(n_652) );
AND2x4_ASAP7_75t_L g395 ( .A(n_370), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g407 ( .A(n_371), .B(n_395), .Y(n_407) );
AND2x4_ASAP7_75t_L g491 ( .A(n_371), .B(n_395), .Y(n_491) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_377), .Y(n_522) );
INVx3_ASAP7_75t_L g1009 ( .A(n_377), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B1(n_384), .B2(n_385), .Y(n_378) );
INVx4_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g483 ( .A(n_382), .Y(n_483) );
BUFx3_ASAP7_75t_L g545 ( .A(n_382), .Y(n_545) );
AND2x4_ASAP7_75t_L g404 ( .A(n_383), .B(n_395), .Y(n_404) );
AND2x4_ASAP7_75t_L g490 ( .A(n_383), .B(n_395), .Y(n_490) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g458 ( .A(n_386), .Y(n_458) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g573 ( .A(n_387), .Y(n_573) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_388), .Y(n_519) );
BUFx3_ASAP7_75t_L g543 ( .A(n_388), .Y(n_543) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_400), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx12f_ASAP7_75t_L g444 ( .A(n_393), .Y(n_444) );
BUFx12f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_394), .Y(n_534) );
BUFx3_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_399), .Y(n_439) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_399), .Y(n_505) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_399), .Y(n_540) );
BUFx4f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g509 ( .A(n_403), .Y(n_509) );
INVx1_ASAP7_75t_L g1002 ( .A(n_403), .Y(n_1002) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx12f_ASAP7_75t_L g538 ( .A(n_404), .Y(n_538) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx5_ASAP7_75t_L g447 ( .A(n_407), .Y(n_447) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_407), .Y(n_510) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI21xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g517 ( .A(n_415), .Y(n_517) );
INVx3_ASAP7_75t_L g577 ( .A(n_415), .Y(n_577) );
BUFx4f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx5_ASAP7_75t_L g451 ( .A(n_418), .Y(n_451) );
BUFx2_ASAP7_75t_L g627 ( .A(n_418), .Y(n_627) );
BUFx2_ASAP7_75t_L g1011 ( .A(n_418), .Y(n_1011) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_423), .Y(n_418) );
AND2x2_ASAP7_75t_L g484 ( .A(n_419), .B(n_423), .Y(n_484) );
AND2x4_ASAP7_75t_L g599 ( .A(n_419), .B(n_423), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
INVx1_ASAP7_75t_L g430 ( .A(n_421), .Y(n_430) );
INVx4_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_427), .B(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_427), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g707 ( .A(n_427), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g722 ( .A(n_427), .B(n_723), .Y(n_722) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g549 ( .A(n_428), .Y(n_549) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_429), .Y(n_461) );
INVx1_ASAP7_75t_L g495 ( .A(n_433), .Y(n_495) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
XNOR2x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_462), .Y(n_434) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_437), .B(n_448), .Y(n_436) );
NAND4xp25_ASAP7_75t_SL g437 ( .A(n_438), .B(n_441), .C(n_443), .D(n_446), .Y(n_437) );
NAND4xp25_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .C(n_457), .D(n_459), .Y(n_448) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx4_ASAP7_75t_L g524 ( .A(n_451), .Y(n_524) );
INVx2_ASAP7_75t_L g574 ( .A(n_451), .Y(n_574) );
INVx2_ASAP7_75t_L g746 ( .A(n_451), .Y(n_746) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_SL g739 ( .A(n_460), .Y(n_739) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_461), .Y(n_479) );
INVx1_ASAP7_75t_L g525 ( .A(n_461), .Y(n_525) );
BUFx6f_ASAP7_75t_L g674 ( .A(n_461), .Y(n_674) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g499 ( .A(n_463), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g464 ( .A(n_465), .B(n_472), .C(n_481), .D(n_488), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_466), .B(n_470), .Y(n_465) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx4f_ASAP7_75t_L g614 ( .A(n_468), .Y(n_614) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_477), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g601 ( .A(n_479), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_479), .B(n_622), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_479), .B(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_479), .B(n_1014), .Y(n_1013) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
INVx1_ASAP7_75t_L g645 ( .A(n_486), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_487), .Y(n_647) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_492), .Y(n_488) );
XOR2xp5_ASAP7_75t_L g496 ( .A(n_497), .B(n_555), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_500), .B1(n_553), .B2(n_554), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_499), .Y(n_554) );
INVx1_ASAP7_75t_L g553 ( .A(n_500), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_527), .B1(n_551), .B2(n_552), .Y(n_500) );
INVx1_ASAP7_75t_SL g551 ( .A(n_501), .Y(n_551) );
XOR2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_526), .Y(n_501) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_513), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .C(n_508), .D(n_511), .Y(n_503) );
NAND4xp25_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .C(n_520), .D(n_523), .Y(n_513) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g595 ( .A(n_516), .Y(n_595) );
INVx1_ASAP7_75t_L g736 ( .A(n_516), .Y(n_736) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g705 ( .A(n_517), .Y(n_705) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g552 ( .A(n_528), .Y(n_552) );
XNOR2x1_ASAP7_75t_L g528 ( .A(n_529), .B(n_550), .Y(n_528) );
NAND4xp75_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .C(n_541), .D(n_546), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_549), .B(n_769), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_604), .B1(n_657), .B2(n_658), .Y(n_555) );
INVx1_ASAP7_75t_L g657 ( .A(n_556), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_581), .B1(n_602), .B2(n_603), .Y(n_556) );
INVx1_ASAP7_75t_L g603 ( .A(n_557), .Y(n_603) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND4xp75_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .C(n_569), .D(n_575), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g625 ( .A(n_577), .Y(n_625) );
INVx2_ASAP7_75t_L g669 ( .A(n_577), .Y(n_669) );
INVx2_ASAP7_75t_L g721 ( .A(n_577), .Y(n_721) );
INVx1_ASAP7_75t_L g602 ( .A(n_581), .Y(n_602) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_582), .Y(n_581) );
NAND4xp75_ASAP7_75t_L g583 ( .A(n_584), .B(n_588), .C(n_591), .D(n_594), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_587), .Y(n_584) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .Y(n_596) );
INVx4_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g658 ( .A(n_604), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_628), .B1(n_655), .B2(n_656), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_SL g655 ( .A(n_608), .Y(n_655) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_610), .B(n_618), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .C(n_615), .D(n_617), .Y(n_610) );
NAND4xp25_ASAP7_75t_SL g618 ( .A(n_619), .B(n_623), .C(n_624), .D(n_626), .Y(n_618) );
INVx2_ASAP7_75t_L g642 ( .A(n_620), .Y(n_642) );
INVx2_ASAP7_75t_L g656 ( .A(n_628), .Y(n_656) );
NAND4xp75_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .C(n_639), .D(n_649), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_644), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_643), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B1(n_647), .B2(n_648), .Y(n_644) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
XOR2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_714), .Y(n_660) );
XOR2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_680), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g665 ( .A(n_666), .B(n_675), .Y(n_665) );
NAND4xp25_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .C(n_670), .D(n_671), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND4xp25_ASAP7_75t_SL g675 ( .A(n_676), .B(n_677), .C(n_678), .D(n_679), .Y(n_675) );
OA22x2_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_682), .B1(n_698), .B2(n_713), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OR2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_691), .Y(n_683) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .C(n_687), .D(n_688), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .C(n_695), .D(n_696), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
XOR2xp5_ASAP7_75t_L g713 ( .A(n_699), .B(n_700), .Y(n_713) );
OR2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_708), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .C(n_704), .D(n_706), .Y(n_701) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .C(n_711), .D(n_712), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_716), .B1(n_752), .B2(n_772), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
XNOR2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_732), .Y(n_717) );
INVx1_ASAP7_75t_L g771 ( .A(n_718), .Y(n_771) );
NAND3x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .C(n_727), .Y(n_719) );
AND2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
AND4x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .C(n_730), .D(n_731), .Y(n_727) );
XOR2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NAND4xp75_ASAP7_75t_L g734 ( .A(n_735), .B(n_740), .C(n_744), .D(n_749), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_743), .Y(n_740) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx1_ASAP7_75t_L g766 ( .A(n_748), .Y(n_766) );
AND2x2_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx1_ASAP7_75t_L g772 ( .A(n_752), .Y(n_772) );
XNOR2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_771), .Y(n_752) );
XOR2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_770), .Y(n_753) );
NOR4xp75_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .C(n_761), .D(n_764), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_762), .B(n_763), .Y(n_761) );
OAI21x1_ASAP7_75t_SL g764 ( .A1(n_765), .A2(n_766), .B(n_767), .Y(n_764) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_993), .B1(n_995), .B2(n_1018), .C(n_1023), .Y(n_773) );
AOI211xp5_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_797), .B(n_865), .C(n_959), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_793), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g891 ( .A1(n_776), .A2(n_834), .B1(n_892), .B2(n_894), .C(n_917), .Y(n_891) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_776), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_776), .B(n_836), .Y(n_938) );
AOI221xp5_ASAP7_75t_L g965 ( .A1(n_776), .A2(n_893), .B1(n_901), .B2(n_906), .C(n_966), .Y(n_965) );
AND2x2_ASAP7_75t_L g776 ( .A(n_777), .B(n_789), .Y(n_776) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx3_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
AND2x4_ASAP7_75t_L g790 ( .A(n_781), .B(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g796 ( .A(n_781), .B(n_791), .Y(n_796) );
AND2x2_ASAP7_75t_L g832 ( .A(n_781), .B(n_791), .Y(n_832) );
AND2x4_ASAP7_75t_L g787 ( .A(n_783), .B(n_788), .Y(n_787) );
AND2x4_ASAP7_75t_L g815 ( .A(n_783), .B(n_788), .Y(n_815) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx2_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
AND2x4_ASAP7_75t_L g792 ( .A(n_788), .B(n_791), .Y(n_792) );
AND2x2_ASAP7_75t_L g808 ( .A(n_788), .B(n_791), .Y(n_808) );
AND2x2_ASAP7_75t_L g817 ( .A(n_788), .B(n_791), .Y(n_817) );
BUFx2_ASAP7_75t_L g994 ( .A(n_790), .Y(n_994) );
INVx1_ASAP7_75t_L g890 ( .A(n_793), .Y(n_890) );
INVx4_ASAP7_75t_L g897 ( .A(n_793), .Y(n_897) );
AND2x2_ASAP7_75t_L g901 ( .A(n_793), .B(n_838), .Y(n_901) );
NAND3xp33_ASAP7_75t_L g903 ( .A(n_793), .B(n_853), .C(n_904), .Y(n_903) );
AND2x2_ASAP7_75t_L g906 ( .A(n_793), .B(n_907), .Y(n_906) );
AND2x2_ASAP7_75t_L g958 ( .A(n_793), .B(n_888), .Y(n_958) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_795), .Y(n_793) );
NAND4xp25_ASAP7_75t_L g797 ( .A(n_798), .B(n_833), .C(n_855), .D(n_861), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_810), .Y(n_798) );
HB1xp67_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
HB1xp67_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_801), .B(n_901), .Y(n_943) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g857 ( .A(n_802), .Y(n_857) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_803), .Y(n_878) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g889 ( .A(n_805), .B(n_837), .Y(n_889) );
INVx2_ASAP7_75t_L g907 ( .A(n_805), .Y(n_907) );
INVx4_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
OR2x2_ASAP7_75t_L g863 ( .A(n_806), .B(n_837), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_806), .B(n_875), .Y(n_874) );
OR2x2_ASAP7_75t_L g898 ( .A(n_806), .B(n_838), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g904 ( .A(n_806), .B(n_821), .Y(n_904) );
AND2x2_ASAP7_75t_L g950 ( .A(n_806), .B(n_837), .Y(n_950) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .Y(n_806) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_818), .Y(n_811) );
AND2x2_ASAP7_75t_L g845 ( .A(n_812), .B(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_812), .B(n_853), .Y(n_852) );
AND2x2_ASAP7_75t_L g871 ( .A(n_812), .B(n_821), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_812), .B(n_854), .Y(n_909) );
AND2x2_ASAP7_75t_L g911 ( .A(n_812), .B(n_880), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_812), .B(n_847), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_812), .B(n_941), .Y(n_962) );
AND2x2_ASAP7_75t_L g976 ( .A(n_812), .B(n_825), .Y(n_976) );
CKINVDCx6p67_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g849 ( .A(n_813), .B(n_827), .Y(n_849) );
AND2x2_ASAP7_75t_L g859 ( .A(n_813), .B(n_819), .Y(n_859) );
AND2x2_ASAP7_75t_L g869 ( .A(n_813), .B(n_846), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_813), .B(n_854), .Y(n_885) );
AND2x2_ASAP7_75t_L g893 ( .A(n_813), .B(n_880), .Y(n_893) );
AND2x2_ASAP7_75t_L g900 ( .A(n_813), .B(n_860), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_813), .B(n_825), .Y(n_930) );
AND2x2_ASAP7_75t_L g940 ( .A(n_813), .B(n_941), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_813), .B(n_847), .Y(n_952) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g990 ( .A(n_818), .Y(n_990) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_824), .Y(n_818) );
AND2x2_ASAP7_75t_L g850 ( .A(n_819), .B(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_819), .B(n_949), .Y(n_973) );
INVx3_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_820), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_820), .B(n_845), .Y(n_882) );
AND2x2_ASAP7_75t_L g936 ( .A(n_820), .B(n_937), .Y(n_936) );
AND2x2_ASAP7_75t_L g941 ( .A(n_820), .B(n_860), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_820), .B(n_952), .Y(n_951) );
INVx3_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g875 ( .A(n_821), .Y(n_875) );
INVx2_ASAP7_75t_L g887 ( .A(n_821), .Y(n_887) );
NOR2xp33_ASAP7_75t_L g929 ( .A(n_821), .B(n_930), .Y(n_929) );
NOR2xp33_ASAP7_75t_L g932 ( .A(n_821), .B(n_933), .Y(n_932) );
AND2x2_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g880 ( .A(n_824), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g980 ( .A(n_824), .B(n_875), .Y(n_980) );
OR2x2_ASAP7_75t_L g824 ( .A(n_825), .B(n_827), .Y(n_824) );
AND2x2_ASAP7_75t_L g846 ( .A(n_825), .B(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g854 ( .A(n_825), .Y(n_854) );
AND2x2_ASAP7_75t_L g860 ( .A(n_825), .B(n_827), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_825), .B(n_859), .Y(n_918) );
INVx1_ASAP7_75t_L g847 ( .A(n_827), .Y(n_847) );
AND2x2_ASAP7_75t_L g853 ( .A(n_827), .B(n_854), .Y(n_853) );
OAI21xp33_ASAP7_75t_L g971 ( .A1(n_827), .A2(n_972), .B(n_974), .Y(n_971) );
AND2x2_ASAP7_75t_L g827 ( .A(n_828), .B(n_831), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .B1(n_841), .B2(n_850), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
OAI21xp33_ASAP7_75t_L g881 ( .A1(n_835), .A2(n_882), .B(n_883), .Y(n_881) );
INVx3_ASAP7_75t_SL g835 ( .A(n_836), .Y(n_835) );
AOI21xp33_ASAP7_75t_L g876 ( .A1(n_836), .A2(n_858), .B(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_836), .B(n_897), .Y(n_978) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVxp67_ASAP7_75t_L g914 ( .A(n_837), .Y(n_914) );
AND2x2_ASAP7_75t_L g970 ( .A(n_837), .B(n_897), .Y(n_970) );
INVx2_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g843 ( .A(n_844), .B(n_848), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g872 ( .A(n_845), .B(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g933 ( .A(n_846), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_846), .B(n_859), .Y(n_967) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_849), .B(n_887), .Y(n_916) );
OAI221xp5_ASAP7_75t_L g920 ( .A1(n_850), .A2(n_921), .B1(n_927), .B2(n_934), .C(n_938), .Y(n_920) );
INVx2_ASAP7_75t_L g864 ( .A(n_851), .Y(n_864) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_853), .B(n_896), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_853), .A2(n_859), .B1(n_873), .B2(n_945), .C(n_980), .Y(n_979) );
INVxp67_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_857), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
AND2x2_ASAP7_75t_L g879 ( .A(n_859), .B(n_880), .Y(n_879) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_860), .B(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g945 ( .A(n_860), .Y(n_945) );
OAI21xp5_ASAP7_75t_L g987 ( .A1(n_860), .A2(n_947), .B(n_988), .Y(n_987) );
INVxp67_ASAP7_75t_SL g861 ( .A(n_862), .Y(n_861) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
A2O1A1Ixp33_ASAP7_75t_L g867 ( .A1(n_863), .A2(n_868), .B(n_870), .C(n_872), .Y(n_867) );
AOI211xp5_ASAP7_75t_L g917 ( .A1(n_863), .A2(n_882), .B(n_918), .C(n_919), .Y(n_917) );
INVx1_ASAP7_75t_L g937 ( .A(n_863), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_863), .B(n_964), .Y(n_963) );
NAND4xp25_ASAP7_75t_L g865 ( .A(n_866), .B(n_891), .C(n_920), .D(n_939), .Y(n_865) );
OAI31xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_876), .A3(n_881), .B(n_890), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g956 ( .A(n_870), .Y(n_956) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g892 ( .A(n_875), .B(n_893), .Y(n_892) );
AND2x2_ASAP7_75t_L g975 ( .A(n_875), .B(n_976), .Y(n_975) );
OAI211xp5_ASAP7_75t_SL g921 ( .A1(n_877), .A2(n_922), .B(n_923), .C(n_926), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_878), .B(n_879), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_880), .B(n_936), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
OAI221xp5_ASAP7_75t_L g961 ( .A1(n_885), .A2(n_957), .B1(n_962), .B2(n_963), .C(n_965), .Y(n_961) );
AND2x2_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
OAI21xp33_ASAP7_75t_L g908 ( .A1(n_887), .A2(n_909), .B(n_910), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_887), .B(n_924), .Y(n_923) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_887), .B(n_898), .Y(n_947) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_887), .B(n_925), .Y(n_954) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
OAI221xp5_ASAP7_75t_L g927 ( .A1(n_889), .A2(n_898), .B1(n_919), .B2(n_928), .C(n_931), .Y(n_927) );
O2A1O1Ixp33_ASAP7_75t_SL g959 ( .A1(n_890), .A2(n_960), .B(n_968), .C(n_982), .Y(n_959) );
INVx1_ASAP7_75t_L g981 ( .A(n_892), .Y(n_981) );
NOR2xp33_ASAP7_75t_SL g955 ( .A(n_893), .B(n_956), .Y(n_955) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_895), .B(n_899), .C(n_905), .Y(n_894) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
OR2x2_ASAP7_75t_L g913 ( .A(n_897), .B(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g964 ( .A(n_897), .Y(n_964) );
AND2x2_ASAP7_75t_L g969 ( .A(n_897), .B(n_907), .Y(n_969) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_897), .B(n_919), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g989 ( .A1(n_898), .A2(n_949), .B1(n_990), .B2(n_991), .C(n_992), .Y(n_989) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_900), .A2(n_901), .B(n_902), .Y(n_899) );
INVx1_ASAP7_75t_L g986 ( .A(n_900), .Y(n_986) );
INVxp67_ASAP7_75t_SL g902 ( .A(n_903), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_908), .B1(n_912), .B2(n_915), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_907), .B(n_954), .Y(n_953) );
A2O1A1Ixp33_ASAP7_75t_L g985 ( .A1(n_907), .A2(n_916), .B(n_986), .C(n_987), .Y(n_985) );
INVx1_ASAP7_75t_L g988 ( .A(n_909), .Y(n_988) );
AOI21xp33_ASAP7_75t_L g944 ( .A1(n_910), .A2(n_945), .B(n_946), .Y(n_944) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
NOR2xp33_ASAP7_75t_L g928 ( .A(n_915), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g926 ( .A(n_919), .Y(n_926) );
AOI221xp5_ASAP7_75t_L g939 ( .A1(n_919), .A2(n_940), .B1(n_942), .B2(n_944), .C(n_948), .Y(n_939) );
INVx1_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
OAI322xp33_ASAP7_75t_L g948 ( .A1(n_926), .A2(n_938), .A3(n_949), .B1(n_951), .B2(n_953), .C1(n_955), .C2(n_957), .Y(n_948) );
OAI211xp5_ASAP7_75t_L g977 ( .A1(n_926), .A2(n_978), .B(n_979), .C(n_981), .Y(n_977) );
INVx1_ASAP7_75t_L g991 ( .A(n_929), .Y(n_991) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVxp67_ASAP7_75t_SL g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_950), .B(n_966), .Y(n_992) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVxp67_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
AOI211xp5_ASAP7_75t_SL g982 ( .A1(n_961), .A2(n_983), .B(n_985), .C(n_989), .Y(n_982) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
O2A1O1Ixp33_ASAP7_75t_L g968 ( .A1(n_969), .A2(n_970), .B(n_971), .C(n_977), .Y(n_968) );
INVxp33_ASAP7_75t_SL g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
CKINVDCx5p33_ASAP7_75t_R g993 ( .A(n_994), .Y(n_993) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
HB1xp67_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
OAI22x1_ASAP7_75t_L g997 ( .A1(n_998), .A2(n_1005), .B1(n_1016), .B2(n_1017), .Y(n_997) );
HB1xp67_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_999), .B(n_1006), .Y(n_1016) );
NAND4xp25_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1001), .C(n_1003), .D(n_1004), .Y(n_999) );
NAND4xp25_ASAP7_75t_L g1006 ( .A(n_1007), .B(n_1010), .C(n_1012), .D(n_1015), .Y(n_1006) );
INVx2_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVxp33_ASAP7_75t_SL g1027 ( .A(n_1016), .Y(n_1027) );
INVx1_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1026), .Y(n_1028) );
HB1xp67_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_1034), .Y(n_1033) );
endmodule