module fake_jpeg_1666_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_23),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_17),
.B(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_14),
.B(n_7),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_80),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_78),
.B(n_71),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_94),
.Y(n_117)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_77),
.A2(n_63),
.B1(n_59),
.B2(n_70),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_97),
.B1(n_79),
.B2(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_71),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_63),
.B1(n_59),
.B2(n_70),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_98),
.B1(n_69),
.B2(n_51),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_73),
.B1(n_57),
.B2(n_61),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_74),
.B1(n_58),
.B2(n_69),
.Y(n_98)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_99),
.Y(n_130)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_52),
.C(n_72),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_105),
.C(n_61),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_65),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_111),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_72),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_109),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_88),
.B(n_86),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_108),
.A2(n_51),
.B(n_56),
.Y(n_123)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_62),
.Y(n_111)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_113),
.Y(n_124)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_105),
.B1(n_110),
.B2(n_108),
.Y(n_131)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_119),
.Y(n_145)
);

OAI32xp33_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_98),
.A3(n_52),
.B1(n_53),
.B2(n_67),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_53),
.B1(n_67),
.B2(n_57),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_131),
.B1(n_133),
.B2(n_1),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_2),
.B(n_3),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_125),
.B(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_64),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_134),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_87),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_45),
.C(n_44),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_68),
.B1(n_66),
.B2(n_87),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_0),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_0),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_135),
.B(n_136),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_1),
.Y(n_136)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_56),
.A3(n_54),
.B1(n_83),
.B2(n_4),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_54),
.C(n_2),
.Y(n_141)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_148),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_143),
.B(n_153),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_144),
.B1(n_120),
.B2(n_133),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_121),
.A2(n_50),
.B1(n_49),
.B2(n_47),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_162),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_43),
.C(n_42),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_154),
.C(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_5),
.B(n_6),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_41),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_40),
.C(n_39),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_123),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_138),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_36),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_157),
.B(n_158),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_159),
.A2(n_119),
.B1(n_12),
.B2(n_13),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_160),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_32),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_137),
.A2(n_9),
.B(n_11),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_166),
.B1(n_172),
.B2(n_146),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_145),
.B1(n_151),
.B2(n_152),
.Y(n_166)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_143),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_127),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_170),
.B(n_175),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_31),
.A3(n_29),
.B1(n_16),
.B2(n_17),
.C(n_18),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_147),
.B(n_11),
.C(n_15),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_154),
.C(n_180),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_15),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_180),
.B(n_162),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_157),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_182),
.B(n_185),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_184),
.C(n_188),
.Y(n_195)
);

NOR2xp67_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_161),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_190),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_19),
.B(n_20),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_171),
.A3(n_178),
.B1(n_168),
.B2(n_177),
.C1(n_176),
.C2(n_174),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_164),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_164),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_183),
.C(n_173),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_199),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_179),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_196),
.B1(n_168),
.B2(n_195),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_200),
.A2(n_193),
.B1(n_173),
.B2(n_21),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

AOI322xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_198),
.A3(n_20),
.B1(n_21),
.B2(n_22),
.C1(n_19),
.C2(n_24),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_22),
.C(n_23),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_205),
.B(n_24),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_25),
.Y(n_208)
);


endmodule