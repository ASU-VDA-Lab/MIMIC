module fake_jpeg_11759_n_70 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_13),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_19),
.A2(n_16),
.B1(n_14),
.B2(n_12),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_30),
.A2(n_19),
.B1(n_22),
.B2(n_21),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_34),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_33),
.B1(n_22),
.B2(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_27),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_49),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_0),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_0),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_40),
.C(n_36),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_53),
.C(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_47),
.C(n_21),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_24),
.C(n_26),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_59),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_26),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_60),
.B(n_61),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_63),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_62),
.B1(n_23),
.B2(n_9),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_67),
.A3(n_64),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_66),
.B(n_5),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_70)
);


endmodule