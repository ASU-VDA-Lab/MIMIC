module fake_jpeg_11461_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_50),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_0),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_64),
.Y(n_72)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_66),
.Y(n_75)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_50),
.B1(n_46),
.B2(n_55),
.Y(n_68)
);

AO22x2_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_48),
.B1(n_51),
.B2(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_77),
.B1(n_5),
.B2(n_7),
.Y(n_89)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_54),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_52),
.B1(n_49),
.B2(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_42),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_47),
.B1(n_2),
.B2(n_3),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_79),
.A2(n_63),
.B1(n_57),
.B2(n_3),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_82),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_1),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_84),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_85),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_73),
.B(n_68),
.C(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_94),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_68),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

OR2x6_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_32),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_16),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_18),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_39),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_76),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_101),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_92),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_29),
.B(n_30),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_100),
.C(n_97),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_34),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_107),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_110),
.B(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_112),
.Y(n_123)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_104),
.Y(n_117)
);

AO221x1_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_107),
.C(n_96),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_101),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_107),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_122),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_124),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_118),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_129),
.B(n_123),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_115),
.Y(n_131)
);


endmodule