module fake_jpeg_31530_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_15),
.B1(n_30),
.B2(n_28),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_14),
.B1(n_32),
.B2(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_47),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_39),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_55),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_42),
.B1(n_38),
.B2(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_57),
.B1(n_58),
.B2(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_37),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_1),
.B(n_3),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_68),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_12),
.C(n_21),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_70),
.Y(n_84)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_72),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_11),
.C(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_75),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_4),
.B(n_5),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_17),
.B1(n_7),
.B2(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_4),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_80),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_10),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_64),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_90),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_91),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_84),
.B(n_76),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_82),
.C(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_85),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_98),
.A2(n_99),
.B(n_81),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_100),
.B(n_95),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_97),
.C(n_93),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_92),
.Y(n_104)
);


endmodule