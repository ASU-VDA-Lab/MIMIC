module fake_jpeg_83_n_208 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_208);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_6),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_58),
.Y(n_96)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_70),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVxp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_89),
.Y(n_101)
);

NOR2x1_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_54),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_79),
.A2(n_60),
.B1(n_55),
.B2(n_69),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_76),
.B1(n_55),
.B2(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_97),
.B(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_88),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_104),
.B1(n_109),
.B2(n_61),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_114),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_90),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g107 ( 
.A(n_92),
.B(n_77),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_87),
.B(n_81),
.Y(n_119)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_81),
.B1(n_82),
.B2(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_112),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_0),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_66),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_53),
.B(n_3),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_67),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_63),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_123),
.B(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_72),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_59),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_61),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_29),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_69),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_143),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_104),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_107),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_139),
.B(n_153),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_140),
.A2(n_152),
.B(n_154),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_56),
.B1(n_57),
.B2(n_93),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_57),
.B1(n_53),
.B2(n_23),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_1),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_57),
.B1(n_53),
.B2(n_4),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_150),
.B1(n_156),
.B2(n_132),
.Y(n_173)
);

AOI21x1_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_9),
.B(n_11),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_2),
.B(n_5),
.Y(n_152)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_27),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_7),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

AO22x1_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_31),
.B1(n_50),
.B2(n_49),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_122),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_157),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_7),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_9),
.B(n_11),
.Y(n_175)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_171),
.C(n_172),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_132),
.B1(n_125),
.B2(n_119),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_143),
.B(n_144),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_173),
.A2(n_175),
.B(n_171),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_179),
.B1(n_182),
.B2(n_185),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_138),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_174),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_168),
.A2(n_154),
.B1(n_158),
.B2(n_156),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_133),
.B1(n_153),
.B2(n_14),
.Y(n_182)
);

OAI322xp33_ASAP7_75t_L g184 ( 
.A1(n_169),
.A2(n_34),
.A3(n_44),
.B1(n_43),
.B2(n_42),
.C1(n_41),
.C2(n_40),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_35),
.C(n_51),
.Y(n_191)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_190),
.B1(n_194),
.B2(n_12),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_189),
.A2(n_191),
.B(n_184),
.Y(n_195)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_160),
.B1(n_173),
.B2(n_159),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_192),
.A2(n_193),
.B1(n_176),
.B2(n_164),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_180),
.A2(n_165),
.B1(n_164),
.B2(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_196),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_SL g197 ( 
.A1(n_189),
.A2(n_165),
.B(n_19),
.C(n_22),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_197),
.A2(n_38),
.B(n_36),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_187),
.A2(n_161),
.B1(n_13),
.B2(n_14),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_198),
.A2(n_199),
.B(n_12),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_200),
.A2(n_18),
.B(n_25),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_197),
.B(n_15),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_204),
.B(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_17),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_13),
.C(n_16),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_16),
.Y(n_208)
);


endmodule