module fake_netlist_6_4105_n_297 (n_52, n_16, n_1, n_46, n_18, n_21, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_5, n_77, n_42, n_8, n_24, n_54, n_0, n_32, n_66, n_78, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_27, n_38, n_61, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_41, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_297);

input n_52;
input n_16;
input n_1;
input n_46;
input n_18;
input n_21;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_5;
input n_77;
input n_42;
input n_8;
input n_24;
input n_54;
input n_0;
input n_32;
input n_66;
input n_78;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_27;
input n_38;
input n_61;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_41;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_297;

wire n_91;
wire n_119;
wire n_146;
wire n_163;
wire n_235;
wire n_256;
wire n_193;
wire n_147;
wire n_269;
wire n_258;
wire n_281;
wire n_154;
wire n_191;
wire n_88;
wire n_209;
wire n_98;
wire n_277;
wire n_260;
wire n_265;
wire n_283;
wire n_113;
wire n_223;
wire n_278;
wire n_270;
wire n_279;
wire n_148;
wire n_199;
wire n_138;
wire n_161;
wire n_208;
wire n_226;
wire n_228;
wire n_252;
wire n_266;
wire n_296;
wire n_166;
wire n_184;
wire n_212;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_216;
wire n_83;
wire n_206;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_227;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_204;
wire n_245;
wire n_87;
wire n_195;
wire n_285;
wire n_261;
wire n_189;
wire n_85;
wire n_99;
wire n_130;
wire n_213;
wire n_84;
wire n_257;
wire n_164;
wire n_292;
wire n_100;
wire n_294;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_203;
wire n_254;
wire n_142;
wire n_286;
wire n_143;
wire n_207;
wire n_242;
wire n_180;
wire n_155;
wire n_219;
wire n_291;
wire n_109;
wire n_150;
wire n_233;
wire n_263;
wire n_122;
wire n_264;
wire n_255;
wire n_284;
wire n_205;
wire n_140;
wire n_218;
wire n_120;
wire n_234;
wire n_251;
wire n_214;
wire n_274;
wire n_82;
wire n_236;
wire n_246;
wire n_110;
wire n_151;
wire n_289;
wire n_112;
wire n_172;
wire n_237;
wire n_81;
wire n_244;
wire n_181;
wire n_182;
wire n_124;
wire n_238;
wire n_239;
wire n_126;
wire n_243;
wire n_202;
wire n_94;
wire n_97;
wire n_108;
wire n_267;
wire n_282;
wire n_116;
wire n_280;
wire n_211;
wire n_287;
wire n_220;
wire n_288;
wire n_290;
wire n_117;
wire n_118;
wire n_175;
wire n_224;
wire n_231;
wire n_230;
wire n_93;
wire n_80;
wire n_141;
wire n_240;
wire n_135;
wire n_200;
wire n_196;
wire n_165;
wire n_139;
wire n_134;
wire n_259;
wire n_177;
wire n_176;
wire n_273;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_222;
wire n_95;
wire n_179;
wire n_248;
wire n_107;
wire n_295;
wire n_229;
wire n_253;
wire n_190;
wire n_123;
wire n_262;
wire n_136;
wire n_187;
wire n_89;
wire n_249;
wire n_173;
wire n_201;
wire n_250;
wire n_103;
wire n_111;
wire n_159;
wire n_272;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_183;
wire n_232;
wire n_115;
wire n_128;
wire n_241;
wire n_275;
wire n_194;
wire n_171;
wire n_293;
wire n_192;
wire n_169;
wire n_276;
wire n_221;

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_48),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_43),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_22),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_18),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_73),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_39),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_70),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_0),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_1),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_2),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_90),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_2),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_3),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_4),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_5),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_6),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_8),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_10),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_11),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_12),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_12),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_13),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_14),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

AND2x4_ASAP7_75t_L g138 ( 
.A(n_91),
.B(n_15),
.Y(n_138)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_16),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_118),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_122),
.B1(n_116),
.B2(n_120),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_84),
.B1(n_87),
.B2(n_80),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_140),
.Y(n_148)
);

AO22x2_ASAP7_75t_L g149 ( 
.A1(n_110),
.A2(n_21),
.B1(n_17),
.B2(n_20),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_23),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_113),
.B(n_23),
.Y(n_151)
);

AO22x2_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_117),
.B1(n_134),
.B2(n_131),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_95),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

NAND3x1_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_25),
.C(n_27),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_148),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_125),
.B(n_123),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_130),
.Y(n_160)
);

AND2x4_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

NAND2x1p5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_130),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_134),
.Y(n_167)
);

NAND2x1p5_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_156),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_149),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_135),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_98),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_137),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_133),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_183),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NOR2x1_ASAP7_75t_SL g190 ( 
.A(n_185),
.B(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_142),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_129),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_182),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_132),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_195),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_198),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_188),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_206),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

INVx4_ASAP7_75t_SL g211 ( 
.A(n_206),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_193),
.B1(n_181),
.B2(n_191),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_213),
.A2(n_202),
.B1(n_205),
.B2(n_204),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_201),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_221),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_222),
.A2(n_190),
.B1(n_214),
.B2(n_212),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_218),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_28),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_224),
.A2(n_196),
.B(n_194),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_126),
.B1(n_196),
.B2(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_33),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_34),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_35),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_36),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_40),
.Y(n_238)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_232),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_237),
.B(n_231),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_236),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_47),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_241),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_248),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_243),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_244),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_251),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_254),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_250),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_253),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_257),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_264),
.A2(n_261),
.B1(n_262),
.B2(n_260),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_273),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_79),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_277),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_276),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_281),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_284),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_285),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_289),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_290),
.A2(n_286),
.B1(n_63),
.B2(n_64),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_291),
.A2(n_62),
.B1(n_65),
.B2(n_66),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_292),
.Y(n_295)
);

AOI221xp5_ASAP7_75t_L g296 ( 
.A1(n_295),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.C(n_76),
.Y(n_296)
);

AOI211xp5_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_294),
.B(n_77),
.C(n_78),
.Y(n_297)
);


endmodule