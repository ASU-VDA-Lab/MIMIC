module fake_jpeg_6303_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_22),
.B(n_9),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_42),
.A2(n_49),
.B1(n_33),
.B2(n_25),
.Y(n_55)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_22),
.B(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_33),
.B1(n_36),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_51),
.A2(n_56),
.B1(n_40),
.B2(n_50),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_46),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_63),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_29),
.B1(n_37),
.B2(n_23),
.Y(n_56)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_65),
.Y(n_93)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_45),
.C(n_49),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_95),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_85),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_41),
.B1(n_43),
.B2(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_77),
.A2(n_83),
.B1(n_102),
.B2(n_42),
.Y(n_122)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_41),
.B1(n_43),
.B2(n_49),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_43),
.B1(n_38),
.B2(n_42),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_89),
.Y(n_124)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_39),
.Y(n_95)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_40),
.B1(n_47),
.B2(n_50),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_58),
.B(n_40),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_60),
.B1(n_94),
.B2(n_49),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_101),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_61),
.A2(n_43),
.B1(n_38),
.B2(n_42),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_39),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_35),
.C(n_32),
.Y(n_161)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_107),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_123),
.B1(n_126),
.B2(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_120),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_85),
.B(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_49),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_36),
.C(n_48),
.Y(n_140)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_72),
.B1(n_92),
.B2(n_100),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_38),
.B1(n_45),
.B2(n_66),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_72),
.A2(n_38),
.B1(n_45),
.B2(n_47),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_132),
.Y(n_147)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_95),
.B(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_129),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_76),
.B(n_48),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_141),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_146),
.B1(n_154),
.B2(n_19),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_95),
.B(n_86),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_137),
.A2(n_140),
.B(n_143),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_110),
.A2(n_75),
.B1(n_84),
.B2(n_78),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_144),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_74),
.B1(n_96),
.B2(n_77),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_120),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_83),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_150),
.C(n_152),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_36),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_159),
.B1(n_113),
.B2(n_128),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_114),
.A2(n_20),
.B(n_37),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_114),
.A2(n_20),
.B(n_23),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_157),
.C(n_161),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_48),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_110),
.A2(n_90),
.B1(n_82),
.B2(n_28),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_112),
.A2(n_35),
.B1(n_28),
.B2(n_32),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_17),
.B1(n_19),
.B2(n_119),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_112),
.B1(n_111),
.B2(n_109),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_168),
.B1(n_171),
.B2(n_180),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_173),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_164),
.Y(n_218)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_166),
.A2(n_177),
.B1(n_192),
.B2(n_174),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_105),
.B1(n_125),
.B2(n_103),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_105),
.B1(n_125),
.B2(n_103),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_107),
.B1(n_119),
.B2(n_80),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_175),
.A2(n_182),
.B1(n_135),
.B2(n_141),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_104),
.Y(n_176)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_176),
.Y(n_212)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_127),
.Y(n_179)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_143),
.A2(n_48),
.B1(n_31),
.B2(n_34),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_48),
.B1(n_130),
.B2(n_34),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_186),
.B1(n_189),
.B2(n_148),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_133),
.Y(n_185)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_146),
.A2(n_48),
.B1(n_34),
.B2(n_26),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_139),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_187),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_48),
.B1(n_26),
.B2(n_24),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_191),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_155),
.A2(n_131),
.B1(n_30),
.B2(n_26),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_149),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_220),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_150),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_199),
.C(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_137),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_224),
.B1(n_175),
.B2(n_166),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_190),
.A2(n_153),
.B1(n_152),
.B2(n_138),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_24),
.B1(n_131),
.B2(n_30),
.Y(n_207)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_131),
.C(n_30),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_210),
.C(n_215),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_30),
.C(n_27),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_214),
.B(n_217),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_182),
.B(n_24),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_27),
.B(n_2),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_27),
.B1(n_9),
.B2(n_10),
.Y(n_220)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_222),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_27),
.C(n_2),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_181),
.C(n_162),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_178),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_233),
.B1(n_246),
.B2(n_202),
.Y(n_259)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_218),
.Y(n_230)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_230),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_232),
.B(n_237),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_173),
.B1(n_176),
.B2(n_167),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_210),
.B(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_200),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_224),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_239),
.Y(n_265)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_245),
.Y(n_251)
);

XNOR2x1_ASAP7_75t_SL g241 ( 
.A(n_195),
.B(n_180),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_241),
.B(n_242),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_186),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_191),
.B1(n_171),
.B2(n_169),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_199),
.B(n_189),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_1),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_209),
.C(n_203),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_254),
.C(n_255),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_241),
.A2(n_194),
.B(n_213),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_244),
.B1(n_227),
.B2(n_243),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_216),
.C(n_208),
.Y(n_254)
);

AOI211xp5_ASAP7_75t_SL g256 ( 
.A1(n_249),
.A2(n_215),
.B(n_217),
.C(n_204),
.Y(n_256)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_184),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_267),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_248),
.B(n_235),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_206),
.C(n_220),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_266),
.C(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_214),
.C(n_217),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_231),
.B(n_219),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_1),
.C(n_3),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_11),
.C(n_15),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_268),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_226),
.B1(n_227),
.B2(n_243),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_274),
.A2(n_284),
.B1(n_286),
.B2(n_290),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_264),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_275),
.B(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_237),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_281),
.B(n_282),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_229),
.Y(n_280)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_229),
.B(n_236),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_238),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_265),
.A2(n_254),
.B(n_261),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_256),
.A2(n_239),
.B1(n_236),
.B2(n_5),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_253),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_289),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_271),
.C(n_263),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_270),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_252),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_296),
.C(n_304),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_270),
.Y(n_296)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_276),
.B(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_267),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_12),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_12),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_306),
.C(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_7),
.C(n_8),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_286),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_310),
.A2(n_313),
.B(n_318),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_287),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_274),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_288),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_278),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_283),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_297),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_294),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_325),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_291),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_299),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_328),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_293),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_327),
.A2(n_307),
.B(n_296),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_308),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_324),
.A2(n_318),
.B(n_311),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_331),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_328),
.A2(n_12),
.B(n_13),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_335),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_323),
.B(n_16),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_330),
.B(n_321),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_337),
.B(n_338),
.C(n_16),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_327),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_336),
.B(n_332),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_341),
.C(n_339),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_16),
.B(n_7),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_343),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_7),
.B1(n_8),
.B2(n_333),
.Y(n_345)
);

AO21x1_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_7),
.B(n_8),
.Y(n_346)
);


endmodule