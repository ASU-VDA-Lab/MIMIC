module real_jpeg_17968_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_382),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_0),
.B(n_383),
.Y(n_382)
);

NAND2x1p5_ASAP7_75t_L g34 ( 
.A(n_1),
.B(n_35),
.Y(n_34)
);

AND2x4_ASAP7_75t_SL g39 ( 
.A(n_1),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_1),
.B(n_65),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g98 ( 
.A(n_1),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_128),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_2),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_3),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_3),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_4),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_4),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_4),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_4),
.B(n_304),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_4),
.B(n_320),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_6),
.B(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_6),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_6),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_6),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_6),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_6),
.B(n_35),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_7),
.Y(n_184)
);

INVxp33_ASAP7_75t_L g383 ( 
.A(n_8),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_9),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_9),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_9),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_9),
.Y(n_241)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g204 ( 
.A(n_12),
.Y(n_204)
);

BUFx4f_ASAP7_75t_L g306 ( 
.A(n_12),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g132 ( 
.A(n_13),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_162),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_161),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_19),
.B(n_136),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_90),
.C(n_105),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_20),
.B(n_90),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_22),
.B(n_37),
.C(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

AO22x1_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_26),
.B1(n_70),
.B2(n_71),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_25),
.A2(n_26),
.B1(n_63),
.B2(n_64),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_67),
.C(n_70),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_26),
.B(n_28),
.C(n_34),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_26),
.A2(n_64),
.B(n_181),
.C(n_219),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_27),
.Y(n_177)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.C(n_51),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_34),
.A2(n_36),
.B1(n_51),
.B2(n_133),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_34),
.A2(n_36),
.B1(n_97),
.B2(n_103),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_34),
.B(n_64),
.C(n_98),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_38),
.B(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.C(n_46),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_39),
.A2(n_42),
.B(n_109),
.Y(n_108)
);

NAND2x1p5_ASAP7_75t_L g109 ( 
.A(n_39),
.B(n_42),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_39),
.B(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_39),
.A2(n_113),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_39),
.A2(n_201),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_39),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_39),
.A2(n_113),
.B1(n_211),
.B2(n_217),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR2x1_ASAP7_75t_R g187 ( 
.A(n_41),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_41),
.A2(n_42),
.B1(n_205),
.B2(n_206),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_42),
.B(n_57),
.C(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_46),
.A2(n_76),
.B1(n_108),
.B2(n_110),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_46),
.A2(n_76),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_46),
.B(n_109),
.C(n_240),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_50),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_51),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_51),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_51),
.B(n_80),
.C(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_51),
.B(n_318),
.C(n_319),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_51),
.B(n_130),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_51),
.A2(n_133),
.B1(n_319),
.B2(n_340),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_66),
.C(n_75),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_55),
.B(n_347),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_56),
.A2(n_57),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_57),
.A2(n_273),
.B(n_279),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_57),
.B(n_273),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_69),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_58),
.B(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_60),
.Y(n_243)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_63),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_63),
.B(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_63),
.B(n_226),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_66),
.B(n_75),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_67),
.A2(n_68),
.B1(n_127),
.B2(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_67),
.A2(n_68),
.B1(n_240),
.B2(n_244),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_67),
.B(n_244),
.C(n_290),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_68),
.B(n_155),
.C(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_80),
.C(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_79),
.A2(n_80),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_79),
.B(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_123),
.C(n_127),
.Y(n_122)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_92),
.B(n_95),
.C(n_96),
.Y(n_160)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_98),
.A2(n_127),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_101),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g215 ( 
.A1(n_98),
.A2(n_193),
.B(n_216),
.C(n_219),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_98),
.B(n_193),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_98),
.A2(n_154),
.B1(n_193),
.B2(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_98),
.A2(n_154),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_104),
.B(n_154),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_104),
.B(n_127),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_105),
.B(n_379),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_120),
.C(n_134),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_106),
.B(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_118),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_107),
.B(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_108),
.A2(n_110),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_109),
.B(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_110),
.A2(n_187),
.B(n_193),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_111),
.B(n_118),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_112),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_113),
.A2(n_188),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_113),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_113),
.A2(n_123),
.B1(n_217),
.B2(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_113),
.B(n_123),
.C(n_253),
.Y(n_309)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_153),
.Y(n_152)
);

XNOR2x1_ASAP7_75t_L g328 ( 
.A(n_117),
.B(n_329),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_120),
.B(n_134),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_130),
.C(n_133),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_121),
.A2(n_122),
.B1(n_322),
.B2(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_123),
.A2(n_127),
.B1(n_155),
.B2(n_267),
.Y(n_332)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_127),
.A2(n_157),
.B(n_158),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_130),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_131),
.B(n_206),
.C(n_303),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_160),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_150),
.B1(n_151),
.B2(n_159),
.Y(n_140)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_141),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_156),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_375),
.B(n_380),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_312),
.A3(n_362),
.B1(n_368),
.B2(n_373),
.C(n_374),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_283),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_257),
.B(n_282),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_234),
.B(n_256),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_213),
.B(n_233),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_196),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_170),
.B(n_196),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_178),
.B2(n_179),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_172),
.B(n_179),
.C(n_185),
.Y(n_235)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_176),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_176),
.A2(n_253),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_181),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_180),
.A2(n_181),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_225),
.B(n_227),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.C(n_209),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_209),
.B1(n_210),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_200),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_200),
.A2(n_201),
.B(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_205),
.A2(n_206),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_223),
.B(n_232),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_220),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_229),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_228),
.B(n_231),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_236),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_246),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_245),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_245),
.C(n_246),
.Y(n_281)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_250),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_251),
.C(n_255),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_281),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_281),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_269),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_261),
.C(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_265),
.C(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_280),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_272),
.C(n_280),
.Y(n_311)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_279),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_284),
.B(n_285),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_298),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_286),
.B(n_299),
.C(n_311),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_292),
.B2(n_293),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_289),
.B(n_292),
.C(n_296),
.Y(n_358)
);

XNOR2x2_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_311),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_307),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_309),
.C(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_350),
.Y(n_312)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_343),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_314),
.B(n_343),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_333),
.C(n_341),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_341),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_326),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_316)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_325),
.C(n_326),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.C(n_331),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_327),
.A2(n_328),
.B1(n_330),
.B2(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

XOR2x2_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.C(n_337),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_337),
.B1(n_338),
.B2(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_336),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_348),
.C(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

AOI31xp67_ASAP7_75t_SL g368 ( 
.A1(n_350),
.A2(n_363),
.A3(n_369),
.B(n_372),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_353),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_358),
.C(n_359),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_354),
.A2(n_355),
.B1(n_359),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_355),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_358),
.B(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_359),
.Y(n_366)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_367),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_371),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_378),
.Y(n_381)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);


endmodule