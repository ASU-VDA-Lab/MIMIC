module real_jpeg_14391_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_202;
wire n_128;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_1),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_58),
.B1(n_61),
.B2(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_69),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_34),
.B1(n_40),
.B2(n_69),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_4),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_63),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_4),
.B(n_189),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_61),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g251 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_178),
.Y(n_251)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_4),
.A2(n_46),
.B(n_49),
.C(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_4),
.B(n_85),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_4),
.B(n_37),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_4),
.B(n_54),
.Y(n_278)
);

AOI21xp33_ASAP7_75t_L g287 ( 
.A1(n_4),
.A2(n_61),
.B(n_237),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_5),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_5),
.A2(n_53),
.B1(n_58),
.B2(n_61),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_5),
.A2(n_34),
.B1(n_40),
.B2(n_53),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_5),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_320)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_7),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_7),
.A2(n_39),
.B1(n_58),
.B2(n_61),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_7),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_8),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_8),
.A2(n_58),
.B1(n_61),
.B2(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_159),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_8),
.A2(n_34),
.B1(n_40),
.B2(n_159),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_9),
.A2(n_44),
.B1(n_58),
.B2(n_61),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_9),
.A2(n_44),
.B1(n_63),
.B2(n_64),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_9),
.A2(n_34),
.B1(n_40),
.B2(n_44),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_11),
.Y(n_339)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_12),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_13),
.A2(n_58),
.B1(n_61),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_13),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_77),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_34),
.B1(n_40),
.B2(n_77),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_16),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_16),
.A2(n_58),
.B1(n_61),
.B2(n_67),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_16),
.A2(n_45),
.B1(n_46),
.B2(n_67),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_16),
.A2(n_34),
.B1(n_40),
.B2(n_67),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_17),
.A2(n_63),
.B1(n_64),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_17),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_17),
.A2(n_58),
.B1(n_61),
.B2(n_123),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_17),
.A2(n_45),
.B1(n_46),
.B2(n_123),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_17),
.A2(n_34),
.B1(n_40),
.B2(n_123),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_21),
.B(n_338),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_18),
.B(n_339),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_19),
.A2(n_63),
.B1(n_64),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_19),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_19),
.A2(n_58),
.B1(n_61),
.B2(n_186),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_19),
.A2(n_45),
.B1(n_46),
.B2(n_186),
.Y(n_252)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_19),
.A2(n_34),
.B1(n_40),
.B2(n_186),
.Y(n_273)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_333),
.B(n_336),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_325),
.B(n_329),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_312),
.B(n_324),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_137),
.B(n_309),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_124),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_100),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_27),
.B(n_100),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_70),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_28),
.B(n_86),
.C(n_98),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_55),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_29),
.A2(n_30),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_41),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_31),
.A2(n_32),
.B1(n_55),
.B2(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_31),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_37),
.B(n_38),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_33),
.A2(n_37),
.B1(n_38),
.B2(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_33),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_33),
.A2(n_37),
.B1(n_150),
.B2(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_33),
.A2(n_37),
.B1(n_174),
.B2(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_33),
.A2(n_37),
.B1(n_216),
.B2(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_33),
.A2(n_37),
.B1(n_240),
.B2(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_33),
.A2(n_37),
.B1(n_178),
.B2(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_33),
.A2(n_37),
.B1(n_266),
.B2(n_273),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_34),
.B(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_36),
.A2(n_114),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_36),
.A2(n_148),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_40),
.A2(n_50),
.B(n_178),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_52),
.B2(n_54),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_43),
.A2(n_47),
.B1(n_54),
.B2(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_46),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_45),
.A2(n_61),
.A3(n_82),
.B1(n_236),
.B2(n_238),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_46),
.B(n_81),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_52),
.B1(n_54),
.B2(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_47),
.A2(n_54),
.B(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_47),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_47),
.A2(n_54),
.B1(n_153),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_47),
.A2(n_54),
.B1(n_204),
.B2(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_47),
.A2(n_54),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_47),
.A2(n_54),
.B1(n_252),
.B2(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_51),
.A2(n_118),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_51),
.A2(n_154),
.B1(n_231),
.B2(n_289),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_55),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_57),
.B1(n_68),
.B2(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_56),
.A2(n_57),
.B1(n_89),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_56),
.A2(n_57),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_56),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_56),
.A2(n_57),
.B1(n_185),
.B2(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_57),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_57)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_61),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_58),
.A2(n_60),
.A3(n_63),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_59),
.B(n_61),
.Y(n_176)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_64),
.B(n_178),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_86),
.B1(n_98),
.B2(n_99),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_71),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_71),
.A2(n_72),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_84),
.B1(n_85),
.B2(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_78),
.A2(n_85),
.B1(n_180),
.B2(n_182),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_78),
.A2(n_85),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_78),
.A2(n_85),
.B(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_79),
.A2(n_80),
.B1(n_96),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_79),
.A2(n_80),
.B1(n_120),
.B2(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_79),
.A2(n_80),
.B1(n_181),
.B2(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_79),
.A2(n_80),
.B1(n_212),
.B2(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_80),
.Y(n_85)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_87),
.A2(n_88),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_92),
.C(n_94),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_88),
.B(n_127),
.C(n_130),
.Y(n_313)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_97),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_97),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_92),
.B(n_133),
.C(n_135),
.Y(n_323)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_106),
.C(n_108),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_101),
.A2(n_102),
.B1(n_106),
.B2(n_107),
.Y(n_161)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_108),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_119),
.C(n_121),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_110),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_121),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_124),
.A2(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_125),
.B(n_126),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_134),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_136),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_162),
.B(n_308),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_160),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_139),
.B(n_160),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_144),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.C(n_157),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_146),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_147),
.B(n_151),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_157),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_192),
.B(n_307),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_190),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_164),
.B(n_190),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_169),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_170),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_179),
.C(n_183),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_183),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_187),
.A2(n_189),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_187),
.A2(n_189),
.B1(n_320),
.B2(n_327),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_187),
.A2(n_189),
.B(n_327),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_223),
.B(n_301),
.C(n_306),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_217),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_194),
.B(n_217),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_207),
.C(n_209),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_195),
.A2(n_196),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_201),
.C(n_206),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_209),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.C(n_215),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_210),
.B(n_228),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_215),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_300),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_244),
.B(n_299),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_241),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_226),
.B(n_241),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_229),
.A2(n_232),
.B1(n_233),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_229),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_234),
.A2(n_235),
.B1(n_239),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_242),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_293),
.B(n_298),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_282),
.B(n_292),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_262),
.B(n_281),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_255),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_248),
.B(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_260),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_258),
.C(n_260),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_270),
.B(n_280),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_268),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_279),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_283),
.B(n_284),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_290),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_288),
.C(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_294),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_313),
.B(n_314),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_318),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_316),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_321),
.C(n_323),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_328),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_326),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_334),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_328),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_335),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_335),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_337),
.Y(n_336)
);


endmodule