module fake_jpeg_5963_n_230 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_230);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_16),
.B(n_7),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_6),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_55),
.Y(n_74)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_19),
.B1(n_23),
.B2(n_16),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_32),
.A2(n_29),
.B1(n_21),
.B2(n_23),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_21),
.B1(n_14),
.B2(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_31),
.B(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_15),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_24),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_57),
.A2(n_20),
.B1(n_15),
.B2(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_14),
.Y(n_58)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_27),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_62),
.B1(n_70),
.B2(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_32),
.B1(n_40),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_30),
.B1(n_40),
.B2(n_21),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_50),
.A2(n_30),
.B1(n_35),
.B2(n_37),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_73),
.B1(n_39),
.B2(n_20),
.Y(n_98)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_35),
.B1(n_39),
.B2(n_21),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_42),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_28),
.B1(n_22),
.B2(n_16),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_70),
.B1(n_55),
.B2(n_58),
.Y(n_94)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_72),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_88),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_47),
.C(n_41),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_85),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_47),
.C(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_18),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_57),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_99),
.B(n_28),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_54),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_74),
.C(n_51),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_103),
.C(n_59),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_100),
.B1(n_102),
.B2(n_19),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_36),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_96),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_36),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_66),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_98),
.A2(n_19),
.B1(n_22),
.B2(n_66),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_27),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_46),
.B1(n_43),
.B2(n_56),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_35),
.B1(n_59),
.B2(n_28),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_18),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_36),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_110),
.B1(n_112),
.B2(n_90),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_120),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_116),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_117),
.B(n_118),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_98),
.B1(n_85),
.B2(n_84),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_95),
.B(n_101),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_38),
.B1(n_36),
.B2(n_71),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_83),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_97),
.A2(n_79),
.B1(n_81),
.B2(n_71),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_119),
.B1(n_123),
.B2(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_103),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_26),
.B(n_24),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_87),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_122),
.B(n_99),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_83),
.A2(n_59),
.B1(n_26),
.B2(n_49),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_86),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_110),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_135),
.A2(n_111),
.B(n_108),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_104),
.C(n_102),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_143),
.C(n_131),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_139),
.B(n_141),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_112),
.B1(n_122),
.B2(n_118),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_93),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_119),
.B1(n_112),
.B2(n_109),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_105),
.B(n_90),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_145),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_140),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_158),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_121),
.C(n_117),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_127),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_155),
.A2(n_132),
.B1(n_130),
.B2(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_161),
.C(n_128),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_160),
.B(n_113),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_116),
.C(n_117),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_129),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_133),
.C(n_131),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_164),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_174),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_160),
.A2(n_155),
.B1(n_147),
.B2(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_148),
.B1(n_26),
.B2(n_49),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_173),
.C(n_178),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_139),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_148),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_175),
.B1(n_151),
.B2(n_149),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_138),
.C(n_140),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_36),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_159),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_182),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_186),
.Y(n_196)
);

OAI322xp33_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_153),
.A3(n_161),
.B1(n_147),
.B2(n_163),
.C1(n_149),
.C2(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_189),
.B1(n_17),
.B2(n_49),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_158),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_191),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_38),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_0),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_167),
.B1(n_170),
.B2(n_169),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_198),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_171),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_199),
.C(n_184),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_167),
.B(n_178),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_6),
.B(n_13),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_184),
.B(n_9),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_9),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_199),
.C(n_194),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_188),
.C(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.Y(n_211)
);

OAI221xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_180),
.B1(n_38),
.B2(n_17),
.C(n_4),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_210),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_5),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_1),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_216),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_215),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_209),
.A2(n_10),
.B(n_13),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_5),
.C(n_12),
.Y(n_216)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_1),
.B(n_2),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_211),
.A2(n_4),
.B1(n_10),
.B2(n_11),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_222),
.C(n_2),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_38),
.B(n_10),
.Y(n_220)
);

NOR4xp25_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_212),
.C(n_2),
.D(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_224),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_219),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_226),
.C(n_3),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_3),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_228),
.Y(n_230)
);


endmodule