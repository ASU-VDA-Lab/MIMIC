module real_aes_7933_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_404;
wire n_288;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_314;
wire n_252;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_0), .B(n_84), .C(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g446 ( .A(n_0), .Y(n_446) );
INVx1_ASAP7_75t_L g478 ( .A(n_1), .Y(n_478) );
INVx1_ASAP7_75t_L g190 ( .A(n_2), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_3), .A2(n_38), .B1(n_151), .B2(n_508), .Y(n_523) );
AOI21xp33_ASAP7_75t_L g158 ( .A1(n_4), .A2(n_132), .B(n_159), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_5), .B(n_125), .Y(n_491) );
AND2x6_ASAP7_75t_L g137 ( .A(n_6), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_8), .B(n_103), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_8), .B(n_39), .Y(n_447) );
INVx1_ASAP7_75t_L g165 ( .A(n_9), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_10), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g130 ( .A(n_11), .Y(n_130) );
INVx1_ASAP7_75t_L g472 ( .A(n_12), .Y(n_472) );
INVx1_ASAP7_75t_L g246 ( .A(n_13), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_14), .B(n_173), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_15), .B(n_126), .Y(n_549) );
AO32x2_ASAP7_75t_L g521 ( .A1(n_16), .A2(n_125), .A3(n_170), .B1(n_500), .B2(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_17), .A2(n_115), .B1(n_116), .B2(n_441), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_17), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_18), .B(n_151), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_19), .B(n_146), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_20), .B(n_126), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_21), .A2(n_50), .B1(n_151), .B2(n_508), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_22), .B(n_132), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_23), .A2(n_75), .B1(n_151), .B2(n_173), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_24), .B(n_151), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_25), .B(n_154), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_26), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_27), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_28), .A2(n_100), .B1(n_108), .B2(n_764), .Y(n_99) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_29), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_30), .B(n_167), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_31), .B(n_163), .Y(n_192) );
INVx1_ASAP7_75t_L g179 ( .A(n_32), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_33), .B(n_167), .Y(n_538) );
INVx2_ASAP7_75t_L g135 ( .A(n_34), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_35), .B(n_151), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_36), .B(n_167), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_37), .A2(n_137), .B(n_141), .C(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g103 ( .A(n_39), .Y(n_103) );
INVx1_ASAP7_75t_L g177 ( .A(n_40), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_41), .B(n_163), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_42), .B(n_151), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_43), .A2(n_85), .B1(n_209), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_44), .B(n_151), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_45), .B(n_151), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_46), .Y(n_180) );
OAI222xp33_ASAP7_75t_L g452 ( .A1(n_47), .A2(n_453), .B1(n_751), .B2(n_752), .C1(n_757), .C2(n_761), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g751 ( .A(n_47), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_48), .B(n_477), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_49), .B(n_132), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_51), .A2(n_60), .B1(n_151), .B2(n_173), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_52), .A2(n_141), .B1(n_173), .B2(n_175), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_53), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_54), .B(n_151), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g187 ( .A(n_55), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_56), .B(n_151), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_57), .A2(n_150), .B(n_162), .C(n_164), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g222 ( .A(n_58), .Y(n_222) );
INVx1_ASAP7_75t_L g160 ( .A(n_59), .Y(n_160) );
INVx1_ASAP7_75t_L g138 ( .A(n_61), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_62), .B(n_151), .Y(n_479) );
INVx1_ASAP7_75t_L g129 ( .A(n_63), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_64), .Y(n_112) );
AO32x2_ASAP7_75t_L g505 ( .A1(n_65), .A2(n_125), .A3(n_226), .B1(n_500), .B2(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g498 ( .A(n_66), .Y(n_498) );
INVx1_ASAP7_75t_L g533 ( .A(n_67), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_68), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_SL g145 ( .A1(n_69), .A2(n_146), .B(n_147), .C(n_150), .Y(n_145) );
INVxp67_ASAP7_75t_L g148 ( .A(n_70), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_71), .B(n_173), .Y(n_534) );
INVx1_ASAP7_75t_L g107 ( .A(n_72), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_73), .Y(n_183) );
INVx1_ASAP7_75t_L g215 ( .A(n_74), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_76), .A2(n_137), .B(n_141), .C(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_77), .B(n_508), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_78), .B(n_173), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_79), .B(n_191), .Y(n_205) );
INVx2_ASAP7_75t_L g127 ( .A(n_80), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_81), .B(n_146), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_82), .B(n_173), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_83), .A2(n_137), .B(n_141), .C(n_189), .Y(n_188) );
OR2x2_ASAP7_75t_L g443 ( .A(n_84), .B(n_444), .Y(n_443) );
OR2x2_ASAP7_75t_L g455 ( .A(n_84), .B(n_445), .Y(n_455) );
INVx2_ASAP7_75t_L g459 ( .A(n_84), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_86), .A2(n_98), .B1(n_173), .B2(n_174), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_87), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_88), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_89), .A2(n_137), .B(n_141), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_90), .Y(n_236) );
INVx1_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_92), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_93), .B(n_191), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_94), .B(n_173), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_95), .B(n_125), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_97), .A2(n_132), .B(n_139), .Y(n_131) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
BUFx4f_ASAP7_75t_SL g764 ( .A(n_101), .Y(n_764) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_104), .Y(n_101) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_113), .B(n_451), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_SL g763 ( .A(n_111), .Y(n_763) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_442), .B(n_448), .Y(n_113) );
INVx2_ASAP7_75t_L g441 ( .A(n_116), .Y(n_441) );
INVx1_ASAP7_75t_SL g456 ( .A(n_116), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_116), .A2(n_753), .B1(n_755), .B2(n_756), .Y(n_752) );
INVx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND4x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_359), .C(n_406), .D(n_426), .Y(n_117) );
NOR3xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_289), .C(n_314), .Y(n_118) );
OAI211xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_197), .B(n_249), .C(n_279), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_168), .Y(n_121) );
INVx3_ASAP7_75t_SL g331 ( .A(n_122), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_122), .B(n_262), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_122), .B(n_184), .Y(n_412) );
AND2x2_ASAP7_75t_L g435 ( .A(n_122), .B(n_301), .Y(n_435) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_156), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g253 ( .A(n_124), .B(n_157), .Y(n_253) );
INVx3_ASAP7_75t_L g266 ( .A(n_124), .Y(n_266) );
AND2x2_ASAP7_75t_L g271 ( .A(n_124), .B(n_156), .Y(n_271) );
OR2x2_ASAP7_75t_L g322 ( .A(n_124), .B(n_263), .Y(n_322) );
BUFx2_ASAP7_75t_L g342 ( .A(n_124), .Y(n_342) );
AND2x2_ASAP7_75t_L g352 ( .A(n_124), .B(n_263), .Y(n_352) );
AND2x2_ASAP7_75t_L g358 ( .A(n_124), .B(n_169), .Y(n_358) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_131), .B(n_153), .Y(n_124) );
INVx4_ASAP7_75t_L g155 ( .A(n_125), .Y(n_155) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_125), .A2(n_484), .B(n_491), .Y(n_483) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_127), .B(n_128), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx2_ASAP7_75t_L g240 ( .A(n_132), .Y(n_240) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_133), .B(n_137), .Y(n_181) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g477 ( .A(n_134), .Y(n_477) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
INVx1_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
INVx1_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx1_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
INVx3_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_136), .Y(n_163) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx4_ASAP7_75t_SL g152 ( .A(n_137), .Y(n_152) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_137), .A2(n_471), .B(n_475), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_137), .A2(n_485), .B(n_488), .Y(n_484) );
BUFx3_ASAP7_75t_L g500 ( .A(n_137), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_137), .A2(n_513), .B(n_517), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_137), .A2(n_532), .B(n_535), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_144), .B(n_145), .C(n_152), .Y(n_139) );
O2A1O1Ixp33_ASAP7_75t_L g159 ( .A1(n_140), .A2(n_152), .B(n_160), .C(n_161), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_140), .A2(n_152), .B(n_242), .C(n_243), .Y(n_241) );
INVx5_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_142), .Y(n_151) );
BUFx3_ASAP7_75t_L g209 ( .A(n_142), .Y(n_209) );
INVx1_ASAP7_75t_L g508 ( .A(n_142), .Y(n_508) );
INVx1_ASAP7_75t_L g516 ( .A(n_146), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_149), .B(n_165), .Y(n_164) );
INVx5_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g506 ( .A1(n_149), .A2(n_163), .B1(n_507), .B2(n_509), .Y(n_506) );
O2A1O1Ixp5_ASAP7_75t_SL g532 ( .A1(n_150), .A2(n_191), .B(n_533), .C(n_534), .Y(n_532) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_151), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g171 ( .A1(n_152), .A2(n_172), .B1(n_180), .B2(n_181), .Y(n_171) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_154), .A2(n_158), .B(n_166), .Y(n_157) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_SL g211 ( .A(n_155), .B(n_212), .Y(n_211) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_155), .A2(n_545), .B(n_548), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g563 ( .A(n_155), .B(n_500), .C(n_545), .Y(n_563) );
INVx1_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_157), .B(n_263), .Y(n_277) );
INVx2_ASAP7_75t_L g287 ( .A(n_157), .Y(n_287) );
AND2x2_ASAP7_75t_L g300 ( .A(n_157), .B(n_266), .Y(n_300) );
OR2x2_ASAP7_75t_L g311 ( .A(n_157), .B(n_263), .Y(n_311) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_157), .B(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g369 ( .A(n_157), .Y(n_369) );
AND2x2_ASAP7_75t_L g415 ( .A(n_157), .B(n_169), .Y(n_415) );
O2A1O1Ixp5_ASAP7_75t_L g497 ( .A1(n_162), .A2(n_476), .B(n_498), .C(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_162), .A2(n_518), .B(n_519), .Y(n_517) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx4_ASAP7_75t_L g232 ( .A(n_163), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_163), .A2(n_480), .B1(n_523), .B2(n_524), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_163), .A2(n_480), .B1(n_546), .B2(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
INVx2_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_167), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_167), .A2(n_512), .B(n_520), .Y(n_511) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_167), .A2(n_531), .B(n_538), .Y(n_530) );
INVx3_ASAP7_75t_SL g288 ( .A(n_168), .Y(n_288) );
OR2x2_ASAP7_75t_L g341 ( .A(n_168), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_184), .Y(n_168) );
INVx3_ASAP7_75t_L g263 ( .A(n_169), .Y(n_263) );
AND2x2_ASAP7_75t_L g330 ( .A(n_169), .B(n_185), .Y(n_330) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_169), .Y(n_398) );
AOI33xp33_ASAP7_75t_L g402 ( .A1(n_169), .A2(n_331), .A3(n_338), .B1(n_347), .B2(n_403), .B3(n_404), .Y(n_402) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_182), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_170), .B(n_183), .Y(n_182) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_170), .A2(n_186), .B(n_194), .Y(n_185) );
INVx2_ASAP7_75t_L g210 ( .A(n_170), .Y(n_210) );
INVx2_ASAP7_75t_L g193 ( .A(n_173), .Y(n_193) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_176), .A2(n_177), .B1(n_178), .B2(n_179), .Y(n_175) );
INVx2_ASAP7_75t_L g178 ( .A(n_176), .Y(n_178) );
INVx4_ASAP7_75t_L g244 ( .A(n_176), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_181), .A2(n_187), .B(n_188), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g214 ( .A1(n_181), .A2(n_215), .B(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g251 ( .A(n_184), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_184), .B(n_266), .Y(n_265) );
NOR3xp33_ASAP7_75t_L g325 ( .A(n_184), .B(n_326), .C(n_328), .Y(n_325) );
AND2x2_ASAP7_75t_L g351 ( .A(n_184), .B(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_184), .B(n_358), .Y(n_361) );
AND2x2_ASAP7_75t_L g414 ( .A(n_184), .B(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx3_ASAP7_75t_L g270 ( .A(n_185), .Y(n_270) );
OR2x2_ASAP7_75t_L g364 ( .A(n_185), .B(n_263), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_192), .C(n_193), .Y(n_189) );
INVx2_ASAP7_75t_L g480 ( .A(n_191), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_191), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_191), .A2(n_495), .B(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_193), .A2(n_472), .B(n_473), .C(n_474), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_196), .B(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_196), .B(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_223), .Y(n_197) );
AOI32xp33_ASAP7_75t_L g315 ( .A1(n_198), .A2(n_316), .A3(n_318), .B1(n_320), .B2(n_323), .Y(n_315) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_198), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g418 ( .A(n_198), .Y(n_418) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g350 ( .A(n_199), .B(n_334), .Y(n_350) );
AND2x2_ASAP7_75t_L g370 ( .A(n_199), .B(n_296), .Y(n_370) );
AND2x2_ASAP7_75t_L g438 ( .A(n_199), .B(n_356), .Y(n_438) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
INVx3_ASAP7_75t_L g259 ( .A(n_200), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_200), .B(n_257), .Y(n_273) );
OR2x2_ASAP7_75t_L g278 ( .A(n_200), .B(n_256), .Y(n_278) );
INVx1_ASAP7_75t_L g285 ( .A(n_200), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_200), .B(n_267), .Y(n_293) );
AND2x2_ASAP7_75t_L g295 ( .A(n_200), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_200), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g348 ( .A(n_200), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_200), .B(n_433), .Y(n_432) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_211), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_210), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_207), .A2(n_218), .B(n_219), .Y(n_217) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
INVx1_ASAP7_75t_L g220 ( .A(n_210), .Y(n_220) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_210), .A2(n_470), .B(n_481), .Y(n_469) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_210), .A2(n_493), .B(n_501), .Y(n_492) );
INVx2_ASAP7_75t_L g257 ( .A(n_213), .Y(n_257) );
AND2x2_ASAP7_75t_L g303 ( .A(n_213), .B(n_224), .Y(n_303) );
AND2x2_ASAP7_75t_L g313 ( .A(n_213), .B(n_238), .Y(n_313) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_220), .B(n_221), .Y(n_213) );
INVx2_ASAP7_75t_L g433 ( .A(n_223), .Y(n_433) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_224), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g274 ( .A(n_224), .Y(n_274) );
AND2x2_ASAP7_75t_L g318 ( .A(n_224), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g334 ( .A(n_224), .B(n_297), .Y(n_334) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
AND2x2_ASAP7_75t_L g296 ( .A(n_225), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g347 ( .A(n_225), .B(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_225), .B(n_257), .Y(n_379) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .Y(n_229) );
AND2x2_ASAP7_75t_L g258 ( .A(n_237), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g319 ( .A(n_237), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_237), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g356 ( .A(n_237), .Y(n_356) );
INVx1_ASAP7_75t_L g389 ( .A(n_237), .Y(n_389) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g267 ( .A(n_238), .B(n_257), .Y(n_267) );
INVx1_ASAP7_75t_L g297 ( .A(n_238), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g474 ( .A(n_244), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_244), .A2(n_536), .B(n_537), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B1(n_260), .B2(n_267), .C(n_268), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_251), .B(n_271), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_251), .B(n_334), .Y(n_411) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_253), .B(n_301), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_253), .B(n_262), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_253), .B(n_276), .Y(n_405) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g327 ( .A(n_257), .Y(n_327) );
AND2x2_ASAP7_75t_L g302 ( .A(n_258), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g380 ( .A(n_258), .Y(n_380) );
AND2x2_ASAP7_75t_L g312 ( .A(n_259), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_259), .B(n_282), .Y(n_328) );
AND2x2_ASAP7_75t_L g392 ( .A(n_259), .B(n_318), .Y(n_392) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g301 ( .A(n_263), .B(n_270), .Y(n_301) );
AND2x2_ASAP7_75t_L g397 ( .A(n_264), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_266), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_267), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_267), .B(n_274), .Y(n_362) );
AND2x2_ASAP7_75t_L g382 ( .A(n_267), .B(n_282), .Y(n_382) );
AND2x2_ASAP7_75t_L g403 ( .A(n_267), .B(n_347), .Y(n_403) );
OAI32xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .A3(n_274), .B1(n_275), .B2(n_278), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
INVx1_ASAP7_75t_SL g276 ( .A(n_270), .Y(n_276) );
NAND2x1_ASAP7_75t_L g317 ( .A(n_270), .B(n_300), .Y(n_317) );
OR2x2_ASAP7_75t_L g321 ( .A(n_270), .B(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_270), .B(n_369), .Y(n_422) );
INVx1_ASAP7_75t_L g290 ( .A(n_271), .Y(n_290) );
OAI221xp5_ASAP7_75t_SL g408 ( .A1(n_272), .A2(n_363), .B1(n_409), .B2(n_412), .C(n_413), .Y(n_408) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g280 ( .A(n_273), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g323 ( .A(n_273), .B(n_296), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_273), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g401 ( .A(n_273), .B(n_334), .Y(n_401) );
INVxp67_ASAP7_75t_L g337 ( .A(n_274), .Y(n_337) );
OR2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
AND2x2_ASAP7_75t_L g407 ( .A(n_276), .B(n_394), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_276), .B(n_357), .Y(n_430) );
INVx1_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_278), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g423 ( .A(n_278), .B(n_424), .Y(n_423) );
OAI21xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_283), .B(n_286), .Y(n_279) );
AND2x2_ASAP7_75t_L g292 ( .A(n_281), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g376 ( .A(n_285), .B(n_296), .Y(n_376) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g394 ( .A(n_287), .B(n_352), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_287), .B(n_351), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_288), .B(n_300), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B(n_294), .C(n_304), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_290), .A2(n_325), .B1(n_329), .B2(n_332), .C(n_335), .Y(n_324) );
AOI31xp33_ASAP7_75t_L g419 ( .A1(n_290), .A2(n_420), .A3(n_421), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_298), .B1(n_300), .B2(n_302), .Y(n_294) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g420 ( .A(n_300), .Y(n_420) );
INVx1_ASAP7_75t_L g383 ( .A(n_301), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_303), .A2(n_427), .B(n_429), .C(n_431), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_308), .B2(n_312), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_309), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_311), .A2(n_345), .B1(n_364), .B2(n_400), .C(n_402), .Y(n_399) );
INVx1_ASAP7_75t_L g395 ( .A(n_312), .Y(n_395) );
INVx1_ASAP7_75t_L g349 ( .A(n_313), .Y(n_349) );
NAND3xp33_ASAP7_75t_SL g314 ( .A(n_315), .B(n_324), .C(n_339), .Y(n_314) );
OAI21xp33_ASAP7_75t_L g365 ( .A1(n_316), .A2(n_366), .B(n_370), .Y(n_365) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_318), .B(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g425 ( .A(n_319), .Y(n_425) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g363 ( .A(n_326), .B(n_346), .Y(n_363) );
INVx1_ASAP7_75t_L g338 ( .A(n_327), .Y(n_338) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g336 ( .A(n_330), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_330), .B(n_368), .Y(n_367) );
NOR4xp25_ASAP7_75t_L g335 ( .A(n_331), .B(n_336), .C(n_337), .D(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AOI222xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_344), .B1(n_350), .B2(n_351), .C1(n_353), .C2(n_357), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g437 ( .A(n_341), .Y(n_437) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_349), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_353), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_358), .A2(n_414), .B(n_416), .Y(n_413) );
NOR4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_371), .C(n_384), .D(n_399), .Y(n_359) );
OAI221xp5_ASAP7_75t_SL g360 ( .A1(n_361), .A2(n_362), .B1(n_363), .B2(n_364), .C(n_365), .Y(n_360) );
INVx1_ASAP7_75t_L g440 ( .A(n_361), .Y(n_440) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_368), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
OAI222xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_375), .B1(n_377), .B2(n_378), .C1(n_381), .C2(n_383), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AOI211xp5_ASAP7_75t_L g406 ( .A1(n_376), .A2(n_407), .B(n_408), .C(n_419), .Y(n_406) );
OR2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_390), .B1(n_391), .B2(n_393), .C1(n_395), .C2(n_396), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_401), .A2(n_404), .B1(n_437), .B2(n_438), .Y(n_436) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI211xp5_ASAP7_75t_SL g431 ( .A1(n_432), .A2(n_434), .B(n_436), .C(n_439), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_443), .Y(n_449) );
NOR2x2_ASAP7_75t_L g760 ( .A(n_444), .B(n_459), .Y(n_760) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g458 ( .A(n_445), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
OAI21xp5_ASAP7_75t_SL g451 ( .A1(n_448), .A2(n_452), .B(n_762), .Y(n_451) );
NOR2xp33_ASAP7_75t_SL g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_456), .B1(n_457), .B2(n_460), .Y(n_453) );
INVx2_ASAP7_75t_L g754 ( .A(n_454), .Y(n_754) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx6_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g755 ( .A(n_458), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_460), .Y(n_756) );
AND2x2_ASAP7_75t_SL g460 ( .A(n_461), .B(n_717), .Y(n_460) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_621), .C(n_705), .Y(n_461) );
NAND4xp25_ASAP7_75t_L g462 ( .A(n_463), .B(n_564), .C(n_586), .D(n_602), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_502), .B1(n_525), .B2(n_543), .C(n_550), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_482), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_466), .B(n_543), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_466), .B(n_604), .C(n_617), .D(n_619), .Y(n_616) );
INVxp67_ASAP7_75t_L g733 ( .A(n_466), .Y(n_733) );
INVx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g615 ( .A(n_467), .B(n_553), .Y(n_615) );
AND2x2_ASAP7_75t_L g639 ( .A(n_467), .B(n_482), .Y(n_639) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AND2x2_ASAP7_75t_L g606 ( .A(n_468), .B(n_542), .Y(n_606) );
AND2x2_ASAP7_75t_L g646 ( .A(n_468), .B(n_627), .Y(n_646) );
AND2x2_ASAP7_75t_L g663 ( .A(n_468), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_468), .B(n_483), .Y(n_687) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g541 ( .A(n_469), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g558 ( .A(n_469), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_483), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_469), .B(n_492), .Y(n_592) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B(n_479), .C(n_480), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_480), .A2(n_489), .B(n_490), .Y(n_488) );
AND2x2_ASAP7_75t_L g573 ( .A(n_482), .B(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_482), .A2(n_623), .B1(n_626), .B2(n_628), .C(n_632), .Y(n_622) );
AND2x2_ASAP7_75t_L g681 ( .A(n_482), .B(n_646), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_482), .B(n_663), .Y(n_715) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_492), .Y(n_482) );
INVx3_ASAP7_75t_L g542 ( .A(n_483), .Y(n_542) );
AND2x2_ASAP7_75t_L g590 ( .A(n_483), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g644 ( .A(n_483), .B(n_559), .Y(n_644) );
AND2x2_ASAP7_75t_L g702 ( .A(n_483), .B(n_703), .Y(n_702) );
AND2x2_ASAP7_75t_L g543 ( .A(n_492), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
INVx1_ASAP7_75t_L g614 ( .A(n_492), .Y(n_614) );
HB1xp67_ASAP7_75t_L g620 ( .A(n_492), .Y(n_620) );
AND2x2_ASAP7_75t_L g665 ( .A(n_492), .B(n_542), .Y(n_665) );
OR2x2_ASAP7_75t_L g704 ( .A(n_492), .B(n_544), .Y(n_704) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_502), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_510), .Y(n_502) );
AND2x2_ASAP7_75t_L g700 ( .A(n_503), .B(n_697), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_503), .B(n_682), .Y(n_732) );
BUFx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g631 ( .A(n_504), .B(n_555), .Y(n_631) );
AND2x2_ASAP7_75t_L g680 ( .A(n_504), .B(n_528), .Y(n_680) );
INVx1_ASAP7_75t_L g726 ( .A(n_504), .Y(n_726) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_505), .Y(n_540) );
AND2x2_ASAP7_75t_L g581 ( .A(n_505), .B(n_555), .Y(n_581) );
INVx1_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
AND2x2_ASAP7_75t_L g604 ( .A(n_505), .B(n_521), .Y(n_604) );
AND2x2_ASAP7_75t_L g672 ( .A(n_510), .B(n_580), .Y(n_672) );
INVx2_ASAP7_75t_L g737 ( .A(n_510), .Y(n_737) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
AND2x2_ASAP7_75t_L g554 ( .A(n_511), .B(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g567 ( .A(n_511), .B(n_529), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_511), .B(n_528), .Y(n_595) );
INVx1_ASAP7_75t_L g601 ( .A(n_511), .Y(n_601) );
INVx1_ASAP7_75t_L g618 ( .A(n_511), .Y(n_618) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_511), .Y(n_630) );
INVx2_ASAP7_75t_L g698 ( .A(n_511), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_516), .Y(n_513) );
INVx2_ASAP7_75t_L g555 ( .A(n_521), .Y(n_555) );
BUFx2_ASAP7_75t_L g652 ( .A(n_521), .Y(n_652) );
AND2x2_ASAP7_75t_L g697 ( .A(n_521), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_539), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_527), .B(n_634), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_527), .A2(n_696), .B(n_710), .Y(n_720) );
AND2x2_ASAP7_75t_L g745 ( .A(n_527), .B(n_631), .Y(n_745) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g667 ( .A(n_529), .Y(n_667) );
AND2x2_ASAP7_75t_L g696 ( .A(n_529), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
INVx2_ASAP7_75t_L g599 ( .A(n_530), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_530), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
INVx2_ASAP7_75t_L g553 ( .A(n_540), .Y(n_553) );
OR2x2_ASAP7_75t_L g566 ( .A(n_540), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g634 ( .A(n_540), .B(n_630), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_540), .B(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g735 ( .A(n_540), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_540), .B(n_672), .Y(n_747) );
AND2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g649 ( .A(n_541), .B(n_543), .Y(n_649) );
INVx2_ASAP7_75t_L g561 ( .A(n_542), .Y(n_561) );
AND2x2_ASAP7_75t_L g589 ( .A(n_542), .B(n_562), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_542), .B(n_614), .Y(n_670) );
AND2x2_ASAP7_75t_L g584 ( .A(n_543), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g731 ( .A(n_543), .Y(n_731) );
AND2x2_ASAP7_75t_L g743 ( .A(n_543), .B(n_606), .Y(n_743) );
AND2x2_ASAP7_75t_L g569 ( .A(n_544), .B(n_559), .Y(n_569) );
INVx1_ASAP7_75t_L g664 ( .A(n_544), .Y(n_664) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g562 ( .A(n_549), .B(n_563), .Y(n_562) );
INVxp67_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_556), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_553), .B(n_600), .Y(n_609) );
OR2x2_ASAP7_75t_L g741 ( .A(n_553), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g658 ( .A(n_554), .B(n_599), .Y(n_658) );
AND2x2_ASAP7_75t_L g666 ( .A(n_554), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g725 ( .A(n_554), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g749 ( .A(n_554), .B(n_596), .Y(n_749) );
NOR2xp67_ASAP7_75t_L g707 ( .A(n_555), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g736 ( .A(n_555), .B(n_599), .Y(n_736) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2x1p5_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
AND2x2_ASAP7_75t_L g588 ( .A(n_558), .B(n_589), .Y(n_588) );
INVxp67_ASAP7_75t_L g750 ( .A(n_558), .Y(n_750) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVx1_ASAP7_75t_L g585 ( .A(n_561), .Y(n_585) );
AND2x2_ASAP7_75t_L g636 ( .A(n_561), .B(n_569), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_561), .B(n_704), .Y(n_730) );
INVx2_ASAP7_75t_L g575 ( .A(n_562), .Y(n_575) );
INVx3_ASAP7_75t_L g627 ( .A(n_562), .Y(n_627) );
OR2x2_ASAP7_75t_L g655 ( .A(n_562), .B(n_656), .Y(n_655) );
AOI311xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_568), .A3(n_570), .B(n_571), .C(n_582), .Y(n_564) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_565), .A2(n_603), .B(n_605), .C(n_607), .Y(n_602) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g587 ( .A(n_567), .Y(n_587) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g605 ( .A(n_569), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_569), .B(n_585), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_569), .B(n_570), .Y(n_738) );
AND2x2_ASAP7_75t_L g660 ( .A(n_570), .B(n_574), .Y(n_660) );
AOI21xp33_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g718 ( .A(n_574), .B(n_606), .Y(n_718) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_575), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
AND2x2_ASAP7_75t_L g603 ( .A(n_579), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g648 ( .A(n_581), .Y(n_648) );
AND2x4_ASAP7_75t_L g710 ( .A(n_581), .B(n_679), .Y(n_710) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_584), .A2(n_650), .B1(n_662), .B2(n_666), .C1(n_668), .C2(n_672), .Y(n_661) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_590), .C(n_593), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_587), .B(n_631), .Y(n_654) );
INVx1_ASAP7_75t_L g676 ( .A(n_589), .Y(n_676) );
INVx1_ASAP7_75t_L g610 ( .A(n_591), .Y(n_610) );
OR2x2_ASAP7_75t_L g675 ( .A(n_592), .B(n_676), .Y(n_675) );
OAI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B(n_600), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_594), .B(n_612), .C(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_594), .A2(n_631), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_598), .Y(n_651) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_599), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g708 ( .A(n_599), .Y(n_708) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_599), .Y(n_724) );
INVx2_ASAP7_75t_L g682 ( .A(n_600), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_604), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g656 ( .A(n_606), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_610), .B1(n_611), .B2(n_615), .C(n_616), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_610), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g744 ( .A(n_610), .Y(n_744) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g625 ( .A(n_617), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_617), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g683 ( .A(n_617), .B(n_631), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_617), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g716 ( .A(n_617), .B(n_651), .Y(n_716) );
BUFx3_ASAP7_75t_L g679 ( .A(n_618), .Y(n_679) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND5xp2_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .C(n_661), .D(n_673), .E(n_688), .Y(n_621) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AOI32xp33_ASAP7_75t_L g713 ( .A1(n_625), .A2(n_652), .A3(n_668), .B1(n_714), .B2(n_716), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_627), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g637 ( .A(n_631), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_647), .B1(n_649), .B2(n_650), .C(n_653), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g712 ( .A(n_644), .B(n_663), .Y(n_712) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_649), .A2(n_710), .B1(n_728), .B2(n_733), .C(n_734), .Y(n_727) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx2_ASAP7_75t_L g693 ( .A(n_652), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_657), .B2(n_659), .Y(n_653) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g671 ( .A(n_663), .Y(n_671) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .B1(n_681), .B2(n_682), .C1(n_683), .C2(n_684), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g728 ( .A1(n_682), .A2(n_729), .B1(n_731), .B2(n_732), .Y(n_728) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_694), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_699), .B(n_701), .Y(n_694) );
INVx2_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g742 ( .A(n_697), .Y(n_742) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_709), .B(n_711), .C(n_713), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI211xp5_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_721), .C(n_746), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_718), .Y(n_722) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
OAI211xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_727), .C(n_739), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B(n_738), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_743), .B1(n_744), .B2(n_745), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
endmodule