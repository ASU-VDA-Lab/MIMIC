module fake_ibex_796_n_4275 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_805, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_232, n_380, n_749, n_281, n_559, n_425, n_4275);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4275;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_3559;
wire n_4158;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_1722;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_2230;
wire n_1782;
wire n_963;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_3904;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2605;
wire n_2343;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_1636;
wire n_939;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3753;
wire n_3896;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3395;
wire n_3242;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3509;
wire n_3472;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3949;
wire n_3507;
wire n_3884;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_2436;
wire n_1663;
wire n_2705;
wire n_1214;
wire n_1274;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_3699;
wire n_1955;
wire n_3668;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_3022;
wire n_3148;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_3973;
wire n_1313;
wire n_4214;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_810;
wire n_1401;
wire n_3764;
wire n_4173;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_1620;
wire n_869;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_4188;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2899;
wire n_2826;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1764;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2625;
wire n_2350;
wire n_1742;
wire n_2444;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2646;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3800;
wire n_3963;
wire n_3461;
wire n_2445;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4103;
wire n_3583;
wire n_2019;
wire n_4126;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_822;
wire n_1042;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2718;
wire n_2377;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_3788;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_4096;
wire n_3634;
wire n_1377;
wire n_2473;
wire n_3524;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_3054;
wire n_2924;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_1140;
wire n_1985;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_3790;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_2573;
wire n_1237;
wire n_2880;
wire n_2390;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_3855;
wire n_4033;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1890;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1990;
wire n_1179;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_2999;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_1345;
wire n_4215;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3470;
wire n_3584;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3797;
wire n_998;
wire n_1395;
wire n_1729;
wire n_1115;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_814;
wire n_3829;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1523;
wire n_1086;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_2570;
wire n_4051;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_3719;
wire n_3948;
wire n_1539;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_2711;
wire n_2842;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_3646;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_2193;
wire n_817;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_2716;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_3735;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_4052;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_836;
wire n_1475;
wire n_3316;
wire n_2465;
wire n_1263;
wire n_3337;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1683;
wire n_1185;
wire n_4256;
wire n_3575;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_831;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1845;
wire n_1667;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2684;
wire n_3284;
wire n_2524;
wire n_2875;
wire n_1437;
wire n_3835;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1941;
wire n_1707;
wire n_3902;
wire n_3927;
wire n_2422;
wire n_4185;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_4133;
wire n_920;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_991;
wire n_961;
wire n_2127;
wire n_1223;
wire n_3747;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_3552;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_3100;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1601;
wire n_1294;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4142;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_4007;
wire n_3960;
wire n_3608;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1348;
wire n_838;
wire n_1289;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_4149;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_3930;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_1396;
wire n_2916;
wire n_1923;
wire n_1224;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_3745;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_3907;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_3746;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_1603;
wire n_935;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_3044;
wire n_2868;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_950;
wire n_3139;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_3619;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_3604;
wire n_833;
wire n_3649;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2093;
wire n_2348;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_2366;
wire n_4229;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_2898;
wire n_2232;
wire n_3121;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1809;
wire n_1206;
wire n_855;
wire n_2367;
wire n_812;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2667;
wire n_1050;
wire n_2218;
wire n_2553;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1542;
wire n_1547;
wire n_1586;
wire n_1362;
wire n_946;
wire n_3497;
wire n_4178;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3586;
wire n_956;
wire n_3561;
wire n_4125;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1887;
wire n_1212;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1584;
wire n_1481;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_4235;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3403;
wire n_1363;
wire n_3863;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_3102;
wire n_2790;
wire n_2872;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_3343;
wire n_3752;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_3543;
wire n_1734;
wire n_3655;
wire n_3742;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_2371;
wire n_914;
wire n_3992;
wire n_4147;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2140;
wire n_2013;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_3296;
wire n_1911;
wire n_2293;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3318;
wire n_3223;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_1193;
wire n_849;
wire n_980;
wire n_3067;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3380;
wire n_1074;
wire n_2928;
wire n_3557;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_2982;
wire n_999;
wire n_2634;
wire n_3124;
wire n_3286;
wire n_1092;
wire n_4038;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1385;
wire n_1142;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_2653;
wire n_2357;
wire n_2303;
wire n_2618;
wire n_2855;
wire n_3938;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_2302;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_3189;
wire n_2443;
wire n_3052;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_2961;
wire n_2996;
wire n_2704;
wire n_2770;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3582;
wire n_3689;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_990;
wire n_1383;
wire n_3675;
wire n_1968;
wire n_4108;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3562;
wire n_3933;
wire n_955;
wire n_1916;
wire n_1333;
wire n_2726;
wire n_2917;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_3758;
wire n_3988;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1696;
wire n_1277;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3635;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1678;
wire n_1780;
wire n_1091;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_1655;
wire n_984;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

INVx1_ASAP7_75t_L g808 ( 
.A(n_153),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_56),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_285),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_7),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_166),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_193),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_180),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_504),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_113),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_464),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_22),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_601),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_779),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_464),
.Y(n_821)
);

BUFx10_ASAP7_75t_L g822 ( 
.A(n_180),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_28),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_638),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_169),
.Y(n_825)
);

CKINVDCx16_ASAP7_75t_R g826 ( 
.A(n_785),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_530),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_201),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_196),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_509),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_761),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_216),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_228),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_426),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_505),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_132),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_118),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_568),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_780),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_252),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_646),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_226),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_94),
.Y(n_843)
);

CKINVDCx20_ASAP7_75t_R g844 ( 
.A(n_191),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_467),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_346),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_110),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_23),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_697),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_86),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_444),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_49),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_538),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_793),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_411),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_423),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_798),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_57),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_153),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_771),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_3),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_175),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_634),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_372),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_314),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_457),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_353),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_252),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_300),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_190),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_561),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_181),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_201),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_304),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_629),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_778),
.Y(n_876)
);

INVx1_ASAP7_75t_SL g877 ( 
.A(n_703),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_659),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_435),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_569),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_786),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_658),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_403),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_435),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_206),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_633),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_523),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_674),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_417),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_223),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_160),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_336),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_681),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_22),
.Y(n_894)
);

BUFx10_ASAP7_75t_L g895 ( 
.A(n_207),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_273),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_564),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_541),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_68),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_228),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_2),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_657),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_670),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_789),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_358),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_597),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_572),
.Y(n_907)
);

CKINVDCx16_ASAP7_75t_R g908 ( 
.A(n_359),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_88),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_767),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_640),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_342),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_807),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_8),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_337),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_689),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_565),
.Y(n_917)
);

BUFx10_ASAP7_75t_L g918 ( 
.A(n_479),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_205),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_38),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_258),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_787),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_498),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_127),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_51),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_31),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_194),
.Y(n_927)
);

BUFx10_ASAP7_75t_L g928 ( 
.A(n_19),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_429),
.Y(n_929)
);

BUFx2_ASAP7_75t_L g930 ( 
.A(n_459),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_107),
.Y(n_931)
);

BUFx8_ASAP7_75t_SL g932 ( 
.A(n_523),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_402),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_727),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_166),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_472),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_324),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_680),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_407),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_608),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_218),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_711),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_674),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_2),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_432),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_187),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_492),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_335),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_394),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_702),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_279),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_534),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_381),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_733),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_425),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_235),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_506),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_76),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_624),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_139),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_100),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_727),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_221),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_771),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_757),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_125),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_732),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_659),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_132),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_588),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_562),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_503),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_617),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_762),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_177),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_571),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_436),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_221),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_63),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_309),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_541),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_119),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_775),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_299),
.Y(n_984)
);

INVx1_ASAP7_75t_SL g985 ( 
.A(n_800),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_699),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_13),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_619),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_143),
.Y(n_989)
);

BUFx5_ASAP7_75t_L g990 ( 
.A(n_694),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_747),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_194),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_756),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_162),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_349),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_798),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_734),
.Y(n_997)
);

CKINVDCx20_ASAP7_75t_R g998 ( 
.A(n_611),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_37),
.Y(n_999)
);

CKINVDCx20_ASAP7_75t_R g1000 ( 
.A(n_338),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_656),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_91),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_362),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_563),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_408),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_45),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_419),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_627),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_162),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_612),
.Y(n_1010)
);

BUFx10_ASAP7_75t_L g1011 ( 
.A(n_331),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_359),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_769),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_586),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_122),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_680),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_368),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_404),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_418),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_770),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_613),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_366),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_560),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_495),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_181),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_297),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_709),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_465),
.Y(n_1028)
);

BUFx10_ASAP7_75t_L g1029 ( 
.A(n_638),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_768),
.Y(n_1030)
);

CKINVDCx20_ASAP7_75t_R g1031 ( 
.A(n_634),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_429),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_748),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_719),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_209),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_737),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_97),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_481),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_117),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_724),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_702),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_65),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_375),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_154),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_310),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_478),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_785),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_371),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_515),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_543),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_148),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_484),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_774),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_27),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_36),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_693),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_58),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_666),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_689),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_772),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_573),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_531),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_40),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_795),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_4),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_802),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_377),
.Y(n_1067)
);

BUFx10_ASAP7_75t_L g1068 ( 
.A(n_690),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_764),
.Y(n_1069)
);

BUFx10_ASAP7_75t_L g1070 ( 
.A(n_307),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_759),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_191),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_489),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_788),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_758),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_129),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_679),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_182),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_443),
.Y(n_1079)
);

BUFx10_ASAP7_75t_L g1080 ( 
.A(n_603),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_447),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_26),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_60),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_753),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_176),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_461),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_721),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_184),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_614),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_516),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_763),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_129),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_282),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_193),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_114),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_85),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_263),
.Y(n_1097)
);

CKINVDCx14_ASAP7_75t_R g1098 ( 
.A(n_239),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_184),
.Y(n_1099)
);

INVx1_ASAP7_75t_SL g1100 ( 
.A(n_399),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_172),
.Y(n_1101)
);

CKINVDCx14_ASAP7_75t_R g1102 ( 
.A(n_353),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_789),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_264),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_458),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_649),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_787),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_449),
.Y(n_1108)
);

BUFx5_ASAP7_75t_L g1109 ( 
.A(n_593),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_79),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_553),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_513),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_212),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_244),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_710),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_519),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_688),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_465),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_66),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_579),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_313),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_676),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_784),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_165),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_569),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_367),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_667),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_633),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_613),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_670),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_652),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_521),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_118),
.Y(n_1133)
);

BUFx5_ASAP7_75t_L g1134 ( 
.A(n_367),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_778),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_547),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_671),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_223),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_782),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_420),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_351),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_321),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_356),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_783),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_402),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_185),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_477),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_421),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_365),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_383),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_760),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_612),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_628),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_87),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_135),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_261),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_556),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_765),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_274),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_597),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_703),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_327),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_664),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_269),
.Y(n_1164)
);

BUFx2_ASAP7_75t_L g1165 ( 
.A(n_63),
.Y(n_1165)
);

BUFx8_ASAP7_75t_SL g1166 ( 
.A(n_678),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_373),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_249),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_700),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_496),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_765),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_556),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_448),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_580),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_254),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_287),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_550),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_155),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_159),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_777),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_44),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_226),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_344),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_19),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_152),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_325),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_713),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_66),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_476),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_23),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_584),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_699),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_90),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_146),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_405),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_535),
.Y(n_1196)
);

CKINVDCx16_ASAP7_75t_R g1197 ( 
.A(n_742),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_107),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_708),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_677),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_90),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_342),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_794),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_536),
.Y(n_1204)
);

CKINVDCx14_ASAP7_75t_R g1205 ( 
.A(n_116),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_408),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_188),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_781),
.Y(n_1208)
);

CKINVDCx14_ASAP7_75t_R g1209 ( 
.A(n_122),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_42),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_732),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_276),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_600),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_220),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_807),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_415),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_790),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_473),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_721),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_520),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_594),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_607),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_329),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_207),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_8),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_729),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_97),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_8),
.Y(n_1228)
);

BUFx5_ASAP7_75t_L g1229 ( 
.A(n_319),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_443),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_400),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_608),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_627),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_35),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_773),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_389),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_481),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_417),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_796),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_454),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_14),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_639),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_497),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_332),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_776),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_321),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_562),
.Y(n_1248)
);

CKINVDCx14_ASAP7_75t_R g1249 ( 
.A(n_729),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_52),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_35),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_30),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_436),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_73),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_660),
.Y(n_1255)
);

CKINVDCx20_ASAP7_75t_R g1256 ( 
.A(n_127),
.Y(n_1256)
);

CKINVDCx14_ASAP7_75t_R g1257 ( 
.A(n_701),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_337),
.Y(n_1258)
);

INVx1_ASAP7_75t_SL g1259 ( 
.A(n_24),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_69),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_276),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_24),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_578),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_88),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_93),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_346),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_790),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_323),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_315),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_576),
.Y(n_1270)
);

BUFx8_ASAP7_75t_SL g1271 ( 
.A(n_296),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_376),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_489),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_147),
.Y(n_1274)
);

BUFx10_ASAP7_75t_L g1275 ( 
.A(n_573),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_488),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_520),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_293),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_755),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_685),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_477),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_365),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_791),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_131),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_766),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_792),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_619),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_479),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_23),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_418),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_563),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_549),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_55),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_327),
.Y(n_1294)
);

BUFx10_ASAP7_75t_L g1295 ( 
.A(n_95),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_14),
.Y(n_1296)
);

BUFx3_ASAP7_75t_L g1297 ( 
.A(n_76),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_137),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_66),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_590),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_781),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_718),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_35),
.Y(n_1303)
);

INVxp67_ASAP7_75t_L g1304 ( 
.A(n_1165),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_861),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_930),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_809),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_829),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_829),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_809),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_924),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1054),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_933),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_990),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_924),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_960),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1184),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_960),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_945),
.B(n_1),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_970),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1098),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_818),
.Y(n_1322)
);

INVxp67_ASAP7_75t_SL g1323 ( 
.A(n_1083),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_970),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_818),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1008),
.B(n_0),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_823),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_823),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1172),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1172),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1113),
.B(n_0),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_852),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1186),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1186),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1214),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_826),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1102),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1214),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1205),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_852),
.Y(n_1340)
);

INVxp33_ASAP7_75t_L g1341 ( 
.A(n_828),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_858),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1272),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1083),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_875),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1272),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_858),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_860),
.B(n_0),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_868),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_1241),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1209),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1241),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_1243),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_811),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1243),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_1249),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_920),
.Y(n_1357)
);

CKINVDCx20_ASAP7_75t_R g1358 ( 
.A(n_1257),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_990),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_928),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_944),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_987),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_908),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1021),
.Y(n_1364)
);

CKINVDCx16_ASAP7_75t_R g1365 ( 
.A(n_928),
.Y(n_1365)
);

CKINVDCx20_ASAP7_75t_R g1366 ( 
.A(n_1197),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1119),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1250),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1250),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1251),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_868),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_928),
.Y(n_1373)
);

INVxp67_ASAP7_75t_L g1374 ( 
.A(n_1251),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_822),
.B(n_1),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1262),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1262),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1293),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_1293),
.Y(n_1379)
);

CKINVDCx20_ASAP7_75t_R g1380 ( 
.A(n_1296),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_1296),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1299),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1299),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_894),
.Y(n_1384)
);

INVxp67_ASAP7_75t_SL g1385 ( 
.A(n_907),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_932),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1166),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1271),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1303),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_907),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_901),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1045),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_914),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_808),
.B(n_3),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_925),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_822),
.B(n_2),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1045),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1090),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_822),
.B(n_3),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_926),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1090),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_979),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_817),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1215),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_990),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_999),
.Y(n_1406)
);

INVxp33_ASAP7_75t_L g1407 ( 
.A(n_810),
.Y(n_1407)
);

CKINVDCx16_ASAP7_75t_R g1408 ( 
.A(n_838),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1215),
.Y(n_1409)
);

CKINVDCx16_ASAP7_75t_R g1410 ( 
.A(n_838),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1006),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1042),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1232),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1232),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1297),
.Y(n_1415)
);

INVxp67_ASAP7_75t_SL g1416 ( 
.A(n_1297),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_820),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_831),
.Y(n_1418)
);

BUFx3_ASAP7_75t_L g1419 ( 
.A(n_990),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_810),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_812),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_812),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1055),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1057),
.Y(n_1424)
);

HB1xp67_ASAP7_75t_L g1425 ( 
.A(n_1063),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_836),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_836),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_846),
.Y(n_1428)
);

INVxp33_ASAP7_75t_SL g1429 ( 
.A(n_1065),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_846),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1082),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_883),
.Y(n_1432)
);

NOR2xp67_ASAP7_75t_L g1433 ( 
.A(n_883),
.B(n_4),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_884),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_844),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1374),
.B(n_1181),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1349),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1323),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1345),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1376),
.B(n_1188),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1371),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1304),
.B(n_838),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1371),
.Y(n_1443)
);

BUFx8_ASAP7_75t_L g1444 ( 
.A(n_1319),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1344),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1308),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1379),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1307),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1379),
.Y(n_1449)
);

XOR2xp5_ASAP7_75t_L g1450 ( 
.A(n_1312),
.B(n_866),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1345),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1360),
.B(n_1210),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1349),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1345),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1309),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1380),
.Y(n_1456)
);

BUFx6f_ASAP7_75t_L g1457 ( 
.A(n_1345),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1380),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_R g1459 ( 
.A(n_1365),
.B(n_1225),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1419),
.Y(n_1460)
);

NOR3xp33_ASAP7_75t_L g1461 ( 
.A(n_1375),
.B(n_1190),
.C(n_848),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1305),
.B(n_884),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1310),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1311),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1341),
.B(n_895),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1419),
.Y(n_1466)
);

NAND2x1_ASAP7_75t_L g1467 ( 
.A(n_1373),
.B(n_936),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_1322),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1314),
.Y(n_1469)
);

BUFx8_ASAP7_75t_L g1470 ( 
.A(n_1394),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1315),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_SL g1472 ( 
.A(n_1341),
.B(n_1228),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1314),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1325),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1359),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1312),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1332),
.B(n_936),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1378),
.B(n_895),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1327),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1316),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1328),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1359),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1306),
.B(n_1313),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1318),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1384),
.B(n_1234),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1340),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1320),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1317),
.A2(n_1288),
.B1(n_897),
.B2(n_912),
.Y(n_1488)
);

BUFx6f_ASAP7_75t_L g1489 ( 
.A(n_1405),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1324),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1342),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1317),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1403),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1405),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1347),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1329),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1400),
.B(n_1406),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1350),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1330),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_R g1500 ( 
.A(n_1321),
.B(n_813),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1333),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_1352),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1354),
.A2(n_966),
.B(n_952),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_R g1504 ( 
.A(n_1337),
.B(n_813),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1425),
.B(n_814),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1334),
.B(n_885),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1403),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1353),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1335),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1355),
.Y(n_1510)
);

AND2x6_ASAP7_75t_L g1511 ( 
.A(n_1396),
.B(n_875),
.Y(n_1511)
);

CKINVDCx20_ASAP7_75t_R g1512 ( 
.A(n_1417),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1420),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1368),
.Y(n_1514)
);

BUFx6f_ASAP7_75t_L g1515 ( 
.A(n_1421),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_1370),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1338),
.Y(n_1517)
);

AND3x2_ASAP7_75t_L g1518 ( 
.A(n_1399),
.B(n_832),
.C(n_824),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1343),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_1377),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1346),
.B(n_952),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1381),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1408),
.B(n_1259),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1390),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1422),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1392),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1382),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1397),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1383),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1398),
.Y(n_1530)
);

BUFx8_ASAP7_75t_L g1531 ( 
.A(n_1410),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1389),
.Y(n_1532)
);

HB1xp67_ASAP7_75t_L g1533 ( 
.A(n_1391),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1429),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1393),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1401),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1417),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1418),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1426),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1404),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1409),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1407),
.B(n_895),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1413),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1414),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1415),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1395),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1427),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1432),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1402),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1411),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1412),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1407),
.B(n_918),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_1418),
.Y(n_1553)
);

BUFx6f_ASAP7_75t_L g1554 ( 
.A(n_1428),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1357),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1430),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1423),
.B(n_990),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1435),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1434),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1336),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1336),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1361),
.B(n_886),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1424),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1362),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1431),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1367),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_R g1567 ( 
.A(n_1339),
.B(n_814),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1369),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1372),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_1363),
.Y(n_1570)
);

CKINVDCx20_ASAP7_75t_R g1571 ( 
.A(n_1363),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1364),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1364),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1385),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1416),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1433),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1366),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1348),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1366),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1326),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1331),
.B(n_966),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1386),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1351),
.B(n_815),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1387),
.B(n_1289),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1356),
.B(n_991),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1388),
.Y(n_1586)
);

NAND2xp33_ASAP7_75t_L g1587 ( 
.A(n_1358),
.B(n_990),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_1371),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1371),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1365),
.B(n_990),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1371),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_R g1592 ( 
.A(n_1365),
.B(n_815),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1323),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1371),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1365),
.B(n_990),
.Y(n_1595)
);

NAND2xp33_ASAP7_75t_R g1596 ( 
.A(n_1310),
.B(n_816),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1310),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1305),
.B(n_991),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1323),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1349),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1349),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1371),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1323),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1371),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1345),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1371),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_1371),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1349),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1323),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1374),
.B(n_816),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1349),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1349),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1304),
.B(n_918),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1323),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1314),
.A2(n_1088),
.B(n_1075),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1371),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1371),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1349),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1323),
.Y(n_1619)
);

AOI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1310),
.A2(n_821),
.B1(n_825),
.B2(n_819),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1310),
.A2(n_821),
.B1(n_825),
.B2(n_819),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1305),
.B(n_1075),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1323),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1323),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1323),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1323),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1349),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1307),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1349),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1323),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1323),
.B(n_1109),
.Y(n_1631)
);

CKINVDCx5p33_ASAP7_75t_R g1632 ( 
.A(n_1371),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1323),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1371),
.Y(n_1634)
);

HB1xp67_ASAP7_75t_L g1635 ( 
.A(n_1310),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1304),
.B(n_1302),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1371),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1349),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1371),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1310),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_1371),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1323),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1349),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1323),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1323),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1349),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1323),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1305),
.B(n_1088),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1310),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1323),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1323),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1578),
.B(n_887),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1513),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1436),
.B(n_888),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1503),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1580),
.A2(n_840),
.B1(n_841),
.B2(n_839),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1503),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1542),
.B(n_918),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1600),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1552),
.Y(n_1661)
);

NOR2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1534),
.B(n_827),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1477),
.B(n_843),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1461),
.B(n_830),
.C(n_827),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1600),
.Y(n_1665)
);

INVx5_ASAP7_75t_L g1666 ( 
.A(n_1513),
.Y(n_1666)
);

INVx3_ASAP7_75t_L g1667 ( 
.A(n_1513),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1465),
.B(n_1011),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1501),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1601),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1523),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1601),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1483),
.B(n_1011),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1459),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1483),
.B(n_830),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1564),
.B(n_1438),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_L g1677 ( 
.A(n_1511),
.B(n_1109),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1509),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1517),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1564),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1446),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1483),
.B(n_1011),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1515),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1455),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1464),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1515),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1440),
.B(n_1452),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1497),
.B(n_833),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1515),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_L g1690 ( 
.A(n_1488),
.B(n_964),
.C(n_877),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1471),
.Y(n_1691)
);

BUFx6f_ASAP7_75t_L g1692 ( 
.A(n_1525),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1445),
.B(n_1109),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1448),
.B(n_1029),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1480),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1484),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1487),
.Y(n_1697)
);

INVx3_ASAP7_75t_L g1698 ( 
.A(n_1525),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1485),
.B(n_1610),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1555),
.B(n_875),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1628),
.B(n_1029),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1490),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1477),
.B(n_1636),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1593),
.B(n_1109),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1496),
.Y(n_1705)
);

BUFx2_ASAP7_75t_L g1706 ( 
.A(n_1592),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1539),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1499),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1532),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1472),
.A2(n_834),
.B1(n_835),
.B2(n_833),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_1594),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1620),
.A2(n_837),
.B1(n_842),
.B2(n_835),
.C(n_834),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_SL g1713 ( 
.A(n_1566),
.B(n_1568),
.Y(n_1713)
);

INVx4_ASAP7_75t_L g1714 ( 
.A(n_1453),
.Y(n_1714)
);

INVx4_ASAP7_75t_SL g1715 ( 
.A(n_1511),
.Y(n_1715)
);

INVx3_ASAP7_75t_L g1716 ( 
.A(n_1539),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1519),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1539),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1442),
.A2(n_1613),
.B1(n_1636),
.B2(n_1478),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1599),
.B(n_1109),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1554),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1581),
.B(n_1650),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1603),
.A2(n_853),
.B1(n_862),
.B2(n_850),
.Y(n_1724)
);

INVx4_ASAP7_75t_L g1725 ( 
.A(n_1627),
.Y(n_1725)
);

NAND2xp33_ASAP7_75t_L g1726 ( 
.A(n_1511),
.B(n_1109),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1609),
.B(n_1109),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1636),
.B(n_1581),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1554),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1569),
.B(n_889),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1584),
.B(n_837),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1614),
.B(n_1109),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1621),
.B(n_1029),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1651),
.B(n_864),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1619),
.B(n_1134),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1528),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1556),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1528),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1531),
.Y(n_1739)
);

INVx3_ASAP7_75t_L g1740 ( 
.A(n_1556),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1596),
.Y(n_1741)
);

INVx3_ASAP7_75t_L g1742 ( 
.A(n_1556),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1623),
.B(n_870),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1505),
.B(n_845),
.C(n_842),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1535),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1624),
.B(n_875),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1530),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1625),
.B(n_874),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1530),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1626),
.B(n_881),
.Y(n_1750)
);

CKINVDCx8_ASAP7_75t_R g1751 ( 
.A(n_1570),
.Y(n_1751)
);

INVx2_ASAP7_75t_SL g1752 ( 
.A(n_1462),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1521),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1521),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1559),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1548),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1630),
.B(n_882),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1526),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1547),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1574),
.B(n_890),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1559),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1633),
.B(n_1134),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1642),
.B(n_1134),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1575),
.B(n_892),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1533),
.B(n_1068),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1644),
.B(n_1134),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1540),
.Y(n_1767)
);

INVx1_ASAP7_75t_SL g1768 ( 
.A(n_1546),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1559),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1645),
.B(n_875),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1647),
.B(n_1590),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1462),
.B(n_898),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1595),
.B(n_893),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1437),
.Y(n_1774)
);

AND2x6_ASAP7_75t_L g1775 ( 
.A(n_1631),
.B(n_1142),
.Y(n_1775)
);

INVx2_ASAP7_75t_SL g1776 ( 
.A(n_1598),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1549),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1598),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1506),
.B(n_896),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1562),
.B(n_1134),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1547),
.Y(n_1781)
);

INVx5_ASAP7_75t_L g1782 ( 
.A(n_1511),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1463),
.A2(n_847),
.B1(n_849),
.B2(n_845),
.Y(n_1783)
);

INVx5_ASAP7_75t_L g1784 ( 
.A(n_1469),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1541),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1545),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1576),
.B(n_1099),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1576),
.B(n_899),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1550),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1467),
.B(n_900),
.Y(n_1790)
);

BUFx4f_ASAP7_75t_L g1791 ( 
.A(n_1582),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1608),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1631),
.B(n_1134),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1611),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1469),
.Y(n_1795)
);

INVx1_ASAP7_75t_SL g1796 ( 
.A(n_1551),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1524),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1612),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1618),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1622),
.B(n_902),
.Y(n_1800)
);

INVxp67_ASAP7_75t_SL g1801 ( 
.A(n_1481),
.Y(n_1801)
);

INVx3_ASAP7_75t_L g1802 ( 
.A(n_1629),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1638),
.Y(n_1803)
);

AND2x6_ASAP7_75t_L g1804 ( 
.A(n_1582),
.B(n_1142),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1622),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1522),
.B(n_1068),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1648),
.B(n_1099),
.Y(n_1807)
);

INVx3_ASAP7_75t_L g1808 ( 
.A(n_1643),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1536),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1543),
.Y(n_1810)
);

INVx3_ASAP7_75t_L g1811 ( 
.A(n_1646),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1544),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1469),
.Y(n_1813)
);

AND2x2_ASAP7_75t_SL g1814 ( 
.A(n_1597),
.B(n_1157),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1648),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1557),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1635),
.Y(n_1817)
);

CKINVDCx11_ASAP7_75t_R g1818 ( 
.A(n_1558),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1640),
.B(n_1068),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1649),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1468),
.B(n_1070),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1583),
.B(n_1474),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1606),
.Y(n_1823)
);

BUFx3_ASAP7_75t_L g1824 ( 
.A(n_1531),
.Y(n_1824)
);

INVx5_ASAP7_75t_L g1825 ( 
.A(n_1475),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1582),
.Y(n_1826)
);

OR2x6_ASAP7_75t_L g1827 ( 
.A(n_1586),
.B(n_1157),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1518),
.Y(n_1828)
);

BUFx4f_ASAP7_75t_L g1829 ( 
.A(n_1585),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1473),
.Y(n_1830)
);

BUFx3_ASAP7_75t_L g1831 ( 
.A(n_1563),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1482),
.B(n_1494),
.Y(n_1832)
);

INVx4_ASAP7_75t_L g1833 ( 
.A(n_1565),
.Y(n_1833)
);

CKINVDCx14_ASAP7_75t_R g1834 ( 
.A(n_1500),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1441),
.B(n_847),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1479),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1475),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1475),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1486),
.B(n_1491),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1585),
.Y(n_1840)
);

AND2x2_ASAP7_75t_SL g1841 ( 
.A(n_1587),
.B(n_1183),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1495),
.A2(n_1502),
.B1(n_1508),
.B2(n_1498),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1489),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1489),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1510),
.B(n_1070),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1489),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1460),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1514),
.Y(n_1848)
);

AND2x6_ASAP7_75t_L g1849 ( 
.A(n_1466),
.B(n_1183),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1516),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1439),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1520),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1527),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1529),
.A2(n_904),
.B1(n_906),
.B2(n_903),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1577),
.B(n_909),
.Y(n_1855)
);

NOR2xp33_ASAP7_75t_L g1856 ( 
.A(n_1579),
.B(n_905),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1470),
.Y(n_1857)
);

NAND3xp33_ASAP7_75t_L g1858 ( 
.A(n_1470),
.B(n_851),
.C(n_849),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1443),
.B(n_917),
.Y(n_1859)
);

BUFx6f_ASAP7_75t_L g1860 ( 
.A(n_1439),
.Y(n_1860)
);

INVx3_ASAP7_75t_L g1861 ( 
.A(n_1439),
.Y(n_1861)
);

BUFx10_ASAP7_75t_L g1862 ( 
.A(n_1641),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1444),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1444),
.A2(n_937),
.B1(n_938),
.B2(n_934),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1447),
.B(n_910),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1451),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1451),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1449),
.B(n_911),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1504),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1567),
.B(n_1134),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1451),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1454),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1454),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1454),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1457),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1457),
.Y(n_1876)
);

INVxp67_ASAP7_75t_SL g1877 ( 
.A(n_1476),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1457),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1605),
.Y(n_1879)
);

INVxp67_ASAP7_75t_SL g1880 ( 
.A(n_1492),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1456),
.B(n_1458),
.Y(n_1881)
);

AO22x2_ASAP7_75t_L g1882 ( 
.A1(n_1450),
.A2(n_985),
.B1(n_1074),
.B2(n_969),
.Y(n_1882)
);

BUFx2_ASAP7_75t_L g1883 ( 
.A(n_1588),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1602),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1604),
.B(n_913),
.Y(n_1886)
);

AND2x6_ASAP7_75t_L g1887 ( 
.A(n_1605),
.B(n_1276),
.Y(n_1887)
);

AND2x6_ASAP7_75t_L g1888 ( 
.A(n_1605),
.B(n_1276),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1607),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1616),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1639),
.B(n_1134),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1617),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1632),
.B(n_915),
.Y(n_1893)
);

INVx4_ASAP7_75t_SL g1894 ( 
.A(n_1488),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1634),
.B(n_1637),
.Y(n_1895)
);

INVxp67_ASAP7_75t_SL g1896 ( 
.A(n_1493),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1560),
.Y(n_1897)
);

BUFx4_ASAP7_75t_L g1898 ( 
.A(n_1561),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1571),
.B(n_947),
.Y(n_1899)
);

INVx5_ASAP7_75t_L g1900 ( 
.A(n_1572),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1573),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1507),
.Y(n_1902)
);

NAND3xp33_ASAP7_75t_L g1903 ( 
.A(n_1512),
.B(n_854),
.C(n_851),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1553),
.Y(n_1904)
);

OR2x6_ASAP7_75t_L g1905 ( 
.A(n_1537),
.B(n_1302),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1538),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1578),
.B(n_916),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1501),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1578),
.B(n_919),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1564),
.B(n_1229),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1501),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1501),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1513),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1501),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1501),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_1459),
.Y(n_1916)
);

INVx4_ASAP7_75t_L g1917 ( 
.A(n_1564),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1459),
.Y(n_1918)
);

AND2x6_ASAP7_75t_L g1919 ( 
.A(n_1578),
.B(n_1099),
.Y(n_1919)
);

INVx3_ASAP7_75t_L g1920 ( 
.A(n_1513),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1578),
.B(n_921),
.Y(n_1921)
);

INVx4_ASAP7_75t_L g1922 ( 
.A(n_1564),
.Y(n_1922)
);

BUFx4f_ASAP7_75t_L g1923 ( 
.A(n_1582),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1501),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1600),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1542),
.B(n_1070),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1503),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1542),
.B(n_1080),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1564),
.Y(n_1929)
);

BUFx10_ASAP7_75t_L g1930 ( 
.A(n_1483),
.Y(n_1930)
);

AND2x6_ASAP7_75t_L g1931 ( 
.A(n_1578),
.B(n_1099),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1503),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1503),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1578),
.B(n_922),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1436),
.B(n_1099),
.Y(n_1935)
);

BUFx6f_ASAP7_75t_L g1936 ( 
.A(n_1615),
.Y(n_1936)
);

INVx4_ASAP7_75t_L g1937 ( 
.A(n_1564),
.Y(n_1937)
);

AND2x6_ASAP7_75t_L g1938 ( 
.A(n_1578),
.B(n_1140),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1503),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1503),
.Y(n_1940)
);

NAND3x1_ASAP7_75t_L g1941 ( 
.A(n_1620),
.B(n_940),
.C(n_891),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1600),
.Y(n_1942)
);

OR2x6_ASAP7_75t_L g1943 ( 
.A(n_1824),
.B(n_949),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1917),
.B(n_854),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1688),
.B(n_855),
.Y(n_1945)
);

BUFx6f_ASAP7_75t_L g1946 ( 
.A(n_1689),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1917),
.B(n_855),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1756),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1922),
.B(n_1937),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1922),
.B(n_856),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1781),
.Y(n_1951)
);

AOI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1728),
.A2(n_1703),
.B1(n_1717),
.B2(n_1720),
.Y(n_1952)
);

INVxp67_ASAP7_75t_SL g1953 ( 
.A(n_1728),
.Y(n_1953)
);

O2A1O1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1723),
.A2(n_961),
.B(n_972),
.C(n_955),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1781),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1681),
.B(n_1294),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1671),
.B(n_856),
.Y(n_1957)
);

AOI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1703),
.A2(n_859),
.B1(n_863),
.B2(n_857),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_SL g1959 ( 
.A(n_1929),
.B(n_857),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1731),
.B(n_859),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1929),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1684),
.B(n_1300),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1676),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1685),
.B(n_1300),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1691),
.B(n_1301),
.Y(n_1965)
);

NOR3xp33_ASAP7_75t_L g1966 ( 
.A(n_1712),
.B(n_1100),
.C(n_1094),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1695),
.B(n_1280),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1696),
.Y(n_1968)
);

INVxp67_ASAP7_75t_SL g1969 ( 
.A(n_1709),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1697),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1937),
.B(n_863),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1687),
.A2(n_978),
.B(n_973),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1734),
.B(n_865),
.Y(n_1973)
);

INVx2_ASAP7_75t_SL g1974 ( 
.A(n_1930),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1820),
.B(n_865),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1734),
.B(n_867),
.Y(n_1976)
);

A2O1A1Ixp33_ASAP7_75t_L g1977 ( 
.A1(n_1702),
.A2(n_995),
.B(n_997),
.C(n_992),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1736),
.B(n_867),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1692),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1736),
.B(n_869),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1743),
.B(n_869),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1745),
.B(n_1291),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1743),
.B(n_871),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1748),
.B(n_1750),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1705),
.Y(n_1985)
);

AOI22xp33_ASAP7_75t_L g1986 ( 
.A1(n_1733),
.A2(n_1775),
.B1(n_1748),
.B2(n_1757),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1750),
.B(n_871),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1708),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1692),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1739),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1757),
.B(n_872),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1718),
.Y(n_1992)
);

A2O1A1Ixp33_ASAP7_75t_L g1993 ( 
.A1(n_1771),
.A2(n_1009),
.B(n_1026),
.C(n_1001),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1747),
.B(n_872),
.Y(n_1994)
);

INVx3_ASAP7_75t_L g1995 ( 
.A(n_1747),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1836),
.B(n_873),
.Y(n_1996)
);

INVx2_ASAP7_75t_SL g1997 ( 
.A(n_1930),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1675),
.B(n_873),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1699),
.A2(n_1028),
.B(n_1027),
.Y(n_1999)
);

BUFx6f_ASAP7_75t_L g2000 ( 
.A(n_1729),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1658),
.B(n_876),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1926),
.B(n_1928),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1775),
.A2(n_1039),
.B1(n_1041),
.B2(n_1037),
.Y(n_2003)
);

OAI22xp5_ASAP7_75t_L g2004 ( 
.A1(n_1655),
.A2(n_1060),
.B1(n_1064),
.B2(n_1053),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1768),
.B(n_876),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1777),
.B(n_878),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1669),
.B(n_878),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1775),
.A2(n_1085),
.B1(n_1086),
.B2(n_1067),
.Y(n_2008)
);

OAI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1655),
.A2(n_1097),
.B1(n_1106),
.B2(n_1089),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1753),
.Y(n_2010)
);

OAI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_1854),
.A2(n_1056),
.B1(n_1238),
.B2(n_880),
.C(n_879),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_SL g2012 ( 
.A(n_1862),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1775),
.A2(n_1107),
.B1(n_1111),
.B2(n_1108),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1657),
.A2(n_1116),
.B1(n_1117),
.B2(n_1115),
.Y(n_2014)
);

AOI22xp33_ASAP7_75t_L g2015 ( 
.A1(n_1652),
.A2(n_1120),
.B1(n_1127),
.B2(n_1126),
.Y(n_2015)
);

NOR2xp67_ASAP7_75t_SL g2016 ( 
.A(n_1782),
.B(n_1290),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1678),
.B(n_879),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1679),
.B(n_880),
.Y(n_2018)
);

NOR2xp33_ASAP7_75t_L g2019 ( 
.A(n_1661),
.B(n_1056),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1754),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1797),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1809),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_1801),
.Y(n_2023)
);

OR2x2_ASAP7_75t_SL g2024 ( 
.A(n_1863),
.B(n_998),
.Y(n_2024)
);

INVxp67_ASAP7_75t_L g2025 ( 
.A(n_1817),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1908),
.B(n_1238),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1789),
.B(n_1796),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1911),
.B(n_1239),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1810),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1912),
.B(n_1239),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1812),
.Y(n_2031)
);

HB1xp67_ASAP7_75t_L g2032 ( 
.A(n_1905),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1905),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1657),
.B(n_1301),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_L g2035 ( 
.A1(n_1907),
.A2(n_1130),
.B1(n_1138),
.B2(n_1137),
.Y(n_2035)
);

INVx4_ASAP7_75t_L g2036 ( 
.A(n_1833),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1729),
.Y(n_2037)
);

AOI22xp5_ASAP7_75t_L g2038 ( 
.A1(n_1668),
.A2(n_1244),
.B1(n_1245),
.B2(n_1240),
.Y(n_2038)
);

AND2x6_ASAP7_75t_SL g2039 ( 
.A(n_1881),
.B(n_1146),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1694),
.B(n_1240),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1927),
.B(n_1283),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1841),
.B(n_1244),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1914),
.B(n_1245),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_SL g2044 ( 
.A(n_1885),
.B(n_1248),
.C(n_1247),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1915),
.B(n_1247),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_SL g2046 ( 
.A(n_1833),
.B(n_1000),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1815),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1829),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1701),
.B(n_1248),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1924),
.B(n_1253),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1909),
.B(n_1253),
.Y(n_2051)
);

BUFx3_ASAP7_75t_L g2052 ( 
.A(n_1826),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1921),
.B(n_1261),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1934),
.B(n_1261),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1759),
.Y(n_2055)
);

AOI21xp5_ASAP7_75t_L g2056 ( 
.A1(n_1659),
.A2(n_1153),
.B(n_1150),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1822),
.A2(n_1266),
.B1(n_1268),
.B2(n_1265),
.Y(n_2057)
);

INVxp33_ASAP7_75t_L g2058 ( 
.A(n_1818),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1769),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1654),
.B(n_1265),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_1829),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1782),
.B(n_1814),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1831),
.A2(n_1007),
.B1(n_1019),
.B2(n_1004),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1785),
.B(n_1266),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1782),
.B(n_1268),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1785),
.B(n_1270),
.Y(n_2066)
);

BUFx3_ASAP7_75t_L g2067 ( 
.A(n_1791),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1758),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1663),
.B(n_1270),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1663),
.B(n_1273),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1673),
.B(n_1273),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1767),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1786),
.Y(n_2073)
);

NOR2xp33_ASAP7_75t_L g2074 ( 
.A(n_1765),
.B(n_1274),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1680),
.Y(n_2075)
);

AOI22xp5_ASAP7_75t_L g2076 ( 
.A1(n_1840),
.A2(n_1277),
.B1(n_1279),
.B2(n_1274),
.Y(n_2076)
);

NOR2xp67_ASAP7_75t_L g2077 ( 
.A(n_1858),
.B(n_4),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1682),
.B(n_1277),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1752),
.B(n_1279),
.Y(n_2079)
);

CKINVDCx5p33_ASAP7_75t_R g2080 ( 
.A(n_1711),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1713),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1776),
.B(n_1280),
.Y(n_2082)
);

CKINVDCx20_ASAP7_75t_R g2083 ( 
.A(n_1823),
.Y(n_2083)
);

INVx2_ASAP7_75t_SL g2084 ( 
.A(n_1791),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1848),
.B(n_1283),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1794),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1778),
.B(n_1285),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_SL g2088 ( 
.A(n_1744),
.B(n_1285),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1805),
.B(n_1290),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_1806),
.A2(n_1292),
.B1(n_1294),
.B2(n_1291),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1730),
.B(n_1292),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1802),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1760),
.B(n_923),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_1764),
.B(n_927),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1693),
.Y(n_2095)
);

OR2x6_ASAP7_75t_L g2096 ( 
.A(n_1857),
.B(n_1941),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_SL g2097 ( 
.A(n_1783),
.B(n_929),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1923),
.B(n_931),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1772),
.B(n_935),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_1819),
.A2(n_941),
.B1(n_942),
.B2(n_939),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1923),
.B(n_943),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1710),
.B(n_946),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1821),
.B(n_1020),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1772),
.B(n_1779),
.Y(n_2104)
);

AOI22xp33_ASAP7_75t_L g2105 ( 
.A1(n_1664),
.A2(n_1155),
.B1(n_1159),
.B2(n_1158),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1656),
.B(n_1800),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1802),
.Y(n_2107)
);

AOI21xp5_ASAP7_75t_L g2108 ( 
.A1(n_1659),
.A2(n_1173),
.B(n_1171),
.Y(n_2108)
);

INVx2_ASAP7_75t_SL g2109 ( 
.A(n_1827),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1870),
.B(n_948),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1724),
.B(n_1773),
.Y(n_2111)
);

AOI22xp5_ASAP7_75t_L g2112 ( 
.A1(n_1662),
.A2(n_951),
.B1(n_953),
.B2(n_950),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1704),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1738),
.B(n_954),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1900),
.Y(n_2115)
);

CKINVDCx5p33_ASAP7_75t_R g2116 ( 
.A(n_1916),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1850),
.B(n_956),
.Y(n_2117)
);

BUFx6f_ASAP7_75t_L g2118 ( 
.A(n_1936),
.Y(n_2118)
);

O2A1O1Ixp33_ASAP7_75t_L g2119 ( 
.A1(n_1721),
.A2(n_1174),
.B(n_1177),
.C(n_1176),
.Y(n_2119)
);

A2O1A1Ixp33_ASAP7_75t_L g2120 ( 
.A1(n_1793),
.A2(n_1180),
.B(n_1192),
.C(n_1187),
.Y(n_2120)
);

NOR2xp33_ASAP7_75t_L g2121 ( 
.A(n_1845),
.B(n_1031),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1727),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1852),
.B(n_1853),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_SL g2124 ( 
.A(n_1674),
.B(n_957),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_SL g2125 ( 
.A(n_1666),
.B(n_958),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_1714),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1732),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1735),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1666),
.B(n_959),
.Y(n_2129)
);

OR2x2_ASAP7_75t_L g2130 ( 
.A(n_1835),
.B(n_1104),
.Y(n_2130)
);

OR2x6_ASAP7_75t_SL g2131 ( 
.A(n_1918),
.B(n_1842),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_1927),
.A2(n_1196),
.B1(n_1198),
.B2(n_1193),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1808),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_1859),
.B(n_1080),
.Y(n_2134)
);

AOI22xp33_ASAP7_75t_L g2135 ( 
.A1(n_1849),
.A2(n_1207),
.B1(n_1211),
.B2(n_1201),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_1834),
.Y(n_2136)
);

NAND2xp33_ASAP7_75t_L g2137 ( 
.A(n_1932),
.B(n_1229),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1762),
.Y(n_2138)
);

INVx5_ASAP7_75t_L g2139 ( 
.A(n_1919),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1763),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_L g2141 ( 
.A1(n_1932),
.A2(n_1230),
.B(n_1237),
.C(n_1227),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1808),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_L g2143 ( 
.A1(n_1849),
.A2(n_1246),
.B1(n_1258),
.B2(n_1254),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1766),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1749),
.B(n_962),
.Y(n_2145)
);

BUFx3_ASAP7_75t_L g2146 ( 
.A(n_1900),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1790),
.B(n_963),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1788),
.B(n_965),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_SL g2149 ( 
.A(n_1933),
.B(n_1032),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1666),
.B(n_967),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_1811),
.Y(n_2151)
);

AOI22xp5_ASAP7_75t_L g2152 ( 
.A1(n_1828),
.A2(n_971),
.B1(n_974),
.B2(n_968),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_SL g2153 ( 
.A(n_1741),
.B(n_975),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1891),
.B(n_976),
.Y(n_2154)
);

BUFx3_ASAP7_75t_L g2155 ( 
.A(n_1900),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1933),
.B(n_1939),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1939),
.B(n_977),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1940),
.B(n_980),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1940),
.B(n_981),
.Y(n_2159)
);

AOI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1849),
.A2(n_1263),
.B1(n_1267),
.B2(n_1264),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1856),
.A2(n_983),
.B1(n_984),
.B2(n_982),
.Y(n_2161)
);

INVx2_ASAP7_75t_L g2162 ( 
.A(n_1811),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1780),
.B(n_986),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1859),
.B(n_1080),
.Y(n_2164)
);

O2A1O1Ixp5_ASAP7_75t_L g2165 ( 
.A1(n_1935),
.A2(n_1269),
.B(n_1282),
.C(n_1281),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1830),
.B(n_988),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1936),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1816),
.B(n_989),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_1910),
.B(n_993),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_1889),
.B(n_1093),
.Y(n_2170)
);

OR2x2_ASAP7_75t_L g2171 ( 
.A(n_1883),
.B(n_1260),
.Y(n_2171)
);

AND2x6_ASAP7_75t_L g2172 ( 
.A(n_1936),
.B(n_1140),
.Y(n_2172)
);

INVx4_ASAP7_75t_L g2173 ( 
.A(n_1804),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1890),
.B(n_1125),
.Y(n_2174)
);

NOR3x1_ASAP7_75t_L g2175 ( 
.A(n_1877),
.B(n_1242),
.C(n_1163),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1807),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1832),
.B(n_994),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1660),
.Y(n_2178)
);

INVx8_ASAP7_75t_L g2179 ( 
.A(n_1827),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1774),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1665),
.B(n_1925),
.Y(n_2181)
);

AOI22xp33_ASAP7_75t_L g2182 ( 
.A1(n_1849),
.A2(n_1284),
.B1(n_1287),
.B2(n_1286),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1670),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1672),
.B(n_996),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1942),
.B(n_1002),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1706),
.B(n_1003),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_1847),
.A2(n_1298),
.B(n_1010),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_L g2188 ( 
.A(n_1714),
.B(n_1005),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_1869),
.B(n_1012),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_SL g2190 ( 
.A(n_1725),
.B(n_1013),
.Y(n_2190)
);

CKINVDCx5p33_ASAP7_75t_R g2191 ( 
.A(n_1751),
.Y(n_2191)
);

CKINVDCx5p33_ASAP7_75t_R g2192 ( 
.A(n_1862),
.Y(n_2192)
);

AND2x4_ASAP7_75t_L g2193 ( 
.A(n_1725),
.B(n_1256),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_1892),
.B(n_1014),
.Y(n_2194)
);

OR2x6_ASAP7_75t_L g2195 ( 
.A(n_1839),
.B(n_1140),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1792),
.B(n_1798),
.Y(n_2196)
);

NOR2x1p5_ASAP7_75t_L g2197 ( 
.A(n_1880),
.B(n_1022),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1799),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_SL g2199 ( 
.A(n_1864),
.B(n_1015),
.Y(n_2199)
);

AND2x6_ASAP7_75t_SL g2200 ( 
.A(n_1884),
.B(n_1178),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_1855),
.B(n_1178),
.Y(n_2201)
);

OR2x6_ASAP7_75t_L g2202 ( 
.A(n_1855),
.B(n_1140),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_1865),
.A2(n_1017),
.B1(n_1018),
.B2(n_1016),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_1715),
.B(n_1903),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1803),
.B(n_1023),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1804),
.B(n_1024),
.Y(n_2206)
);

O2A1O1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_1690),
.A2(n_1278),
.B(n_1275),
.C(n_1178),
.Y(n_2207)
);

AND2x2_ASAP7_75t_L g2208 ( 
.A(n_1868),
.B(n_1275),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1886),
.B(n_1275),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_SL g2210 ( 
.A(n_1715),
.B(n_1025),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_1804),
.B(n_1030),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1746),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1653),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1804),
.Y(n_2214)
);

NOR2xp33_ASAP7_75t_L g2215 ( 
.A(n_1893),
.B(n_1033),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1653),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_1667),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_SL g2218 ( 
.A(n_1919),
.B(n_1295),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_1770),
.B(n_1034),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_SL g2220 ( 
.A(n_1784),
.B(n_1035),
.Y(n_2220)
);

NAND2xp5_ASAP7_75t_L g2221 ( 
.A(n_1784),
.B(n_1036),
.Y(n_2221)
);

OAI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_1896),
.A2(n_1236),
.B1(n_1235),
.B2(n_1040),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1667),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_SL g2224 ( 
.A(n_1784),
.B(n_1038),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_1899),
.A2(n_1726),
.B1(n_1677),
.B2(n_1895),
.Y(n_2225)
);

INVxp33_ASAP7_75t_L g2226 ( 
.A(n_1902),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_1898),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1825),
.B(n_1043),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_1825),
.B(n_1044),
.Y(n_2229)
);

AOI22xp5_ASAP7_75t_L g2230 ( 
.A1(n_1899),
.A2(n_1047),
.B1(n_1048),
.B2(n_1046),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1825),
.B(n_1049),
.Y(n_2231)
);

NOR2x1p5_ASAP7_75t_L g2232 ( 
.A(n_1897),
.B(n_1221),
.Y(n_2232)
);

INVxp67_ASAP7_75t_L g2233 ( 
.A(n_1904),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_1698),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_L g2235 ( 
.A(n_1698),
.B(n_1050),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_SL g2236 ( 
.A(n_1716),
.B(n_1051),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_1882),
.B(n_1295),
.Y(n_2237)
);

BUFx3_ASAP7_75t_L g2238 ( 
.A(n_1901),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_1716),
.B(n_1719),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_1719),
.B(n_1052),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1787),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_1722),
.B(n_1058),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_SL g2243 ( 
.A(n_1737),
.B(n_1059),
.Y(n_2243)
);

AOI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_1843),
.A2(n_1062),
.B(n_1061),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_SL g2245 ( 
.A(n_1919),
.B(n_1931),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_1938),
.A2(n_1229),
.B1(n_1295),
.B2(n_1191),
.Y(n_2246)
);

NAND2x1p5_ASAP7_75t_L g2247 ( 
.A(n_1740),
.B(n_1140),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_1882),
.A2(n_1742),
.B1(n_1755),
.B2(n_1740),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_SL g2249 ( 
.A(n_1742),
.B(n_1066),
.Y(n_2249)
);

BUFx3_ASAP7_75t_L g2250 ( 
.A(n_1906),
.Y(n_2250)
);

AOI21xp5_ASAP7_75t_L g2251 ( 
.A1(n_1844),
.A2(n_1071),
.B(n_1069),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1700),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1755),
.B(n_1072),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1913),
.B(n_1920),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1913),
.B(n_1073),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1920),
.B(n_1076),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_1683),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1686),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_1938),
.A2(n_1229),
.B1(n_1255),
.B2(n_1191),
.Y(n_2259)
);

AND2x6_ASAP7_75t_SL g2260 ( 
.A(n_1894),
.B(n_5),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_SL g2261 ( 
.A(n_1795),
.B(n_1077),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1938),
.B(n_1078),
.Y(n_2262)
);

CKINVDCx5p33_ASAP7_75t_R g2263 ( 
.A(n_1894),
.Y(n_2263)
);

BUFx8_ASAP7_75t_L g2264 ( 
.A(n_1919),
.Y(n_2264)
);

INVxp67_ASAP7_75t_L g2265 ( 
.A(n_1931),
.Y(n_2265)
);

OAI22x1_ASAP7_75t_L g2266 ( 
.A1(n_1931),
.A2(n_1081),
.B1(n_1084),
.B2(n_1079),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_1707),
.B(n_1087),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_1931),
.B(n_1091),
.Y(n_2268)
);

AOI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_1938),
.A2(n_1095),
.B1(n_1096),
.B2(n_1092),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1761),
.Y(n_2270)
);

BUFx6f_ASAP7_75t_L g2271 ( 
.A(n_1795),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1887),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_1948),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1968),
.Y(n_2274)
);

INVxp67_ASAP7_75t_SL g2275 ( 
.A(n_2156),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1970),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1963),
.B(n_1837),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1985),
.B(n_1838),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_1988),
.B(n_1846),
.Y(n_2279)
);

NOR2xp33_ASAP7_75t_R g2280 ( 
.A(n_2046),
.B(n_1101),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_2149),
.B(n_1813),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2027),
.B(n_1103),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1992),
.Y(n_2283)
);

BUFx3_ASAP7_75t_L g2284 ( 
.A(n_2083),
.Y(n_2284)
);

INVx1_ASAP7_75t_SL g2285 ( 
.A(n_2156),
.Y(n_2285)
);

BUFx4f_ASAP7_75t_L g2286 ( 
.A(n_2179),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1955),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2021),
.B(n_2022),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2029),
.Y(n_2289)
);

AOI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2149),
.A2(n_1110),
.B1(n_1112),
.B2(n_1105),
.Y(n_2290)
);

BUFx3_ASAP7_75t_L g2291 ( 
.A(n_1990),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2202),
.Y(n_2292)
);

OR2x6_ASAP7_75t_L g2293 ( 
.A(n_2179),
.B(n_2227),
.Y(n_2293)
);

AOI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2046),
.A2(n_1118),
.B1(n_1121),
.B2(n_1114),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_1957),
.A2(n_1123),
.B1(n_1124),
.B2(n_1122),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2031),
.B(n_1795),
.Y(n_2296)
);

INVx5_ASAP7_75t_L g2297 ( 
.A(n_2172),
.Y(n_2297)
);

NOR2xp33_ASAP7_75t_L g2298 ( 
.A(n_2103),
.B(n_1128),
.Y(n_2298)
);

BUFx3_ASAP7_75t_L g2299 ( 
.A(n_2179),
.Y(n_2299)
);

BUFx3_ASAP7_75t_L g2300 ( 
.A(n_2115),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2111),
.B(n_1813),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2095),
.B(n_1813),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_SL g2303 ( 
.A(n_2245),
.B(n_1887),
.Y(n_2303)
);

NAND2xp5_ASAP7_75t_L g2304 ( 
.A(n_2113),
.B(n_1229),
.Y(n_2304)
);

CKINVDCx5p33_ASAP7_75t_R g2305 ( 
.A(n_2012),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2122),
.B(n_1229),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_2271),
.Y(n_2307)
);

INVx3_ASAP7_75t_SL g2308 ( 
.A(n_2192),
.Y(n_2308)
);

NAND2xp5_ASAP7_75t_L g2309 ( 
.A(n_2127),
.B(n_1229),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2036),
.B(n_1887),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1984),
.Y(n_2311)
);

INVx6_ASAP7_75t_L g2312 ( 
.A(n_2036),
.Y(n_2312)
);

BUFx6f_ASAP7_75t_L g2313 ( 
.A(n_2271),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_2023),
.B(n_1129),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2075),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_2055),
.Y(n_2316)
);

NAND2xp33_ASAP7_75t_R g2317 ( 
.A(n_2080),
.B(n_5),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2068),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_1955),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2072),
.Y(n_2320)
);

BUFx3_ASAP7_75t_L g2321 ( 
.A(n_2146),
.Y(n_2321)
);

HB1xp67_ASAP7_75t_L g2322 ( 
.A(n_2202),
.Y(n_2322)
);

AND2x2_ASAP7_75t_SL g2323 ( 
.A(n_2173),
.B(n_1191),
.Y(n_2323)
);

INVx1_ASAP7_75t_SL g2324 ( 
.A(n_2202),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2128),
.B(n_1229),
.Y(n_2325)
);

OAI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2063),
.A2(n_1132),
.B1(n_1133),
.B2(n_1131),
.Y(n_2326)
);

BUFx2_ASAP7_75t_SL g2327 ( 
.A(n_2012),
.Y(n_2327)
);

AND2x4_ASAP7_75t_L g2328 ( 
.A(n_2061),
.B(n_1887),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_1952),
.A2(n_1255),
.B1(n_1191),
.B2(n_1136),
.Y(n_2329)
);

INVxp67_ASAP7_75t_SL g2330 ( 
.A(n_1953),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2138),
.B(n_1135),
.Y(n_2331)
);

BUFx6f_ASAP7_75t_L g2332 ( 
.A(n_2271),
.Y(n_2332)
);

AO21x1_ASAP7_75t_L g2333 ( 
.A1(n_2248),
.A2(n_1874),
.B(n_1871),
.Y(n_2333)
);

AND3x1_ASAP7_75t_SL g2334 ( 
.A(n_2197),
.B(n_1141),
.C(n_1139),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2140),
.B(n_2144),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2073),
.Y(n_2336)
);

BUFx2_ASAP7_75t_L g2337 ( 
.A(n_1943),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2180),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2025),
.B(n_1143),
.Y(n_2339)
);

NOR3xp33_ASAP7_75t_SL g2340 ( 
.A(n_2136),
.B(n_1145),
.C(n_1144),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_1943),
.A2(n_1148),
.B1(n_1149),
.B2(n_1147),
.Y(n_2341)
);

INVx3_ASAP7_75t_L g2342 ( 
.A(n_1961),
.Y(n_2342)
);

NOR3xp33_ASAP7_75t_SL g2343 ( 
.A(n_2263),
.B(n_2191),
.C(n_2116),
.Y(n_2343)
);

OR2x6_ASAP7_75t_L g2344 ( 
.A(n_1943),
.B(n_1191),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_R g2345 ( 
.A(n_2264),
.B(n_1151),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2010),
.Y(n_2346)
);

INVxp67_ASAP7_75t_L g2347 ( 
.A(n_1969),
.Y(n_2347)
);

OR2x6_ASAP7_75t_L g2348 ( 
.A(n_2096),
.B(n_1255),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2020),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2034),
.B(n_1152),
.Y(n_2350)
);

AND2x4_ASAP7_75t_L g2351 ( 
.A(n_1974),
.B(n_1888),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2034),
.B(n_1154),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2041),
.B(n_2106),
.Y(n_2353)
);

INVx3_ASAP7_75t_L g2354 ( 
.A(n_1961),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_1996),
.B(n_1156),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2198),
.Y(n_2356)
);

NAND3xp33_ASAP7_75t_SL g2357 ( 
.A(n_2225),
.B(n_1161),
.C(n_1160),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2041),
.B(n_1162),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2178),
.Y(n_2359)
);

BUFx2_ASAP7_75t_L g2360 ( 
.A(n_2193),
.Y(n_2360)
);

AND2x2_ASAP7_75t_L g2361 ( 
.A(n_2005),
.B(n_1164),
.Y(n_2361)
);

INVx3_ASAP7_75t_L g2362 ( 
.A(n_1995),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2006),
.B(n_1167),
.Y(n_2363)
);

BUFx4f_ASAP7_75t_L g2364 ( 
.A(n_2195),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_1960),
.B(n_1168),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_1998),
.B(n_1169),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2183),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1986),
.B(n_1170),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2157),
.B(n_1175),
.Y(n_2369)
);

BUFx3_ASAP7_75t_L g2370 ( 
.A(n_2155),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2200),
.Y(n_2371)
);

AOI21xp5_ASAP7_75t_L g2372 ( 
.A1(n_2137),
.A2(n_1878),
.B(n_1876),
.Y(n_2372)
);

BUFx2_ASAP7_75t_L g2373 ( 
.A(n_2193),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_2157),
.B(n_1179),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2047),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_1997),
.B(n_1888),
.Y(n_2376)
);

NOR3xp33_ASAP7_75t_SL g2377 ( 
.A(n_2248),
.B(n_1185),
.C(n_1182),
.Y(n_2377)
);

OR2x6_ASAP7_75t_L g2378 ( 
.A(n_2096),
.B(n_1255),
.Y(n_2378)
);

NAND2xp5_ASAP7_75t_L g2379 ( 
.A(n_2158),
.B(n_1189),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2204),
.B(n_1888),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2002),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_2032),
.Y(n_2382)
);

BUFx3_ASAP7_75t_L g2383 ( 
.A(n_2052),
.Y(n_2383)
);

NOR3xp33_ASAP7_75t_SL g2384 ( 
.A(n_2121),
.B(n_1195),
.C(n_1194),
.Y(n_2384)
);

AO22x1_ASAP7_75t_L g2385 ( 
.A1(n_2058),
.A2(n_1888),
.B1(n_1200),
.B2(n_1202),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_L g2386 ( 
.A(n_2033),
.B(n_1199),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2181),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_2109),
.Y(n_2388)
);

HB1xp67_ASAP7_75t_L g2389 ( 
.A(n_1982),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2081),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_2181),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2196),
.Y(n_2392)
);

BUFx10_ASAP7_75t_L g2393 ( 
.A(n_2195),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2064),
.Y(n_2394)
);

BUFx10_ASAP7_75t_L g2395 ( 
.A(n_2195),
.Y(n_2395)
);

NOR2x1_ASAP7_75t_L g2396 ( 
.A(n_2096),
.B(n_1255),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2057),
.B(n_1203),
.Y(n_2397)
);

OR2x2_ASAP7_75t_L g2398 ( 
.A(n_2130),
.B(n_1204),
.Y(n_2398)
);

OR2x6_ASAP7_75t_L g2399 ( 
.A(n_2173),
.B(n_1851),
.Y(n_2399)
);

INVx4_ASAP7_75t_L g2400 ( 
.A(n_2067),
.Y(n_2400)
);

CKINVDCx6p67_ASAP7_75t_R g2401 ( 
.A(n_2238),
.Y(n_2401)
);

NAND2xp33_ASAP7_75t_SL g2402 ( 
.A(n_2016),
.B(n_1206),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_2222),
.B(n_1208),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2085),
.B(n_1212),
.Y(n_2404)
);

OR2x6_ASAP7_75t_L g2405 ( 
.A(n_2048),
.B(n_1851),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2066),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2038),
.B(n_1213),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_1946),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1956),
.Y(n_2409)
);

OR2x6_ASAP7_75t_L g2410 ( 
.A(n_2084),
.B(n_1851),
.Y(n_2410)
);

BUFx3_ASAP7_75t_L g2411 ( 
.A(n_2250),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2247),
.Y(n_2412)
);

AOI221xp5_ASAP7_75t_SL g2413 ( 
.A1(n_2141),
.A2(n_1879),
.B1(n_1867),
.B2(n_1860),
.C(n_1872),
.Y(n_2413)
);

INVx3_ASAP7_75t_L g2414 ( 
.A(n_1995),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2158),
.B(n_1216),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2237),
.B(n_1217),
.Y(n_2416)
);

INVxp67_ASAP7_75t_L g2417 ( 
.A(n_2171),
.Y(n_2417)
);

INVx5_ASAP7_75t_L g2418 ( 
.A(n_2172),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_1966),
.A2(n_1219),
.B1(n_1220),
.B2(n_1218),
.Y(n_2419)
);

AND2x4_ASAP7_75t_L g2420 ( 
.A(n_2204),
.B(n_5),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_1945),
.B(n_1222),
.Y(n_2421)
);

OR2x6_ASAP7_75t_L g2422 ( 
.A(n_2214),
.B(n_1860),
.Y(n_2422)
);

AOI22xp5_ASAP7_75t_SL g2423 ( 
.A1(n_2170),
.A2(n_1224),
.B1(n_1226),
.B2(n_1223),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2159),
.B(n_1231),
.Y(n_2424)
);

BUFx8_ASAP7_75t_SL g2425 ( 
.A(n_2134),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2159),
.B(n_1233),
.Y(n_2426)
);

OAI22xp5_ASAP7_75t_SL g2427 ( 
.A1(n_2024),
.A2(n_2174),
.B1(n_2011),
.B2(n_2230),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_2074),
.A2(n_1861),
.B1(n_1867),
.B2(n_1860),
.Y(n_2428)
);

A2O1A1Ixp33_ASAP7_75t_L g2429 ( 
.A1(n_2119),
.A2(n_1861),
.B(n_1873),
.C(n_1866),
.Y(n_2429)
);

INVxp67_ASAP7_75t_L g2430 ( 
.A(n_1950),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_2126),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_SL g2432 ( 
.A(n_2269),
.B(n_1867),
.Y(n_2432)
);

BUFx2_ASAP7_75t_L g2433 ( 
.A(n_2264),
.Y(n_2433)
);

AND2x6_ASAP7_75t_L g2434 ( 
.A(n_1951),
.B(n_1875),
.Y(n_2434)
);

AND2x6_ASAP7_75t_SL g2435 ( 
.A(n_2175),
.B(n_6),
.Y(n_2435)
);

NAND2xp33_ASAP7_75t_SL g2436 ( 
.A(n_2104),
.B(n_6),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_1956),
.Y(n_2437)
);

AOI211xp5_ASAP7_75t_L g2438 ( 
.A1(n_2207),
.A2(n_9),
.B(n_6),
.C(n_7),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2247),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_SL g2440 ( 
.A1(n_2131),
.A2(n_10),
.B1(n_7),
.B2(n_9),
.Y(n_2440)
);

BUFx2_ASAP7_75t_L g2441 ( 
.A(n_2039),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2123),
.B(n_9),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_1962),
.Y(n_2443)
);

INVx2_ASAP7_75t_L g2444 ( 
.A(n_2176),
.Y(n_2444)
);

AOI21xp5_ASAP7_75t_L g2445 ( 
.A1(n_2056),
.A2(n_10),
.B(n_11),
.Y(n_2445)
);

AND2x4_ASAP7_75t_L g2446 ( 
.A(n_2190),
.B(n_10),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_1958),
.B(n_12),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_1962),
.B(n_11),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_1964),
.B(n_11),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_1964),
.B(n_12),
.Y(n_2450)
);

INVx2_ASAP7_75t_SL g2451 ( 
.A(n_2232),
.Y(n_2451)
);

AND2x6_ASAP7_75t_SL g2452 ( 
.A(n_2164),
.B(n_12),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1965),
.Y(n_2453)
);

BUFx4f_ASAP7_75t_SL g2454 ( 
.A(n_2071),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_1965),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_2126),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1967),
.Y(n_2457)
);

BUFx12f_ASAP7_75t_L g2458 ( 
.A(n_2260),
.Y(n_2458)
);

BUFx8_ASAP7_75t_L g2459 ( 
.A(n_2201),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_1967),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_1993),
.B(n_2108),
.Y(n_2461)
);

HB1xp67_ASAP7_75t_L g2462 ( 
.A(n_2266),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_1954),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_2463)
);

BUFx12f_ASAP7_75t_L g2464 ( 
.A(n_2208),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_R g2465 ( 
.A(n_2218),
.B(n_13),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2086),
.Y(n_2466)
);

AO22x1_ASAP7_75t_L g2467 ( 
.A1(n_2139),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2120),
.B(n_15),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2007),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_SL g2470 ( 
.A(n_1973),
.B(n_16),
.Y(n_2470)
);

INVx4_ASAP7_75t_L g2471 ( 
.A(n_2139),
.Y(n_2471)
);

BUFx8_ASAP7_75t_L g2472 ( 
.A(n_2209),
.Y(n_2472)
);

BUFx3_ASAP7_75t_L g2473 ( 
.A(n_2092),
.Y(n_2473)
);

INVx5_ASAP7_75t_L g2474 ( 
.A(n_2172),
.Y(n_2474)
);

BUFx3_ASAP7_75t_L g2475 ( 
.A(n_2107),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2168),
.B(n_15),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2040),
.B(n_16),
.Y(n_2477)
);

BUFx4f_ASAP7_75t_L g2478 ( 
.A(n_2172),
.Y(n_2478)
);

BUFx3_ASAP7_75t_L g2479 ( 
.A(n_2133),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2004),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2142),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2062),
.B(n_17),
.Y(n_2482)
);

AND2x4_ASAP7_75t_L g2483 ( 
.A(n_2184),
.B(n_18),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2017),
.Y(n_2484)
);

OAI221xp5_ASAP7_75t_L g2485 ( 
.A1(n_2015),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.C(n_24),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_2168),
.B(n_20),
.Y(n_2486)
);

BUFx6f_ASAP7_75t_L g2487 ( 
.A(n_2000),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2018),
.Y(n_2488)
);

AND2x4_ASAP7_75t_L g2489 ( 
.A(n_2184),
.B(n_20),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_2035),
.B(n_21),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_L g2491 ( 
.A(n_2166),
.B(n_21),
.Y(n_2491)
);

BUFx12f_ASAP7_75t_L g2492 ( 
.A(n_2139),
.Y(n_2492)
);

OAI22xp5_ASAP7_75t_L g2493 ( 
.A1(n_2004),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2151),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2026),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2162),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_2000),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2000),
.Y(n_2498)
);

NOR2xp67_ASAP7_75t_L g2499 ( 
.A(n_2112),
.B(n_25),
.Y(n_2499)
);

BUFx2_ASAP7_75t_L g2500 ( 
.A(n_2221),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2028),
.Y(n_2501)
);

NAND2xp33_ASAP7_75t_SL g2502 ( 
.A(n_2044),
.B(n_25),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_R g2503 ( 
.A(n_2218),
.B(n_26),
.Y(n_2503)
);

AO22x1_ASAP7_75t_L g2504 ( 
.A1(n_2139),
.A2(n_29),
.B1(n_30),
.B2(n_28),
.Y(n_2504)
);

BUFx2_ASAP7_75t_L g2505 ( 
.A(n_2228),
.Y(n_2505)
);

CKINVDCx5p33_ASAP7_75t_R g2506 ( 
.A(n_2078),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2257),
.Y(n_2507)
);

OAI22xp5_ASAP7_75t_L g2508 ( 
.A1(n_2009),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2508)
);

NOR3xp33_ASAP7_75t_SL g2509 ( 
.A(n_1977),
.B(n_29),
.C(n_30),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2166),
.B(n_31),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_1999),
.B(n_31),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2030),
.Y(n_2512)
);

AOI211xp5_ASAP7_75t_L g2513 ( 
.A1(n_2049),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_2513)
);

HB1xp67_ASAP7_75t_L g2514 ( 
.A(n_2233),
.Y(n_2514)
);

CKINVDCx5p33_ASAP7_75t_R g2515 ( 
.A(n_2090),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_SL g2516 ( 
.A(n_1976),
.B(n_33),
.Y(n_2516)
);

INVx4_ASAP7_75t_L g2517 ( 
.A(n_2118),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_1972),
.B(n_32),
.Y(n_2518)
);

OR2x2_ASAP7_75t_L g2519 ( 
.A(n_1981),
.B(n_32),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_1975),
.B(n_33),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2185),
.B(n_34),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2043),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2045),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2258),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2050),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2118),
.Y(n_2526)
);

NOR3xp33_ASAP7_75t_SL g2527 ( 
.A(n_2199),
.B(n_34),
.C(n_36),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2118),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2177),
.B(n_36),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_1983),
.B(n_38),
.Y(n_2530)
);

HB1xp67_ASAP7_75t_L g2531 ( 
.A(n_2069),
.Y(n_2531)
);

INVx3_ASAP7_75t_L g2532 ( 
.A(n_2223),
.Y(n_2532)
);

BUFx3_ASAP7_75t_L g2533 ( 
.A(n_2229),
.Y(n_2533)
);

NOR3xp33_ASAP7_75t_SL g2534 ( 
.A(n_2215),
.B(n_37),
.C(n_38),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_2177),
.B(n_37),
.Y(n_2535)
);

NOR3xp33_ASAP7_75t_SL g2536 ( 
.A(n_2097),
.B(n_39),
.C(n_40),
.Y(n_2536)
);

BUFx4f_ASAP7_75t_L g2537 ( 
.A(n_2272),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2185),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_SL g2539 ( 
.A(n_1987),
.B(n_40),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2009),
.B(n_39),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2014),
.Y(n_2541)
);

INVx5_ASAP7_75t_L g2542 ( 
.A(n_2167),
.Y(n_2542)
);

HB1xp67_ASAP7_75t_L g2543 ( 
.A(n_2070),
.Y(n_2543)
);

HB1xp67_ASAP7_75t_L g2544 ( 
.A(n_1944),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2014),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2132),
.B(n_39),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2132),
.Y(n_2547)
);

INVx2_ASAP7_75t_L g2548 ( 
.A(n_2270),
.Y(n_2548)
);

BUFx3_ASAP7_75t_L g2549 ( 
.A(n_2231),
.Y(n_2549)
);

INVx4_ASAP7_75t_L g2550 ( 
.A(n_2167),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_1979),
.Y(n_2551)
);

NAND2xp5_ASAP7_75t_L g2552 ( 
.A(n_2169),
.B(n_2163),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2235),
.Y(n_2553)
);

NOR3xp33_ASAP7_75t_SL g2554 ( 
.A(n_2042),
.B(n_2102),
.C(n_2088),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2169),
.B(n_41),
.Y(n_2555)
);

OR2x6_ASAP7_75t_L g2556 ( 
.A(n_2098),
.B(n_41),
.Y(n_2556)
);

NOR3xp33_ASAP7_75t_SL g2557 ( 
.A(n_2189),
.B(n_2210),
.C(n_2153),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2242),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_L g2559 ( 
.A(n_2163),
.B(n_41),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_2105),
.B(n_42),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2255),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2256),
.Y(n_2562)
);

AND2x4_ASAP7_75t_L g2563 ( 
.A(n_1947),
.B(n_42),
.Y(n_2563)
);

HB1xp67_ASAP7_75t_L g2564 ( 
.A(n_1959),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2003),
.B(n_43),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_2008),
.B(n_43),
.Y(n_2566)
);

BUFx6f_ASAP7_75t_L g2567 ( 
.A(n_2167),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2205),
.Y(n_2568)
);

BUFx4f_ASAP7_75t_L g2569 ( 
.A(n_2223),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2013),
.B(n_43),
.Y(n_2570)
);

INVx5_ASAP7_75t_L g2571 ( 
.A(n_1989),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_SL g2572 ( 
.A(n_1991),
.B(n_45),
.Y(n_2572)
);

AND2x4_ASAP7_75t_L g2573 ( 
.A(n_1971),
.B(n_44),
.Y(n_2573)
);

NAND2xp33_ASAP7_75t_SL g2574 ( 
.A(n_1949),
.B(n_44),
.Y(n_2574)
);

CKINVDCx5p33_ASAP7_75t_R g2575 ( 
.A(n_2100),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2079),
.Y(n_2576)
);

NAND2xp5_ASAP7_75t_L g2577 ( 
.A(n_2091),
.B(n_45),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2051),
.B(n_46),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2053),
.B(n_46),
.Y(n_2579)
);

AND2x6_ASAP7_75t_L g2580 ( 
.A(n_2241),
.B(n_46),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2082),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_1978),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2001),
.B(n_47),
.Y(n_2583)
);

INVx4_ASAP7_75t_L g2584 ( 
.A(n_2037),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2087),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2089),
.Y(n_2586)
);

BUFx2_ASAP7_75t_L g2587 ( 
.A(n_2206),
.Y(n_2587)
);

AOI22xp33_ASAP7_75t_L g2588 ( 
.A1(n_2226),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2211),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2076),
.B(n_47),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2019),
.B(n_48),
.Y(n_2591)
);

INVxp67_ASAP7_75t_SL g2592 ( 
.A(n_2245),
.Y(n_2592)
);

BUFx6f_ASAP7_75t_L g2593 ( 
.A(n_2059),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2054),
.B(n_48),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2114),
.Y(n_2595)
);

INVx3_ASAP7_75t_SL g2596 ( 
.A(n_2220),
.Y(n_2596)
);

BUFx3_ASAP7_75t_L g2597 ( 
.A(n_2188),
.Y(n_2597)
);

NOR3xp33_ASAP7_75t_SL g2598 ( 
.A(n_2186),
.B(n_49),
.C(n_50),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2145),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2219),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2219),
.Y(n_2601)
);

BUFx2_ASAP7_75t_L g2602 ( 
.A(n_2268),
.Y(n_2602)
);

AND2x6_ASAP7_75t_L g2603 ( 
.A(n_2212),
.B(n_50),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_1980),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_R g2605 ( 
.A(n_2268),
.B(n_50),
.Y(n_2605)
);

O2A1O1Ixp33_ASAP7_75t_L g2606 ( 
.A1(n_2060),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2187),
.B(n_51),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2093),
.B(n_52),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_1994),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2094),
.B(n_53),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2147),
.B(n_2154),
.Y(n_2611)
);

AND2x4_ASAP7_75t_L g2612 ( 
.A(n_2117),
.B(n_53),
.Y(n_2612)
);

BUFx3_ASAP7_75t_L g2613 ( 
.A(n_2213),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_2099),
.B(n_55),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2077),
.Y(n_2615)
);

INVx1_ASAP7_75t_SL g2616 ( 
.A(n_2262),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2161),
.B(n_54),
.Y(n_2617)
);

AND3x2_ASAP7_75t_SL g2618 ( 
.A(n_2216),
.B(n_62),
.C(n_54),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2236),
.Y(n_2619)
);

AND2x4_ASAP7_75t_L g2620 ( 
.A(n_2125),
.B(n_54),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2240),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2243),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2249),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2253),
.Y(n_2624)
);

CKINVDCx5p33_ASAP7_75t_R g2625 ( 
.A(n_2152),
.Y(n_2625)
);

NAND2xp5_ASAP7_75t_L g2626 ( 
.A(n_2148),
.B(n_55),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2267),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2194),
.B(n_56),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2165),
.Y(n_2629)
);

BUFx6f_ASAP7_75t_L g2630 ( 
.A(n_2239),
.Y(n_2630)
);

AND2x2_ASAP7_75t_SL g2631 ( 
.A(n_2135),
.B(n_56),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2261),
.Y(n_2632)
);

INVx2_ASAP7_75t_L g2633 ( 
.A(n_2217),
.Y(n_2633)
);

INVx3_ASAP7_75t_L g2634 ( 
.A(n_2234),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2244),
.B(n_2251),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2203),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_R g2637 ( 
.A(n_2252),
.B(n_57),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2143),
.B(n_58),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2065),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2129),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2150),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2224),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2160),
.B(n_59),
.Y(n_2643)
);

OR2x6_ASAP7_75t_L g2644 ( 
.A(n_2101),
.B(n_59),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2182),
.B(n_60),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2254),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2110),
.B(n_2124),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_R g2648 ( 
.A(n_2246),
.B(n_60),
.Y(n_2648)
);

NOR2xp33_ASAP7_75t_L g2649 ( 
.A(n_2265),
.B(n_61),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2259),
.Y(n_2650)
);

AOI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2149),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_2651)
);

BUFx6f_ASAP7_75t_L g2652 ( 
.A(n_2271),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_1948),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_SL g2654 ( 
.A(n_2149),
.B(n_62),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_1948),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_1955),
.Y(n_2656)
);

INVx2_ASAP7_75t_L g2657 ( 
.A(n_2156),
.Y(n_2657)
);

INVx3_ASAP7_75t_L g2658 ( 
.A(n_1955),
.Y(n_2658)
);

BUFx6f_ASAP7_75t_L g2659 ( 
.A(n_2271),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2156),
.Y(n_2660)
);

NOR3xp33_ASAP7_75t_SL g2661 ( 
.A(n_2136),
.B(n_61),
.C(n_64),
.Y(n_2661)
);

AOI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_1966),
.A2(n_67),
.B1(n_64),
.B2(n_65),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_1948),
.Y(n_2663)
);

OR2x6_ASAP7_75t_L g2664 ( 
.A(n_2179),
.B(n_64),
.Y(n_2664)
);

AOI22xp5_ASAP7_75t_L g2665 ( 
.A1(n_2149),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_2665)
);

INVx4_ASAP7_75t_L g2666 ( 
.A(n_2179),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1948),
.Y(n_2667)
);

HB1xp67_ASAP7_75t_L g2668 ( 
.A(n_2027),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_1948),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_1948),
.Y(n_2670)
);

AOI22xp5_ASAP7_75t_SL g2671 ( 
.A1(n_2083),
.A2(n_67),
.B1(n_70),
.B2(n_69),
.Y(n_2671)
);

BUFx3_ASAP7_75t_L g2672 ( 
.A(n_2083),
.Y(n_2672)
);

NOR2xp67_ASAP7_75t_L g2673 ( 
.A(n_2227),
.B(n_70),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_1963),
.B(n_71),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_1948),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2156),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_1948),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_1963),
.B(n_71),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2027),
.B(n_72),
.Y(n_2679)
);

BUFx3_ASAP7_75t_L g2680 ( 
.A(n_2083),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2156),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_2179),
.Y(n_2682)
);

BUFx6f_ASAP7_75t_L g2683 ( 
.A(n_2271),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_1948),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_1963),
.B(n_72),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2149),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_1948),
.Y(n_2687)
);

BUFx2_ASAP7_75t_L g2688 ( 
.A(n_2027),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_1948),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2149),
.B(n_74),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_1963),
.B(n_75),
.Y(n_2691)
);

BUFx4f_ASAP7_75t_L g2692 ( 
.A(n_2179),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_1948),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_1948),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_L g2695 ( 
.A(n_2103),
.B(n_797),
.Y(n_2695)
);

INVx5_ASAP7_75t_L g2696 ( 
.A(n_2172),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_1948),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_1955),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2156),
.Y(n_2699)
);

BUFx6f_ASAP7_75t_L g2700 ( 
.A(n_2271),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_1966),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2156),
.Y(n_2702)
);

BUFx8_ASAP7_75t_L g2703 ( 
.A(n_2012),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2103),
.B(n_799),
.Y(n_2704)
);

AND2x4_ASAP7_75t_L g2705 ( 
.A(n_2036),
.B(n_77),
.Y(n_2705)
);

BUFx2_ASAP7_75t_L g2706 ( 
.A(n_2027),
.Y(n_2706)
);

BUFx3_ASAP7_75t_L g2707 ( 
.A(n_2083),
.Y(n_2707)
);

BUFx2_ASAP7_75t_L g2708 ( 
.A(n_2027),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_1948),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2027),
.Y(n_2710)
);

NOR2x1_ASAP7_75t_R g2711 ( 
.A(n_2036),
.B(n_78),
.Y(n_2711)
);

NOR3xp33_ASAP7_75t_SL g2712 ( 
.A(n_2136),
.B(n_80),
.C(n_81),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_1963),
.B(n_80),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_SL g2714 ( 
.A(n_2136),
.B(n_81),
.C(n_82),
.Y(n_2714)
);

CKINVDCx5p33_ASAP7_75t_R g2715 ( 
.A(n_2012),
.Y(n_2715)
);

AOI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2149),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2716)
);

AOI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2149),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_1948),
.Y(n_2718)
);

INVx3_ASAP7_75t_L g2719 ( 
.A(n_1955),
.Y(n_2719)
);

BUFx3_ASAP7_75t_L g2720 ( 
.A(n_2083),
.Y(n_2720)
);

OR2x2_ASAP7_75t_SL g2721 ( 
.A(n_2046),
.B(n_86),
.Y(n_2721)
);

INVx2_ASAP7_75t_SL g2722 ( 
.A(n_2179),
.Y(n_2722)
);

NOR3xp33_ASAP7_75t_SL g2723 ( 
.A(n_2136),
.B(n_87),
.C(n_89),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2027),
.B(n_89),
.Y(n_2724)
);

NOR3xp33_ASAP7_75t_SL g2725 ( 
.A(n_2136),
.B(n_91),
.C(n_92),
.Y(n_2725)
);

AOI22xp5_ASAP7_75t_L g2726 ( 
.A1(n_2149),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_2726)
);

INVx2_ASAP7_75t_L g2727 ( 
.A(n_2156),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_SL g2728 ( 
.A(n_2149),
.B(n_95),
.Y(n_2728)
);

INVx3_ASAP7_75t_L g2729 ( 
.A(n_1955),
.Y(n_2729)
);

AND2x4_ASAP7_75t_L g2730 ( 
.A(n_2036),
.B(n_96),
.Y(n_2730)
);

INVx4_ASAP7_75t_L g2731 ( 
.A(n_2179),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_1948),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_1963),
.B(n_96),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2156),
.Y(n_2734)
);

AND2x4_ASAP7_75t_L g2735 ( 
.A(n_2036),
.B(n_98),
.Y(n_2735)
);

NOR3xp33_ASAP7_75t_SL g2736 ( 
.A(n_2136),
.B(n_98),
.C(n_99),
.Y(n_2736)
);

INVx2_ASAP7_75t_L g2737 ( 
.A(n_2156),
.Y(n_2737)
);

AOI22xp5_ASAP7_75t_L g2738 ( 
.A1(n_2149),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2738)
);

NOR2x1_ASAP7_75t_L g2739 ( 
.A(n_2036),
.B(n_101),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_R g2740 ( 
.A(n_2046),
.B(n_804),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2156),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_1948),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2103),
.B(n_804),
.Y(n_2743)
);

BUFx2_ASAP7_75t_L g2744 ( 
.A(n_2027),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2156),
.Y(n_2745)
);

BUFx3_ASAP7_75t_L g2746 ( 
.A(n_2083),
.Y(n_2746)
);

AND2x6_ASAP7_75t_L g2747 ( 
.A(n_2214),
.B(n_102),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2547),
.B(n_102),
.Y(n_2748)
);

OR2x6_ASAP7_75t_L g2749 ( 
.A(n_2344),
.B(n_103),
.Y(n_2749)
);

BUFx2_ASAP7_75t_L g2750 ( 
.A(n_2344),
.Y(n_2750)
);

AOI21xp5_ASAP7_75t_L g2751 ( 
.A1(n_2275),
.A2(n_103),
.B(n_104),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2381),
.Y(n_2752)
);

BUFx3_ASAP7_75t_L g2753 ( 
.A(n_2703),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2285),
.B(n_104),
.Y(n_2754)
);

NOR2xp67_ASAP7_75t_L g2755 ( 
.A(n_2297),
.B(n_105),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2285),
.B(n_105),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2703),
.Y(n_2757)
);

NAND3xp33_ASAP7_75t_L g2758 ( 
.A(n_2534),
.B(n_106),
.C(n_108),
.Y(n_2758)
);

AOI21x1_ASAP7_75t_L g2759 ( 
.A1(n_2333),
.A2(n_106),
.B(n_108),
.Y(n_2759)
);

INVx2_ASAP7_75t_L g2760 ( 
.A(n_2657),
.Y(n_2760)
);

OR2x6_ASAP7_75t_L g2761 ( 
.A(n_2344),
.B(n_109),
.Y(n_2761)
);

OAI21x1_ASAP7_75t_L g2762 ( 
.A1(n_2372),
.A2(n_111),
.B(n_112),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2541),
.B(n_114),
.Y(n_2763)
);

AO21x2_ASAP7_75t_L g2764 ( 
.A1(n_2301),
.A2(n_115),
.B(n_116),
.Y(n_2764)
);

AO22x1_ASAP7_75t_L g2765 ( 
.A1(n_2396),
.A2(n_119),
.B1(n_115),
.B2(n_117),
.Y(n_2765)
);

OAI21x1_ASAP7_75t_L g2766 ( 
.A1(n_2372),
.A2(n_120),
.B(n_121),
.Y(n_2766)
);

OAI21x1_ASAP7_75t_L g2767 ( 
.A1(n_2301),
.A2(n_120),
.B(n_121),
.Y(n_2767)
);

AO31x2_ASAP7_75t_L g2768 ( 
.A1(n_2329),
.A2(n_2353),
.A3(n_2429),
.B(n_2660),
.Y(n_2768)
);

AND2x2_ASAP7_75t_L g2769 ( 
.A(n_2688),
.B(n_2706),
.Y(n_2769)
);

OAI22xp5_ASAP7_75t_L g2770 ( 
.A1(n_2364),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2770)
);

OAI21x1_ASAP7_75t_L g2771 ( 
.A1(n_2412),
.A2(n_123),
.B(n_124),
.Y(n_2771)
);

AND2x4_ASAP7_75t_L g2772 ( 
.A(n_2335),
.B(n_126),
.Y(n_2772)
);

AOI21x1_ASAP7_75t_SL g2773 ( 
.A1(n_2628),
.A2(n_126),
.B(n_128),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2708),
.B(n_128),
.Y(n_2774)
);

OAI21x1_ASAP7_75t_L g2775 ( 
.A1(n_2439),
.A2(n_130),
.B(n_131),
.Y(n_2775)
);

OAI21xp5_ASAP7_75t_L g2776 ( 
.A1(n_2353),
.A2(n_130),
.B(n_133),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2545),
.B(n_133),
.Y(n_2777)
);

OAI21x1_ASAP7_75t_L g2778 ( 
.A1(n_2296),
.A2(n_134),
.B(n_135),
.Y(n_2778)
);

OAI21x1_ASAP7_75t_L g2779 ( 
.A1(n_2296),
.A2(n_134),
.B(n_136),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2744),
.B(n_136),
.Y(n_2780)
);

OA21x2_ASAP7_75t_L g2781 ( 
.A1(n_2413),
.A2(n_137),
.B(n_138),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2280),
.B(n_138),
.Y(n_2782)
);

OAI21x1_ASAP7_75t_L g2783 ( 
.A1(n_2432),
.A2(n_139),
.B(n_140),
.Y(n_2783)
);

INVx1_ASAP7_75t_SL g2784 ( 
.A(n_2676),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2681),
.Y(n_2785)
);

AOI21xp5_ASAP7_75t_L g2786 ( 
.A1(n_2552),
.A2(n_140),
.B(n_141),
.Y(n_2786)
);

AO22x1_ASAP7_75t_L g2787 ( 
.A1(n_2603),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2273),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2552),
.A2(n_142),
.B(n_144),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_2409),
.B(n_144),
.Y(n_2790)
);

BUFx3_ASAP7_75t_L g2791 ( 
.A(n_2291),
.Y(n_2791)
);

BUFx2_ASAP7_75t_L g2792 ( 
.A(n_2337),
.Y(n_2792)
);

A2O1A1Ixp33_ASAP7_75t_L g2793 ( 
.A1(n_2364),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2699),
.A2(n_145),
.B(n_148),
.Y(n_2794)
);

OR2x2_ASAP7_75t_L g2795 ( 
.A(n_2417),
.B(n_149),
.Y(n_2795)
);

OAI21x1_ASAP7_75t_SL g2796 ( 
.A1(n_2702),
.A2(n_149),
.B(n_150),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2274),
.Y(n_2797)
);

NOR2x1_ASAP7_75t_SL g2798 ( 
.A(n_2348),
.B(n_150),
.Y(n_2798)
);

AOI21xp33_ASAP7_75t_L g2799 ( 
.A1(n_2461),
.A2(n_151),
.B(n_152),
.Y(n_2799)
);

AOI21x1_ASAP7_75t_L g2800 ( 
.A1(n_2281),
.A2(n_151),
.B(n_154),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2437),
.B(n_155),
.Y(n_2801)
);

AOI21xp5_ASAP7_75t_L g2802 ( 
.A1(n_2727),
.A2(n_156),
.B(n_157),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2276),
.Y(n_2803)
);

OAI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2461),
.A2(n_156),
.B(n_157),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2631),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.Y(n_2805)
);

OAI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2555),
.A2(n_2559),
.B(n_2535),
.Y(n_2806)
);

NOR2x1_ASAP7_75t_SL g2807 ( 
.A(n_2348),
.B(n_2378),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2283),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2734),
.Y(n_2809)
);

AND2x2_ASAP7_75t_L g2810 ( 
.A(n_2668),
.B(n_158),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2443),
.B(n_161),
.Y(n_2811)
);

OAI21x1_ASAP7_75t_L g2812 ( 
.A1(n_2302),
.A2(n_161),
.B(n_163),
.Y(n_2812)
);

AO21x1_ASAP7_75t_L g2813 ( 
.A1(n_2513),
.A2(n_163),
.B(n_164),
.Y(n_2813)
);

AO32x2_ASAP7_75t_L g2814 ( 
.A1(n_2329),
.A2(n_167),
.A3(n_164),
.B1(n_165),
.B2(n_168),
.Y(n_2814)
);

OAI21x1_ASAP7_75t_L g2815 ( 
.A1(n_2302),
.A2(n_167),
.B(n_168),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2737),
.A2(n_169),
.B(n_170),
.Y(n_2816)
);

INVx3_ASAP7_75t_L g2817 ( 
.A(n_2492),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2453),
.B(n_170),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2455),
.B(n_171),
.Y(n_2819)
);

OAI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2555),
.A2(n_171),
.B(n_172),
.Y(n_2820)
);

INVx4_ASAP7_75t_L g2821 ( 
.A(n_2664),
.Y(n_2821)
);

OAI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2741),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2457),
.B(n_2460),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2289),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2653),
.Y(n_2825)
);

AOI21x1_ASAP7_75t_L g2826 ( 
.A1(n_2628),
.A2(n_173),
.B(n_174),
.Y(n_2826)
);

INVx3_ASAP7_75t_L g2827 ( 
.A(n_2478),
.Y(n_2827)
);

OAI21x1_ASAP7_75t_L g2828 ( 
.A1(n_2592),
.A2(n_176),
.B(n_177),
.Y(n_2828)
);

OAI21x1_ASAP7_75t_L g2829 ( 
.A1(n_2592),
.A2(n_178),
.B(n_179),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2745),
.A2(n_2611),
.B(n_2635),
.Y(n_2830)
);

OAI21x1_ASAP7_75t_L g2831 ( 
.A1(n_2304),
.A2(n_2309),
.B(n_2306),
.Y(n_2831)
);

INVx4_ASAP7_75t_L g2832 ( 
.A(n_2664),
.Y(n_2832)
);

OAI21x1_ASAP7_75t_L g2833 ( 
.A1(n_2304),
.A2(n_178),
.B(n_179),
.Y(n_2833)
);

AO31x2_ASAP7_75t_L g2834 ( 
.A1(n_2629),
.A2(n_185),
.A3(n_182),
.B(n_183),
.Y(n_2834)
);

OR2x6_ASAP7_75t_L g2835 ( 
.A(n_2664),
.B(n_183),
.Y(n_2835)
);

AOI21xp33_ASAP7_75t_L g2836 ( 
.A1(n_2626),
.A2(n_186),
.B(n_187),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2710),
.B(n_186),
.Y(n_2837)
);

NAND2x1p5_ASAP7_75t_L g2838 ( 
.A(n_2286),
.B(n_188),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2655),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2311),
.B(n_189),
.Y(n_2840)
);

NAND2xp5_ASAP7_75t_L g2841 ( 
.A(n_2347),
.B(n_189),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2478),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2347),
.B(n_190),
.Y(n_2843)
);

OAI21x1_ASAP7_75t_L g2844 ( 
.A1(n_2309),
.A2(n_192),
.B(n_195),
.Y(n_2844)
);

OAI21x1_ASAP7_75t_L g2845 ( 
.A1(n_2325),
.A2(n_192),
.B(n_195),
.Y(n_2845)
);

OAI21xp33_ASAP7_75t_L g2846 ( 
.A1(n_2465),
.A2(n_196),
.B(n_197),
.Y(n_2846)
);

CKINVDCx8_ASAP7_75t_R g2847 ( 
.A(n_2327),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2394),
.B(n_197),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2663),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2667),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2406),
.B(n_198),
.Y(n_2851)
);

AND3x4_ASAP7_75t_L g2852 ( 
.A(n_2284),
.B(n_199),
.C(n_200),
.Y(n_2852)
);

HB1xp67_ASAP7_75t_L g2853 ( 
.A(n_2514),
.Y(n_2853)
);

AOI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2626),
.A2(n_200),
.B(n_202),
.Y(n_2854)
);

NOR2x1_ASAP7_75t_SL g2855 ( 
.A(n_2348),
.B(n_202),
.Y(n_2855)
);

CKINVDCx5p33_ASAP7_75t_R g2856 ( 
.A(n_2305),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2515),
.B(n_203),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2417),
.B(n_203),
.Y(n_2858)
);

AOI221xp5_ASAP7_75t_SL g2859 ( 
.A1(n_2606),
.A2(n_206),
.B1(n_204),
.B2(n_205),
.C(n_208),
.Y(n_2859)
);

AOI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2559),
.A2(n_204),
.B(n_208),
.Y(n_2860)
);

OAI22xp5_ASAP7_75t_L g2861 ( 
.A1(n_2378),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2861)
);

OAI21x1_ASAP7_75t_L g2862 ( 
.A1(n_2646),
.A2(n_210),
.B(n_211),
.Y(n_2862)
);

OA21x2_ASAP7_75t_L g2863 ( 
.A1(n_2413),
.A2(n_212),
.B(n_213),
.Y(n_2863)
);

A2O1A1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2436),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_2864)
);

AOI211x1_ASAP7_75t_L g2865 ( 
.A1(n_2485),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_SL g2866 ( 
.A(n_2323),
.B(n_217),
.Y(n_2866)
);

OAI22xp5_ASAP7_75t_L g2867 ( 
.A1(n_2330),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2538),
.B(n_219),
.Y(n_2868)
);

OAI21x1_ASAP7_75t_SL g2869 ( 
.A1(n_2540),
.A2(n_220),
.B(n_222),
.Y(n_2869)
);

INVx2_ASAP7_75t_L g2870 ( 
.A(n_2387),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2469),
.B(n_222),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2669),
.Y(n_2872)
);

AND2x4_ASAP7_75t_L g2873 ( 
.A(n_2666),
.B(n_224),
.Y(n_2873)
);

NOR2x1_ASAP7_75t_L g2874 ( 
.A(n_2378),
.B(n_224),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2484),
.B(n_225),
.Y(n_2875)
);

BUFx2_ASAP7_75t_L g2876 ( 
.A(n_2401),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_2740),
.B(n_225),
.Y(n_2877)
);

AO31x2_ASAP7_75t_L g2878 ( 
.A1(n_2517),
.A2(n_230),
.A3(n_227),
.B(n_229),
.Y(n_2878)
);

OAI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2529),
.A2(n_227),
.B(n_229),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2670),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2529),
.A2(n_230),
.B(n_231),
.Y(n_2881)
);

AOI21xp5_ASAP7_75t_L g2882 ( 
.A1(n_2535),
.A2(n_2610),
.B(n_2608),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2488),
.B(n_231),
.Y(n_2883)
);

INVxp67_ASAP7_75t_SL g2884 ( 
.A(n_2330),
.Y(n_2884)
);

AO31x2_ASAP7_75t_L g2885 ( 
.A1(n_2517),
.A2(n_234),
.A3(n_232),
.B(n_233),
.Y(n_2885)
);

AOI21xp5_ASAP7_75t_L g2886 ( 
.A1(n_2608),
.A2(n_232),
.B(n_233),
.Y(n_2886)
);

OA22x2_ASAP7_75t_L g2887 ( 
.A1(n_2427),
.A2(n_2651),
.B1(n_2665),
.B2(n_2644),
.Y(n_2887)
);

OR2x6_ASAP7_75t_L g2888 ( 
.A(n_2666),
.B(n_234),
.Y(n_2888)
);

OAI22xp5_ASAP7_75t_L g2889 ( 
.A1(n_2391),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2889)
);

AO21x2_ASAP7_75t_L g2890 ( 
.A1(n_2491),
.A2(n_2510),
.B(n_2449),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2495),
.B(n_236),
.Y(n_2891)
);

OAI21x1_ASAP7_75t_L g2892 ( 
.A1(n_2551),
.A2(n_237),
.B(n_238),
.Y(n_2892)
);

AOI21xp5_ASAP7_75t_L g2893 ( 
.A1(n_2610),
.A2(n_238),
.B(n_239),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2577),
.A2(n_240),
.B(n_241),
.Y(n_2894)
);

AO31x2_ASAP7_75t_L g2895 ( 
.A1(n_2550),
.A2(n_2463),
.A3(n_2448),
.B(n_2450),
.Y(n_2895)
);

CKINVDCx5p33_ASAP7_75t_R g2896 ( 
.A(n_2715),
.Y(n_2896)
);

OAI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2324),
.A2(n_2721),
.B1(n_2392),
.B2(n_2733),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2675),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2677),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2501),
.B(n_242),
.Y(n_2900)
);

OAI21xp5_ASAP7_75t_L g2901 ( 
.A1(n_2448),
.A2(n_242),
.B(n_243),
.Y(n_2901)
);

AOI21x1_ASAP7_75t_L g2902 ( 
.A1(n_2450),
.A2(n_243),
.B(n_244),
.Y(n_2902)
);

OAI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2476),
.A2(n_245),
.B(n_246),
.Y(n_2903)
);

AND2x4_ASAP7_75t_L g2904 ( 
.A(n_2731),
.B(n_245),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2512),
.B(n_246),
.Y(n_2905)
);

NAND3xp33_ASAP7_75t_SL g2906 ( 
.A(n_2637),
.B(n_247),
.C(n_248),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_L g2907 ( 
.A1(n_2324),
.A2(n_2678),
.B1(n_2685),
.B2(n_2674),
.Y(n_2907)
);

OAI21x1_ASAP7_75t_SL g2908 ( 
.A1(n_2540),
.A2(n_247),
.B(n_248),
.Y(n_2908)
);

BUFx6f_ASAP7_75t_L g2909 ( 
.A(n_2307),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_2522),
.B(n_249),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_SL g2911 ( 
.A(n_2503),
.B(n_250),
.Y(n_2911)
);

AOI21xp5_ASAP7_75t_L g2912 ( 
.A1(n_2577),
.A2(n_251),
.B(n_253),
.Y(n_2912)
);

HB1xp67_ASAP7_75t_L g2913 ( 
.A(n_2411),
.Y(n_2913)
);

INVxp67_ASAP7_75t_L g2914 ( 
.A(n_2711),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2523),
.B(n_2525),
.Y(n_2915)
);

OAI22xp5_ASAP7_75t_L g2916 ( 
.A1(n_2546),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_2288),
.B(n_255),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2288),
.B(n_2576),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2581),
.B(n_256),
.Y(n_2919)
);

AND2x4_ASAP7_75t_L g2920 ( 
.A(n_2731),
.B(n_257),
.Y(n_2920)
);

AND2x2_ASAP7_75t_L g2921 ( 
.A(n_2282),
.B(n_258),
.Y(n_2921)
);

NAND2x1_ASAP7_75t_L g2922 ( 
.A(n_2399),
.B(n_259),
.Y(n_2922)
);

OAI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2476),
.A2(n_259),
.B(n_260),
.Y(n_2923)
);

BUFx6f_ASAP7_75t_L g2924 ( 
.A(n_2307),
.Y(n_2924)
);

CKINVDCx5p33_ASAP7_75t_R g2925 ( 
.A(n_2345),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2356),
.Y(n_2926)
);

AO31x2_ASAP7_75t_L g2927 ( 
.A1(n_2550),
.A2(n_262),
.A3(n_260),
.B(n_261),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2585),
.B(n_262),
.Y(n_2928)
);

OAI21xp33_ASAP7_75t_L g2929 ( 
.A1(n_2534),
.A2(n_263),
.B(n_264),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_SL g2930 ( 
.A(n_2341),
.B(n_265),
.Y(n_2930)
);

AO31x2_ASAP7_75t_L g2931 ( 
.A1(n_2486),
.A2(n_267),
.A3(n_265),
.B(n_266),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_L g2932 ( 
.A(n_2586),
.B(n_2595),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2389),
.B(n_266),
.Y(n_2933)
);

A2O1A1Ixp33_ASAP7_75t_L g2934 ( 
.A1(n_2606),
.A2(n_2599),
.B(n_2430),
.C(n_2568),
.Y(n_2934)
);

NAND3x1_ASAP7_75t_L g2935 ( 
.A(n_2739),
.B(n_268),
.C(n_269),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2286),
.Y(n_2936)
);

OA21x2_ASAP7_75t_L g2937 ( 
.A1(n_2486),
.A2(n_270),
.B(n_271),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2684),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2578),
.A2(n_270),
.B(n_271),
.Y(n_2939)
);

OAI22xp5_ASAP7_75t_L g2940 ( 
.A1(n_2546),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2355),
.B(n_272),
.Y(n_2941)
);

AND2x4_ASAP7_75t_L g2942 ( 
.A(n_2553),
.B(n_275),
.Y(n_2942)
);

OAI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2511),
.A2(n_275),
.B(n_277),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2575),
.B(n_277),
.Y(n_2944)
);

NAND3xp33_ASAP7_75t_SL g2945 ( 
.A(n_2605),
.B(n_278),
.C(n_279),
.Y(n_2945)
);

AND2x2_ASAP7_75t_L g2946 ( 
.A(n_2361),
.B(n_2363),
.Y(n_2946)
);

OAI21x1_ASAP7_75t_L g2947 ( 
.A1(n_2278),
.A2(n_280),
.B(n_281),
.Y(n_2947)
);

AOI21x1_ASAP7_75t_L g2948 ( 
.A1(n_2462),
.A2(n_282),
.B(n_283),
.Y(n_2948)
);

BUFx2_ASAP7_75t_L g2949 ( 
.A(n_2692),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2687),
.Y(n_2950)
);

OR2x2_ASAP7_75t_L g2951 ( 
.A(n_2398),
.B(n_283),
.Y(n_2951)
);

OAI21x1_ASAP7_75t_L g2952 ( 
.A1(n_2279),
.A2(n_284),
.B(n_285),
.Y(n_2952)
);

INVx1_ASAP7_75t_SL g2953 ( 
.A(n_2292),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2689),
.B(n_284),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2393),
.B(n_286),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2693),
.B(n_286),
.Y(n_2956)
);

BUFx4_ASAP7_75t_SL g2957 ( 
.A(n_2293),
.Y(n_2957)
);

OR2x2_ASAP7_75t_L g2958 ( 
.A(n_2360),
.B(n_287),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2694),
.Y(n_2959)
);

AOI21xp5_ASAP7_75t_L g2960 ( 
.A1(n_2578),
.A2(n_288),
.B(n_289),
.Y(n_2960)
);

OAI21x1_ASAP7_75t_L g2961 ( 
.A1(n_2532),
.A2(n_288),
.B(n_289),
.Y(n_2961)
);

OAI22x1_ASAP7_75t_L g2962 ( 
.A1(n_2441),
.A2(n_2705),
.B1(n_2735),
.B2(n_2730),
.Y(n_2962)
);

AO31x2_ASAP7_75t_L g2963 ( 
.A1(n_2674),
.A2(n_2678),
.A3(n_2691),
.B(n_2685),
.Y(n_2963)
);

BUFx6f_ASAP7_75t_L g2964 ( 
.A(n_2307),
.Y(n_2964)
);

AO21x2_ASAP7_75t_L g2965 ( 
.A1(n_2579),
.A2(n_290),
.B(n_291),
.Y(n_2965)
);

BUFx2_ASAP7_75t_L g2966 ( 
.A(n_2692),
.Y(n_2966)
);

OAI21x1_ASAP7_75t_L g2967 ( 
.A1(n_2428),
.A2(n_290),
.B(n_291),
.Y(n_2967)
);

AOI21xp5_ASAP7_75t_L g2968 ( 
.A1(n_2579),
.A2(n_292),
.B(n_293),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2316),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2697),
.B(n_292),
.Y(n_2970)
);

OAI21x1_ASAP7_75t_L g2971 ( 
.A1(n_2615),
.A2(n_294),
.B(n_295),
.Y(n_2971)
);

NOR2xp67_ASAP7_75t_SL g2972 ( 
.A(n_2297),
.B(n_294),
.Y(n_2972)
);

BUFx2_ASAP7_75t_L g2973 ( 
.A(n_2672),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2625),
.B(n_2373),
.Y(n_2974)
);

OAI21xp5_ASAP7_75t_L g2975 ( 
.A1(n_2511),
.A2(n_2518),
.B(n_2445),
.Y(n_2975)
);

BUFx2_ASAP7_75t_L g2976 ( 
.A(n_2680),
.Y(n_2976)
);

NAND2x1_ASAP7_75t_L g2977 ( 
.A(n_2399),
.B(n_298),
.Y(n_2977)
);

NAND3xp33_ASAP7_75t_SL g2978 ( 
.A(n_2438),
.B(n_298),
.C(n_299),
.Y(n_2978)
);

OAI21xp5_ASAP7_75t_L g2979 ( 
.A1(n_2518),
.A2(n_300),
.B(n_301),
.Y(n_2979)
);

OAI21x1_ASAP7_75t_L g2980 ( 
.A1(n_2634),
.A2(n_301),
.B(n_302),
.Y(n_2980)
);

BUFx12f_ASAP7_75t_L g2981 ( 
.A(n_2458),
.Y(n_2981)
);

AND2x4_ASAP7_75t_L g2982 ( 
.A(n_2558),
.B(n_302),
.Y(n_2982)
);

AO31x2_ASAP7_75t_L g2983 ( 
.A1(n_2713),
.A2(n_305),
.A3(n_303),
.B(n_304),
.Y(n_2983)
);

OAI21x1_ASAP7_75t_L g2984 ( 
.A1(n_2634),
.A2(n_303),
.B(n_305),
.Y(n_2984)
);

OAI22x1_ASAP7_75t_L g2985 ( 
.A1(n_2705),
.A2(n_308),
.B1(n_306),
.B2(n_307),
.Y(n_2985)
);

BUFx3_ASAP7_75t_L g2986 ( 
.A(n_2299),
.Y(n_2986)
);

OAI21x1_ASAP7_75t_L g2987 ( 
.A1(n_2277),
.A2(n_306),
.B(n_308),
.Y(n_2987)
);

INVx5_ASAP7_75t_L g2988 ( 
.A(n_2747),
.Y(n_2988)
);

AOI21x1_ASAP7_75t_SL g2989 ( 
.A1(n_2468),
.A2(n_309),
.B(n_310),
.Y(n_2989)
);

OAI21x1_ASAP7_75t_L g2990 ( 
.A1(n_2277),
.A2(n_311),
.B(n_312),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2709),
.B(n_311),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2718),
.B(n_312),
.Y(n_2992)
);

AND2x4_ASAP7_75t_L g2993 ( 
.A(n_2561),
.B(n_313),
.Y(n_2993)
);

NOR2x1_ASAP7_75t_L g2994 ( 
.A(n_2399),
.B(n_314),
.Y(n_2994)
);

OAI21xp5_ASAP7_75t_L g2995 ( 
.A1(n_2445),
.A2(n_315),
.B(n_316),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_L g2996 ( 
.A(n_2313),
.Y(n_2996)
);

A2O1A1Ixp33_ASAP7_75t_L g2997 ( 
.A1(n_2499),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_2997)
);

AO22x2_ASAP7_75t_L g2998 ( 
.A1(n_2480),
.A2(n_319),
.B1(n_317),
.B2(n_318),
.Y(n_2998)
);

OAI21x1_ASAP7_75t_L g2999 ( 
.A1(n_2287),
.A2(n_2342),
.B(n_2319),
.Y(n_2999)
);

OAI21x1_ASAP7_75t_L g3000 ( 
.A1(n_2287),
.A2(n_320),
.B(n_322),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_L g3001 ( 
.A1(n_2322),
.A2(n_323),
.B1(n_320),
.B2(n_322),
.Y(n_3001)
);

OAI21x1_ASAP7_75t_L g3002 ( 
.A1(n_2319),
.A2(n_324),
.B(n_325),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2732),
.Y(n_3003)
);

AOI21xp33_ASAP7_75t_L g3004 ( 
.A1(n_2594),
.A2(n_326),
.B(n_328),
.Y(n_3004)
);

INVx1_ASAP7_75t_SL g3005 ( 
.A(n_2730),
.Y(n_3005)
);

NAND3xp33_ASAP7_75t_L g3006 ( 
.A(n_2527),
.B(n_326),
.C(n_328),
.Y(n_3006)
);

AND2x2_ASAP7_75t_L g3007 ( 
.A(n_2416),
.B(n_329),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_2742),
.B(n_330),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2369),
.A2(n_330),
.B(n_331),
.Y(n_3009)
);

A2O1A1Ixp33_ASAP7_75t_L g3010 ( 
.A1(n_2695),
.A2(n_334),
.B(n_332),
.C(n_333),
.Y(n_3010)
);

OAI21x1_ASAP7_75t_L g3011 ( 
.A1(n_2342),
.A2(n_333),
.B(n_334),
.Y(n_3011)
);

A2O1A1Ixp33_ASAP7_75t_L g3012 ( 
.A1(n_2704),
.A2(n_338),
.B(n_335),
.C(n_336),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2397),
.B(n_339),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2407),
.B(n_339),
.Y(n_3014)
);

OAI21x1_ASAP7_75t_L g3015 ( 
.A1(n_2354),
.A2(n_340),
.B(n_341),
.Y(n_3015)
);

CKINVDCx8_ASAP7_75t_R g3016 ( 
.A(n_2435),
.Y(n_3016)
);

BUFx6f_ASAP7_75t_L g3017 ( 
.A(n_2313),
.Y(n_3017)
);

AOI21xp5_ASAP7_75t_L g3018 ( 
.A1(n_2369),
.A2(n_340),
.B(n_341),
.Y(n_3018)
);

OAI21x1_ASAP7_75t_L g3019 ( 
.A1(n_2354),
.A2(n_343),
.B(n_344),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2318),
.B(n_343),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2320),
.B(n_345),
.Y(n_3021)
);

AND2x2_ASAP7_75t_L g3022 ( 
.A(n_2679),
.B(n_2724),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2365),
.B(n_2590),
.Y(n_3023)
);

BUFx2_ASAP7_75t_L g3024 ( 
.A(n_2707),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2336),
.B(n_347),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2346),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2531),
.B(n_347),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2543),
.B(n_348),
.Y(n_3028)
);

AO31x2_ASAP7_75t_L g3029 ( 
.A1(n_2607),
.A2(n_350),
.A3(n_348),
.B(n_349),
.Y(n_3029)
);

OAI21x1_ASAP7_75t_L g3030 ( 
.A1(n_2362),
.A2(n_350),
.B(n_351),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2404),
.B(n_352),
.Y(n_3031)
);

OAI21x1_ASAP7_75t_L g3032 ( 
.A1(n_2362),
.A2(n_352),
.B(n_354),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2349),
.Y(n_3033)
);

INVx3_ASAP7_75t_L g3034 ( 
.A(n_2393),
.Y(n_3034)
);

AOI22xp5_ASAP7_75t_L g3035 ( 
.A1(n_2480),
.A2(n_356),
.B1(n_354),
.B2(n_355),
.Y(n_3035)
);

INVx2_ASAP7_75t_SL g3036 ( 
.A(n_2312),
.Y(n_3036)
);

INVx2_ASAP7_75t_SL g3037 ( 
.A(n_2312),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2375),
.B(n_355),
.Y(n_3038)
);

AOI21xp5_ASAP7_75t_L g3039 ( 
.A1(n_2374),
.A2(n_357),
.B(n_358),
.Y(n_3039)
);

AND2x4_ASAP7_75t_L g3040 ( 
.A(n_2562),
.B(n_357),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2315),
.Y(n_3041)
);

OAI21x1_ASAP7_75t_L g3042 ( 
.A1(n_2414),
.A2(n_360),
.B(n_361),
.Y(n_3042)
);

OAI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2607),
.A2(n_360),
.B(n_361),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2366),
.B(n_362),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2395),
.Y(n_3045)
);

AOI21xp5_ASAP7_75t_L g3046 ( 
.A1(n_2374),
.A2(n_363),
.B(n_364),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2359),
.Y(n_3047)
);

AO31x2_ASAP7_75t_L g3048 ( 
.A1(n_2468),
.A2(n_366),
.A3(n_363),
.B(n_364),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2583),
.B(n_2477),
.Y(n_3049)
);

A2O1A1Ixp33_ASAP7_75t_L g3050 ( 
.A1(n_2743),
.A2(n_371),
.B(n_369),
.C(n_370),
.Y(n_3050)
);

AOI21xp5_ASAP7_75t_SL g3051 ( 
.A1(n_2422),
.A2(n_370),
.B(n_372),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2617),
.B(n_373),
.Y(n_3052)
);

AO22x2_ASAP7_75t_L g3053 ( 
.A1(n_2493),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_3053)
);

INVx1_ASAP7_75t_SL g3054 ( 
.A(n_2735),
.Y(n_3054)
);

BUFx2_ASAP7_75t_SL g3055 ( 
.A(n_2682),
.Y(n_3055)
);

AO31x2_ASAP7_75t_L g3056 ( 
.A1(n_2493),
.A2(n_378),
.A3(n_374),
.B(n_377),
.Y(n_3056)
);

OA22x2_ASAP7_75t_L g3057 ( 
.A1(n_2556),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_3057)
);

NAND2xp5_ASAP7_75t_L g3058 ( 
.A(n_2490),
.B(n_379),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2367),
.Y(n_3059)
);

BUFx6f_ASAP7_75t_L g3060 ( 
.A(n_2313),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2490),
.B(n_380),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2331),
.B(n_381),
.Y(n_3062)
);

BUFx3_ASAP7_75t_L g3063 ( 
.A(n_2383),
.Y(n_3063)
);

OAI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2485),
.A2(n_2377),
.B1(n_2508),
.B2(n_2420),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_SL g3065 ( 
.A(n_2395),
.B(n_382),
.Y(n_3065)
);

AND2x2_ASAP7_75t_L g3066 ( 
.A(n_2421),
.B(n_382),
.Y(n_3066)
);

OAI21x1_ASAP7_75t_L g3067 ( 
.A1(n_2656),
.A2(n_383),
.B(n_384),
.Y(n_3067)
);

OR2x6_ASAP7_75t_L g3068 ( 
.A(n_2293),
.B(n_384),
.Y(n_3068)
);

AOI21x1_ASAP7_75t_L g3069 ( 
.A1(n_2467),
.A2(n_385),
.B(n_386),
.Y(n_3069)
);

AO21x1_ASAP7_75t_L g3070 ( 
.A1(n_2508),
.A2(n_385),
.B(n_386),
.Y(n_3070)
);

AOI21xp33_ASAP7_75t_L g3071 ( 
.A1(n_2627),
.A2(n_387),
.B(n_388),
.Y(n_3071)
);

BUFx6f_ASAP7_75t_L g3072 ( 
.A(n_2332),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2331),
.B(n_387),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_L g3074 ( 
.A(n_2600),
.B(n_388),
.Y(n_3074)
);

NOR2xp33_ASAP7_75t_L g3075 ( 
.A(n_2464),
.B(n_389),
.Y(n_3075)
);

OA21x2_ASAP7_75t_L g3076 ( 
.A1(n_2527),
.A2(n_390),
.B(n_391),
.Y(n_3076)
);

OAI21x1_ASAP7_75t_L g3077 ( 
.A1(n_2656),
.A2(n_390),
.B(n_391),
.Y(n_3077)
);

OR2x2_ASAP7_75t_L g3078 ( 
.A(n_2720),
.B(n_392),
.Y(n_3078)
);

INVx1_ASAP7_75t_SL g3079 ( 
.A(n_2312),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2390),
.Y(n_3080)
);

OAI21xp5_ASAP7_75t_SL g3081 ( 
.A1(n_2290),
.A2(n_392),
.B(n_393),
.Y(n_3081)
);

INVx1_ASAP7_75t_SL g3082 ( 
.A(n_2648),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2423),
.B(n_393),
.Y(n_3083)
);

INVx1_ASAP7_75t_SL g3084 ( 
.A(n_2574),
.Y(n_3084)
);

AOI21xp5_ASAP7_75t_L g3085 ( 
.A1(n_2379),
.A2(n_394),
.B(n_395),
.Y(n_3085)
);

OA21x2_ASAP7_75t_L g3086 ( 
.A1(n_2650),
.A2(n_395),
.B(n_396),
.Y(n_3086)
);

AOI21xp5_ASAP7_75t_L g3087 ( 
.A1(n_2379),
.A2(n_396),
.B(n_397),
.Y(n_3087)
);

OAI21xp5_ASAP7_75t_L g3088 ( 
.A1(n_2565),
.A2(n_397),
.B(n_398),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_L g3089 ( 
.A1(n_2565),
.A2(n_398),
.B(n_399),
.Y(n_3089)
);

OA22x2_ASAP7_75t_L g3090 ( 
.A1(n_2556),
.A2(n_404),
.B1(n_401),
.B2(n_403),
.Y(n_3090)
);

O2A1O1Ixp5_ASAP7_75t_L g3091 ( 
.A1(n_2470),
.A2(n_406),
.B(n_401),
.C(n_405),
.Y(n_3091)
);

AOI221xp5_ASAP7_75t_L g3092 ( 
.A1(n_2326),
.A2(n_2298),
.B1(n_2419),
.B2(n_2662),
.C(n_2520),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2519),
.Y(n_3093)
);

OR2x6_ASAP7_75t_L g3094 ( 
.A(n_2293),
.B(n_406),
.Y(n_3094)
);

AOI21xp5_ASAP7_75t_L g3095 ( 
.A1(n_2415),
.A2(n_407),
.B(n_409),
.Y(n_3095)
);

BUFx6f_ASAP7_75t_L g3096 ( 
.A(n_2332),
.Y(n_3096)
);

CKINVDCx5p33_ASAP7_75t_R g3097 ( 
.A(n_2746),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_SL g3098 ( 
.A(n_2294),
.B(n_409),
.Y(n_3098)
);

OAI21x1_ASAP7_75t_L g3099 ( 
.A1(n_2658),
.A2(n_410),
.B(n_411),
.Y(n_3099)
);

AOI21x1_ASAP7_75t_SL g3100 ( 
.A1(n_2483),
.A2(n_410),
.B(n_412),
.Y(n_3100)
);

OAI21x1_ASAP7_75t_SL g3101 ( 
.A1(n_2471),
.A2(n_412),
.B(n_413),
.Y(n_3101)
);

AND2x2_ASAP7_75t_L g3102 ( 
.A(n_2509),
.B(n_413),
.Y(n_3102)
);

OAI21x1_ASAP7_75t_L g3103 ( 
.A1(n_2658),
.A2(n_414),
.B(n_415),
.Y(n_3103)
);

OAI21x1_ASAP7_75t_L g3104 ( 
.A1(n_2698),
.A2(n_414),
.B(n_416),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2601),
.B(n_416),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_2591),
.B(n_419),
.Y(n_3106)
);

OAI21x1_ASAP7_75t_L g3107 ( 
.A1(n_2698),
.A2(n_2729),
.B(n_2719),
.Y(n_3107)
);

OA21x2_ASAP7_75t_L g3108 ( 
.A1(n_2377),
.A2(n_422),
.B(n_423),
.Y(n_3108)
);

A2O1A1Ixp33_ASAP7_75t_L g3109 ( 
.A1(n_2536),
.A2(n_425),
.B(n_422),
.C(n_424),
.Y(n_3109)
);

NOR4xp25_ASAP7_75t_L g3110 ( 
.A(n_2654),
.B(n_2728),
.C(n_2690),
.D(n_2447),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2350),
.B(n_424),
.Y(n_3111)
);

OAI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2566),
.A2(n_426),
.B(n_427),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_2350),
.B(n_427),
.Y(n_3113)
);

AOI21xp5_ASAP7_75t_L g3114 ( 
.A1(n_2415),
.A2(n_428),
.B(n_430),
.Y(n_3114)
);

INVx2_ASAP7_75t_L g3115 ( 
.A(n_2338),
.Y(n_3115)
);

AO21x1_ASAP7_75t_L g3116 ( 
.A1(n_2502),
.A2(n_431),
.B(n_432),
.Y(n_3116)
);

OAI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2570),
.A2(n_431),
.B(n_433),
.Y(n_3117)
);

AOI21xp5_ASAP7_75t_L g3118 ( 
.A1(n_2424),
.A2(n_434),
.B(n_437),
.Y(n_3118)
);

OAI21x1_ASAP7_75t_L g3119 ( 
.A1(n_2729),
.A2(n_434),
.B(n_437),
.Y(n_3119)
);

INVx1_ASAP7_75t_SL g3120 ( 
.A(n_2563),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2352),
.B(n_438),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2332),
.Y(n_3122)
);

OAI21x1_ASAP7_75t_L g3123 ( 
.A1(n_2431),
.A2(n_438),
.B(n_439),
.Y(n_3123)
);

OAI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2570),
.A2(n_439),
.B(n_440),
.Y(n_3124)
);

AO31x2_ASAP7_75t_L g3125 ( 
.A1(n_2638),
.A2(n_442),
.A3(n_440),
.B(n_441),
.Y(n_3125)
);

OAI21x1_ASAP7_75t_L g3126 ( 
.A1(n_2431),
.A2(n_441),
.B(n_442),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2418),
.B(n_444),
.Y(n_3127)
);

OAI21x1_ASAP7_75t_L g3128 ( 
.A1(n_2456),
.A2(n_445),
.B(n_446),
.Y(n_3128)
);

AOI21xp5_ASAP7_75t_SL g3129 ( 
.A1(n_2422),
.A2(n_445),
.B(n_446),
.Y(n_3129)
);

OAI21x1_ASAP7_75t_L g3130 ( 
.A1(n_2456),
.A2(n_447),
.B(n_448),
.Y(n_3130)
);

A2O1A1Ixp33_ASAP7_75t_L g3131 ( 
.A1(n_2636),
.A2(n_451),
.B(n_449),
.C(n_450),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2352),
.B(n_450),
.Y(n_3132)
);

OAI21x1_ASAP7_75t_L g3133 ( 
.A1(n_2507),
.A2(n_451),
.B(n_452),
.Y(n_3133)
);

AO21x1_ASAP7_75t_L g3134 ( 
.A1(n_2686),
.A2(n_452),
.B(n_453),
.Y(n_3134)
);

NAND2xp5_ASAP7_75t_L g3135 ( 
.A(n_2358),
.B(n_453),
.Y(n_3135)
);

INVx3_ASAP7_75t_L g3136 ( 
.A(n_2310),
.Y(n_3136)
);

AOI21x1_ASAP7_75t_L g3137 ( 
.A1(n_2504),
.A2(n_454),
.B(n_455),
.Y(n_3137)
);

AOI21xp5_ASAP7_75t_L g3138 ( 
.A1(n_2424),
.A2(n_455),
.B(n_456),
.Y(n_3138)
);

NOR2xp33_ASAP7_75t_L g3139 ( 
.A(n_2425),
.B(n_2454),
.Y(n_3139)
);

OAI21x1_ASAP7_75t_SL g3140 ( 
.A1(n_2471),
.A2(n_456),
.B(n_457),
.Y(n_3140)
);

AOI21xp5_ASAP7_75t_L g3141 ( 
.A1(n_2426),
.A2(n_458),
.B(n_459),
.Y(n_3141)
);

INVx6_ASAP7_75t_L g3142 ( 
.A(n_2400),
.Y(n_3142)
);

AO31x2_ASAP7_75t_L g3143 ( 
.A1(n_2638),
.A2(n_462),
.A3(n_460),
.B(n_461),
.Y(n_3143)
);

NOR2xp67_ASAP7_75t_L g3144 ( 
.A(n_2418),
.B(n_460),
.Y(n_3144)
);

AO21x2_ASAP7_75t_L g3145 ( 
.A1(n_2357),
.A2(n_462),
.B(n_463),
.Y(n_3145)
);

OAI22xp5_ASAP7_75t_L g3146 ( 
.A1(n_2420),
.A2(n_467),
.B1(n_463),
.B2(n_466),
.Y(n_3146)
);

AO21x2_ASAP7_75t_L g3147 ( 
.A1(n_2975),
.A2(n_2357),
.B(n_2716),
.Y(n_3147)
);

OAI21x1_ASAP7_75t_SL g3148 ( 
.A1(n_2807),
.A2(n_2726),
.B(n_2717),
.Y(n_3148)
);

AOI22x1_ASAP7_75t_L g3149 ( 
.A1(n_2962),
.A2(n_2440),
.B1(n_2671),
.B2(n_2433),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_3023),
.B(n_2483),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_L g3151 ( 
.A(n_2806),
.B(n_2489),
.Y(n_3151)
);

HB1xp67_ASAP7_75t_L g3152 ( 
.A(n_2884),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2946),
.B(n_2835),
.Y(n_3153)
);

BUFx2_ASAP7_75t_SL g3154 ( 
.A(n_2847),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2988),
.B(n_2418),
.Y(n_3155)
);

NOR2xp33_ASAP7_75t_L g3156 ( 
.A(n_2821),
.B(n_2832),
.Y(n_3156)
);

AO21x2_ASAP7_75t_L g3157 ( 
.A1(n_2975),
.A2(n_2738),
.B(n_2530),
.Y(n_3157)
);

AOI22xp5_ASAP7_75t_L g3158 ( 
.A1(n_3064),
.A2(n_2509),
.B1(n_2521),
.B2(n_2489),
.Y(n_3158)
);

AO21x2_ASAP7_75t_L g3159 ( 
.A1(n_2882),
.A2(n_2539),
.B(n_2516),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2752),
.Y(n_3160)
);

OAI21x1_ASAP7_75t_L g3161 ( 
.A1(n_2999),
.A2(n_2524),
.B(n_2633),
.Y(n_3161)
);

OAI21x1_ASAP7_75t_L g3162 ( 
.A1(n_3107),
.A2(n_2548),
.B(n_2444),
.Y(n_3162)
);

OAI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2934),
.A2(n_2560),
.B(n_2358),
.Y(n_3163)
);

O2A1O1Ixp33_ASAP7_75t_SL g3164 ( 
.A1(n_2997),
.A2(n_2614),
.B(n_2560),
.C(n_2572),
.Y(n_3164)
);

AND2x2_ASAP7_75t_L g3165 ( 
.A(n_2835),
.B(n_2521),
.Y(n_3165)
);

AND2x4_ASAP7_75t_L g3166 ( 
.A(n_2988),
.B(n_2474),
.Y(n_3166)
);

NAND2xp5_ASAP7_75t_L g3167 ( 
.A(n_2806),
.B(n_2442),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2830),
.B(n_2442),
.Y(n_3168)
);

INVx2_ASAP7_75t_L g3169 ( 
.A(n_2784),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2932),
.Y(n_3170)
);

OA21x2_ASAP7_75t_L g3171 ( 
.A1(n_2767),
.A2(n_2701),
.B(n_2598),
.Y(n_3171)
);

OR2x2_ASAP7_75t_L g3172 ( 
.A(n_2918),
.B(n_2382),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_2988),
.B(n_2474),
.Y(n_3173)
);

OAI21x1_ASAP7_75t_L g3174 ( 
.A1(n_2773),
.A2(n_2481),
.B(n_2466),
.Y(n_3174)
);

AOI22xp33_ASAP7_75t_L g3175 ( 
.A1(n_2887),
.A2(n_2603),
.B1(n_2580),
.B2(n_2482),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2788),
.Y(n_3176)
);

OAI21x1_ASAP7_75t_L g3177 ( 
.A1(n_2989),
.A2(n_2496),
.B(n_2494),
.Y(n_3177)
);

OAI21x1_ASAP7_75t_L g3178 ( 
.A1(n_2831),
.A2(n_2639),
.B(n_2528),
.Y(n_3178)
);

OA21x2_ASAP7_75t_L g3179 ( 
.A1(n_2759),
.A2(n_2426),
.B(n_2588),
.Y(n_3179)
);

A2O1A1Ixp33_ASAP7_75t_L g3180 ( 
.A1(n_3081),
.A2(n_2712),
.B(n_2725),
.C(n_2714),
.Y(n_3180)
);

OAI21x1_ASAP7_75t_L g3181 ( 
.A1(n_3100),
.A2(n_2528),
.B(n_2526),
.Y(n_3181)
);

OAI21x1_ASAP7_75t_L g3182 ( 
.A1(n_2783),
.A2(n_2567),
.B(n_2526),
.Y(n_3182)
);

CKINVDCx20_ASAP7_75t_R g3183 ( 
.A(n_2753),
.Y(n_3183)
);

OAI21x1_ASAP7_75t_L g3184 ( 
.A1(n_2812),
.A2(n_2567),
.B(n_2542),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2797),
.Y(n_3185)
);

INVx3_ASAP7_75t_L g3186 ( 
.A(n_2749),
.Y(n_3186)
);

AOI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_3064),
.A2(n_2644),
.B1(n_2556),
.B2(n_2580),
.Y(n_3187)
);

AOI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_3082),
.A2(n_3092),
.B1(n_2835),
.B2(n_2821),
.Y(n_3188)
);

AO21x2_ASAP7_75t_L g3189 ( 
.A1(n_2804),
.A2(n_2661),
.B(n_2712),
.Y(n_3189)
);

NAND2xp5_ASAP7_75t_L g3190 ( 
.A(n_2890),
.B(n_2630),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2890),
.B(n_2630),
.Y(n_3191)
);

BUFx2_ASAP7_75t_L g3192 ( 
.A(n_2749),
.Y(n_3192)
);

NAND2xp5_ASAP7_75t_L g3193 ( 
.A(n_2963),
.B(n_2630),
.Y(n_3193)
);

BUFx3_ASAP7_75t_L g3194 ( 
.A(n_2791),
.Y(n_3194)
);

AO21x2_ASAP7_75t_L g3195 ( 
.A1(n_2804),
.A2(n_2661),
.B(n_2714),
.Y(n_3195)
);

BUFx8_ASAP7_75t_L g3196 ( 
.A(n_2981),
.Y(n_3196)
);

CKINVDCx5p33_ASAP7_75t_R g3197 ( 
.A(n_2757),
.Y(n_3197)
);

OR2x2_ASAP7_75t_L g3198 ( 
.A(n_2853),
.B(n_2482),
.Y(n_3198)
);

AND2x2_ASAP7_75t_L g3199 ( 
.A(n_2769),
.B(n_2612),
.Y(n_3199)
);

AOI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_2978),
.A2(n_2603),
.B1(n_2580),
.B2(n_2573),
.Y(n_3200)
);

OAI21x1_ASAP7_75t_L g3201 ( 
.A1(n_2815),
.A2(n_2567),
.B(n_2542),
.Y(n_3201)
);

AOI21x1_ASAP7_75t_L g3202 ( 
.A1(n_2897),
.A2(n_2385),
.B(n_2422),
.Y(n_3202)
);

HB1xp67_ASAP7_75t_L g3203 ( 
.A(n_2749),
.Y(n_3203)
);

OAI21xp5_ASAP7_75t_L g3204 ( 
.A1(n_2907),
.A2(n_2645),
.B(n_2643),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_2761),
.A2(n_2303),
.B(n_2542),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_2870),
.Y(n_3206)
);

OR2x2_ASAP7_75t_L g3207 ( 
.A(n_2951),
.B(n_2795),
.Y(n_3207)
);

OAI21x1_ASAP7_75t_L g3208 ( 
.A1(n_2778),
.A2(n_2542),
.B(n_2632),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_2761),
.A2(n_2303),
.B(n_2474),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2761),
.A2(n_2696),
.B(n_2474),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_2963),
.B(n_2760),
.Y(n_3211)
);

OA21x2_ASAP7_75t_L g3212 ( 
.A1(n_2762),
.A2(n_2649),
.B(n_2602),
.Y(n_3212)
);

CKINVDCx20_ASAP7_75t_R g3213 ( 
.A(n_2925),
.Y(n_3213)
);

AOI22xp33_ASAP7_75t_L g3214 ( 
.A1(n_3082),
.A2(n_2603),
.B1(n_2580),
.B2(n_2573),
.Y(n_3214)
);

OA21x2_ASAP7_75t_L g3215 ( 
.A1(n_2766),
.A2(n_2554),
.B(n_2604),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_3142),
.Y(n_3216)
);

AO21x2_ASAP7_75t_L g3217 ( 
.A1(n_2796),
.A2(n_2725),
.B(n_2368),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2803),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2963),
.B(n_2616),
.Y(n_3219)
);

HB1xp67_ASAP7_75t_L g3220 ( 
.A(n_3005),
.Y(n_3220)
);

OA21x2_ASAP7_75t_L g3221 ( 
.A1(n_2779),
.A2(n_2554),
.B(n_2609),
.Y(n_3221)
);

BUFx12f_ASAP7_75t_L g3222 ( 
.A(n_3097),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2785),
.B(n_2616),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_2808),
.Y(n_3224)
);

BUFx12f_ASAP7_75t_L g3225 ( 
.A(n_2856),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_2748),
.B(n_2612),
.Y(n_3226)
);

A2O1A1Ixp33_ASAP7_75t_L g3227 ( 
.A1(n_3081),
.A2(n_2723),
.B(n_2736),
.C(n_2563),
.Y(n_3227)
);

AOI32xp33_ASAP7_75t_L g3228 ( 
.A1(n_3083),
.A2(n_2446),
.A3(n_2620),
.B1(n_2371),
.B2(n_2402),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2824),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_2957),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2809),
.Y(n_3231)
);

CKINVDCx16_ASAP7_75t_R g3232 ( 
.A(n_2888),
.Y(n_3232)
);

NAND2x1p5_ASAP7_75t_L g3233 ( 
.A(n_2832),
.B(n_2696),
.Y(n_3233)
);

OAI21x1_ASAP7_75t_L g3234 ( 
.A1(n_2987),
.A2(n_2642),
.B(n_2640),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_2969),
.Y(n_3235)
);

BUFx3_ASAP7_75t_L g3236 ( 
.A(n_2876),
.Y(n_3236)
);

BUFx2_ASAP7_75t_L g3237 ( 
.A(n_2936),
.Y(n_3237)
);

INVx6_ASAP7_75t_L g3238 ( 
.A(n_3142),
.Y(n_3238)
);

AND2x4_ASAP7_75t_L g3239 ( 
.A(n_2772),
.B(n_2696),
.Y(n_3239)
);

BUFx4f_ASAP7_75t_SL g3240 ( 
.A(n_2949),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2825),
.Y(n_3241)
);

OAI21x1_ASAP7_75t_L g3242 ( 
.A1(n_2990),
.A2(n_2696),
.B(n_2621),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2839),
.Y(n_3243)
);

OAI21x1_ASAP7_75t_L g3244 ( 
.A1(n_2947),
.A2(n_2952),
.B(n_2800),
.Y(n_3244)
);

BUFx3_ASAP7_75t_L g3245 ( 
.A(n_3063),
.Y(n_3245)
);

OR2x2_ASAP7_75t_L g3246 ( 
.A(n_2858),
.B(n_2644),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_2768),
.B(n_2587),
.Y(n_3247)
);

OAI21x1_ASAP7_75t_L g3248 ( 
.A1(n_2892),
.A2(n_2622),
.B(n_2619),
.Y(n_3248)
);

AO21x2_ASAP7_75t_L g3249 ( 
.A1(n_2764),
.A2(n_2368),
.B(n_2620),
.Y(n_3249)
);

CKINVDCx8_ASAP7_75t_R g3250 ( 
.A(n_2966),
.Y(n_3250)
);

OAI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3058),
.A2(n_2446),
.B(n_2623),
.Y(n_3251)
);

OA21x2_ASAP7_75t_L g3252 ( 
.A1(n_2833),
.A2(n_2647),
.B(n_2624),
.Y(n_3252)
);

O2A1O1Ixp33_ASAP7_75t_L g3253 ( 
.A1(n_3109),
.A2(n_2403),
.B(n_2564),
.C(n_2544),
.Y(n_3253)
);

OA21x2_ASAP7_75t_L g3254 ( 
.A1(n_2844),
.A2(n_2647),
.B(n_2589),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3014),
.B(n_2384),
.Y(n_3255)
);

AO21x2_ASAP7_75t_L g3256 ( 
.A1(n_2764),
.A2(n_2673),
.B(n_2557),
.Y(n_3256)
);

INVx1_ASAP7_75t_SL g3257 ( 
.A(n_3005),
.Y(n_3257)
);

AND2x4_ASAP7_75t_L g3258 ( 
.A(n_2772),
.B(n_2380),
.Y(n_3258)
);

BUFx2_ASAP7_75t_L g3259 ( 
.A(n_2986),
.Y(n_3259)
);

AOI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_2929),
.A2(n_2747),
.B1(n_2597),
.B2(n_2472),
.Y(n_3260)
);

INVx3_ASAP7_75t_SL g3261 ( 
.A(n_2896),
.Y(n_3261)
);

BUFx2_ASAP7_75t_L g3262 ( 
.A(n_2913),
.Y(n_3262)
);

BUFx4_ASAP7_75t_SL g3263 ( 
.A(n_2888),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_2849),
.Y(n_3264)
);

BUFx3_ASAP7_75t_L g3265 ( 
.A(n_2817),
.Y(n_3265)
);

INVx2_ASAP7_75t_L g3266 ( 
.A(n_2926),
.Y(n_3266)
);

BUFx4f_ASAP7_75t_L g3267 ( 
.A(n_2888),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_2850),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_2914),
.B(n_2472),
.Y(n_3269)
);

BUFx2_ASAP7_75t_R g3270 ( 
.A(n_3016),
.Y(n_3270)
);

AO21x2_ASAP7_75t_L g3271 ( 
.A1(n_2869),
.A2(n_2557),
.B(n_2380),
.Y(n_3271)
);

OA21x2_ASAP7_75t_L g3272 ( 
.A1(n_2845),
.A2(n_2376),
.B(n_2351),
.Y(n_3272)
);

OAI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3061),
.A2(n_2582),
.B(n_2537),
.Y(n_3273)
);

A2O1A1Ixp33_ASAP7_75t_L g3274 ( 
.A1(n_2929),
.A2(n_2805),
.B(n_2846),
.C(n_2758),
.Y(n_3274)
);

OAI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2995),
.A2(n_2537),
.B(n_2747),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2768),
.B(n_2872),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_L g3277 ( 
.A(n_2768),
.B(n_2584),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_2880),
.Y(n_3278)
);

NAND2xp5_ASAP7_75t_L g3279 ( 
.A(n_2898),
.B(n_2584),
.Y(n_3279)
);

AOI21x1_ASAP7_75t_L g3280 ( 
.A1(n_2781),
.A2(n_2410),
.B(n_2376),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_2899),
.B(n_2571),
.Y(n_3281)
);

AND2x4_ASAP7_75t_L g3282 ( 
.A(n_3136),
.B(n_2310),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2974),
.B(n_2973),
.Y(n_3283)
);

INVx2_ASAP7_75t_L g3284 ( 
.A(n_3003),
.Y(n_3284)
);

BUFx3_ASAP7_75t_L g3285 ( 
.A(n_2817),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_2938),
.B(n_2571),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2950),
.Y(n_3287)
);

INVx4_ASAP7_75t_L g3288 ( 
.A(n_3068),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_2959),
.Y(n_3289)
);

INVx1_ASAP7_75t_SL g3290 ( 
.A(n_3054),
.Y(n_3290)
);

CKINVDCx20_ASAP7_75t_R g3291 ( 
.A(n_2976),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_2774),
.B(n_2500),
.Y(n_3292)
);

AND2x4_ASAP7_75t_L g3293 ( 
.A(n_2827),
.B(n_2351),
.Y(n_3293)
);

NOR2xp67_ASAP7_75t_L g3294 ( 
.A(n_3139),
.B(n_2451),
.Y(n_3294)
);

A2O1A1Ixp33_ASAP7_75t_L g3295 ( 
.A1(n_2805),
.A2(n_2569),
.B(n_2533),
.C(n_2549),
.Y(n_3295)
);

INVx3_ASAP7_75t_L g3296 ( 
.A(n_2827),
.Y(n_3296)
);

NOR2x1_ASAP7_75t_L g3297 ( 
.A(n_3068),
.B(n_2400),
.Y(n_3297)
);

INVx2_ASAP7_75t_L g3298 ( 
.A(n_3047),
.Y(n_3298)
);

A2O1A1Ixp33_ASAP7_75t_L g3299 ( 
.A1(n_2846),
.A2(n_2569),
.B(n_2505),
.C(n_2473),
.Y(n_3299)
);

AND2x2_ASAP7_75t_L g3300 ( 
.A(n_2780),
.B(n_2340),
.Y(n_3300)
);

INVx3_ASAP7_75t_L g3301 ( 
.A(n_2842),
.Y(n_3301)
);

OAI21x1_ASAP7_75t_L g3302 ( 
.A1(n_3133),
.A2(n_2487),
.B(n_2408),
.Y(n_3302)
);

AND2x4_ASAP7_75t_L g3303 ( 
.A(n_2842),
.B(n_2405),
.Y(n_3303)
);

INVx3_ASAP7_75t_L g3304 ( 
.A(n_3034),
.Y(n_3304)
);

NOR2xp67_ASAP7_75t_L g3305 ( 
.A(n_2873),
.B(n_2722),
.Y(n_3305)
);

OAI22xp33_ASAP7_75t_L g3306 ( 
.A1(n_3035),
.A2(n_2317),
.B1(n_2618),
.B2(n_2596),
.Y(n_3306)
);

OAI21x1_ASAP7_75t_L g3307 ( 
.A1(n_2828),
.A2(n_2487),
.B(n_2408),
.Y(n_3307)
);

INVx2_ASAP7_75t_L g3308 ( 
.A(n_3059),
.Y(n_3308)
);

OAI21x1_ASAP7_75t_L g3309 ( 
.A1(n_2829),
.A2(n_2498),
.B(n_2497),
.Y(n_3309)
);

OR2x2_ASAP7_75t_L g3310 ( 
.A(n_2915),
.B(n_2388),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_L g3311 ( 
.A1(n_2862),
.A2(n_2498),
.B(n_2497),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3026),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_3054),
.Y(n_3313)
);

NOR2xp67_ASAP7_75t_L g3314 ( 
.A(n_2873),
.B(n_2904),
.Y(n_3314)
);

OAI21x1_ASAP7_75t_L g3315 ( 
.A1(n_2980),
.A2(n_2984),
.B(n_2967),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3033),
.Y(n_3316)
);

AO31x2_ASAP7_75t_L g3317 ( 
.A1(n_3134),
.A2(n_2618),
.A3(n_2386),
.B(n_2498),
.Y(n_3317)
);

AND2x4_ASAP7_75t_L g3318 ( 
.A(n_3068),
.B(n_2405),
.Y(n_3318)
);

BUFx2_ASAP7_75t_L g3319 ( 
.A(n_3094),
.Y(n_3319)
);

OAI21x1_ASAP7_75t_L g3320 ( 
.A1(n_2771),
.A2(n_2652),
.B(n_2497),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3080),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_3115),
.Y(n_3322)
);

AO21x2_ASAP7_75t_L g3323 ( 
.A1(n_2908),
.A2(n_2328),
.B(n_2314),
.Y(n_3323)
);

AND2x2_ASAP7_75t_L g3324 ( 
.A(n_3013),
.B(n_2300),
.Y(n_3324)
);

AND2x4_ASAP7_75t_L g3325 ( 
.A(n_3094),
.B(n_2405),
.Y(n_3325)
);

AND2x4_ASAP7_75t_L g3326 ( 
.A(n_3094),
.B(n_2613),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_2921),
.B(n_2321),
.Y(n_3327)
);

A2O1A1Ixp33_ASAP7_75t_L g3328 ( 
.A1(n_2758),
.A2(n_2479),
.B(n_2475),
.C(n_2641),
.Y(n_3328)
);

AOI21xp5_ASAP7_75t_L g3329 ( 
.A1(n_2750),
.A2(n_2700),
.B(n_2659),
.Y(n_3329)
);

OAI21x1_ASAP7_75t_SL g3330 ( 
.A1(n_2798),
.A2(n_2334),
.B(n_2452),
.Y(n_3330)
);

OAI21x1_ASAP7_75t_L g3331 ( 
.A1(n_2775),
.A2(n_2863),
.B(n_2781),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_2792),
.Y(n_3332)
);

AOI21x1_ASAP7_75t_L g3333 ( 
.A1(n_2863),
.A2(n_2410),
.B(n_2328),
.Y(n_3333)
);

NOR2xp33_ASAP7_75t_L g3334 ( 
.A(n_3024),
.B(n_2459),
.Y(n_3334)
);

OAI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_2995),
.A2(n_2434),
.B(n_2339),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_2904),
.Y(n_3336)
);

AOI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_2874),
.A2(n_2700),
.B(n_2659),
.Y(n_3337)
);

OA21x2_ASAP7_75t_L g3338 ( 
.A1(n_2859),
.A2(n_2659),
.B(n_2652),
.Y(n_3338)
);

INVx5_ASAP7_75t_L g3339 ( 
.A(n_2909),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_SL g3340 ( 
.A(n_2920),
.Y(n_3340)
);

OA21x2_ASAP7_75t_L g3341 ( 
.A1(n_2859),
.A2(n_2683),
.B(n_2652),
.Y(n_3341)
);

OAI221xp5_ASAP7_75t_L g3342 ( 
.A1(n_3035),
.A2(n_2295),
.B1(n_2506),
.B2(n_2370),
.C(n_2343),
.Y(n_3342)
);

OAI21x1_ASAP7_75t_L g3343 ( 
.A1(n_3000),
.A2(n_2700),
.B(n_2683),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3041),
.Y(n_3344)
);

BUFx8_ASAP7_75t_SL g3345 ( 
.A(n_2920),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_2857),
.B(n_2459),
.Y(n_3346)
);

AO21x2_ASAP7_75t_L g3347 ( 
.A1(n_2776),
.A2(n_2434),
.B(n_2410),
.Y(n_3347)
);

OAI21x1_ASAP7_75t_L g3348 ( 
.A1(n_3002),
.A2(n_2593),
.B(n_2434),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_2823),
.Y(n_3349)
);

INVx2_ASAP7_75t_L g3350 ( 
.A(n_3086),
.Y(n_3350)
);

OAI21x1_ASAP7_75t_L g3351 ( 
.A1(n_3011),
.A2(n_3019),
.B(n_3015),
.Y(n_3351)
);

AOI22xp33_ASAP7_75t_L g3352 ( 
.A1(n_2813),
.A2(n_2434),
.B1(n_2571),
.B2(n_2593),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_2998),
.Y(n_3353)
);

OAI21x1_ASAP7_75t_L g3354 ( 
.A1(n_3030),
.A2(n_2593),
.B(n_2571),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_3086),
.Y(n_3355)
);

AOI22xp33_ASAP7_75t_SL g3356 ( 
.A1(n_2998),
.A2(n_2308),
.B1(n_469),
.B2(n_466),
.Y(n_3356)
);

OAI21x1_ASAP7_75t_L g3357 ( 
.A1(n_3032),
.A2(n_468),
.B(n_469),
.Y(n_3357)
);

BUFx3_ASAP7_75t_L g3358 ( 
.A(n_3036),
.Y(n_3358)
);

CKINVDCx5p33_ASAP7_75t_R g3359 ( 
.A(n_3075),
.Y(n_3359)
);

INVx3_ASAP7_75t_L g3360 ( 
.A(n_3034),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3031),
.B(n_468),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3053),
.Y(n_3362)
);

BUFx3_ASAP7_75t_L g3363 ( 
.A(n_3037),
.Y(n_3363)
);

INVx3_ASAP7_75t_L g3364 ( 
.A(n_3045),
.Y(n_3364)
);

OAI21x1_ASAP7_75t_L g3365 ( 
.A1(n_3042),
.A2(n_470),
.B(n_471),
.Y(n_3365)
);

OA21x2_ASAP7_75t_L g3366 ( 
.A1(n_3067),
.A2(n_470),
.B(n_471),
.Y(n_3366)
);

OAI21x1_ASAP7_75t_L g3367 ( 
.A1(n_3077),
.A2(n_3103),
.B(n_3099),
.Y(n_3367)
);

BUFx8_ASAP7_75t_L g3368 ( 
.A(n_3078),
.Y(n_3368)
);

NAND2x1p5_ASAP7_75t_L g3369 ( 
.A(n_3079),
.B(n_2994),
.Y(n_3369)
);

O2A1O1Ixp33_ASAP7_75t_L g3370 ( 
.A1(n_3010),
.A2(n_474),
.B(n_472),
.C(n_473),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_2944),
.B(n_474),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3053),
.Y(n_3372)
);

AO21x2_ASAP7_75t_L g3373 ( 
.A1(n_2776),
.A2(n_806),
.B(n_475),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3029),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3029),
.Y(n_3375)
);

OAI21x1_ASAP7_75t_L g3376 ( 
.A1(n_3104),
.A2(n_475),
.B(n_476),
.Y(n_3376)
);

NOR2x1_ASAP7_75t_SL g3377 ( 
.A(n_2861),
.B(n_478),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_3049),
.B(n_480),
.Y(n_3378)
);

OAI21x1_ASAP7_75t_L g3379 ( 
.A1(n_3119),
.A2(n_480),
.B(n_482),
.Y(n_3379)
);

AOI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_2916),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_3380)
);

OAI21x1_ASAP7_75t_L g3381 ( 
.A1(n_3123),
.A2(n_483),
.B(n_485),
.Y(n_3381)
);

INVx2_ASAP7_75t_L g3382 ( 
.A(n_3126),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3029),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2942),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_2941),
.B(n_485),
.Y(n_3385)
);

NAND2x1p5_ASAP7_75t_L g3386 ( 
.A(n_3079),
.B(n_486),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_2895),
.B(n_486),
.Y(n_3387)
);

NOR2xp33_ASAP7_75t_L g3388 ( 
.A(n_3022),
.B(n_487),
.Y(n_3388)
);

OA21x2_ASAP7_75t_L g3389 ( 
.A1(n_3128),
.A2(n_3130),
.B(n_2961),
.Y(n_3389)
);

AO21x2_ASAP7_75t_L g3390 ( 
.A1(n_2901),
.A2(n_487),
.B(n_488),
.Y(n_3390)
);

INVx3_ASAP7_75t_L g3391 ( 
.A(n_3045),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_2942),
.Y(n_3392)
);

OAI22xp5_ASAP7_75t_L g3393 ( 
.A1(n_3120),
.A2(n_492),
.B1(n_490),
.B2(n_491),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_2982),
.Y(n_3394)
);

OAI21x1_ASAP7_75t_L g3395 ( 
.A1(n_2902),
.A2(n_490),
.B(n_491),
.Y(n_3395)
);

OAI21x1_ASAP7_75t_L g3396 ( 
.A1(n_2826),
.A2(n_493),
.B(n_494),
.Y(n_3396)
);

OAI21x1_ASAP7_75t_L g3397 ( 
.A1(n_2994),
.A2(n_493),
.B(n_494),
.Y(n_3397)
);

AO21x2_ASAP7_75t_L g3398 ( 
.A1(n_2901),
.A2(n_806),
.B(n_495),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3084),
.A2(n_2855),
.B(n_2866),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_2982),
.Y(n_3400)
);

INVx1_ASAP7_75t_L g3401 ( 
.A(n_2993),
.Y(n_3401)
);

OA21x2_ASAP7_75t_L g3402 ( 
.A1(n_2903),
.A2(n_496),
.B(n_497),
.Y(n_3402)
);

OAI21x1_ASAP7_75t_L g3403 ( 
.A1(n_2971),
.A2(n_498),
.B(n_499),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_2937),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2993),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3040),
.Y(n_3406)
);

OAI21x1_ASAP7_75t_L g3407 ( 
.A1(n_2922),
.A2(n_499),
.B(n_500),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_3052),
.B(n_500),
.Y(n_3408)
);

OR2x2_ASAP7_75t_L g3409 ( 
.A(n_2958),
.B(n_501),
.Y(n_3409)
);

AOI21x1_ASAP7_75t_L g3410 ( 
.A1(n_2972),
.A2(n_501),
.B(n_502),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3040),
.Y(n_3411)
);

OAI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_3120),
.A2(n_504),
.B1(n_502),
.B2(n_503),
.Y(n_3412)
);

OAI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_2763),
.A2(n_505),
.B(n_506),
.Y(n_3413)
);

AOI22xp33_ASAP7_75t_L g3414 ( 
.A1(n_3070),
.A2(n_509),
.B1(n_507),
.B2(n_508),
.Y(n_3414)
);

OAI21xp5_ASAP7_75t_L g3415 ( 
.A1(n_2777),
.A2(n_507),
.B(n_508),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_2931),
.Y(n_3416)
);

AND2x4_ASAP7_75t_L g3417 ( 
.A(n_2755),
.B(n_510),
.Y(n_3417)
);

AOI222xp33_ASAP7_75t_L g3418 ( 
.A1(n_2906),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.C1(n_513),
.C2(n_514),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_2931),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_2931),
.Y(n_3420)
);

AOI22xp33_ASAP7_75t_L g3421 ( 
.A1(n_2945),
.A2(n_514),
.B1(n_511),
.B2(n_512),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3066),
.B(n_515),
.Y(n_3422)
);

NOR2xp33_ASAP7_75t_L g3423 ( 
.A(n_3093),
.B(n_516),
.Y(n_3423)
);

AO31x2_ASAP7_75t_L g3424 ( 
.A1(n_3116),
.A2(n_519),
.A3(n_517),
.B(n_518),
.Y(n_3424)
);

INVx3_ASAP7_75t_L g3425 ( 
.A(n_2909),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_2895),
.B(n_517),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2954),
.Y(n_3427)
);

AND2x4_ASAP7_75t_L g3428 ( 
.A(n_2755),
.B(n_518),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_2895),
.B(n_521),
.Y(n_3429)
);

AOI22xp33_ASAP7_75t_L g3430 ( 
.A1(n_3057),
.A2(n_525),
.B1(n_522),
.B2(n_524),
.Y(n_3430)
);

NOR2xp33_ASAP7_75t_L g3431 ( 
.A(n_3007),
.B(n_522),
.Y(n_3431)
);

OR2x6_ASAP7_75t_L g3432 ( 
.A(n_3051),
.B(n_524),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2956),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_2937),
.Y(n_3434)
);

OA21x2_ASAP7_75t_L g3435 ( 
.A1(n_2903),
.A2(n_525),
.B(n_526),
.Y(n_3435)
);

NOR2xp67_ASAP7_75t_L g3436 ( 
.A(n_2861),
.B(n_526),
.Y(n_3436)
);

AO31x2_ASAP7_75t_L g3437 ( 
.A1(n_3131),
.A2(n_529),
.A3(n_527),
.B(n_528),
.Y(n_3437)
);

INVx1_ASAP7_75t_SL g3438 ( 
.A(n_2953),
.Y(n_3438)
);

INVx3_ASAP7_75t_L g3439 ( 
.A(n_2924),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_2970),
.Y(n_3440)
);

AOI21x1_ASAP7_75t_L g3441 ( 
.A1(n_3144),
.A2(n_527),
.B(n_528),
.Y(n_3441)
);

INVx1_ASAP7_75t_SL g3442 ( 
.A(n_2953),
.Y(n_3442)
);

OAI21xp5_ASAP7_75t_L g3443 ( 
.A1(n_3009),
.A2(n_529),
.B(n_530),
.Y(n_3443)
);

OAI21x1_ASAP7_75t_L g3444 ( 
.A1(n_2977),
.A2(n_531),
.B(n_532),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_2838),
.B(n_532),
.Y(n_3445)
);

INVx8_ASAP7_75t_L g3446 ( 
.A(n_2924),
.Y(n_3446)
);

BUFx6f_ASAP7_75t_L g3447 ( 
.A(n_2924),
.Y(n_3447)
);

INVx1_ASAP7_75t_L g3448 ( 
.A(n_2991),
.Y(n_3448)
);

OAI21x1_ASAP7_75t_L g3449 ( 
.A1(n_3069),
.A2(n_533),
.B(n_534),
.Y(n_3449)
);

OAI21x1_ASAP7_75t_L g3450 ( 
.A1(n_3137),
.A2(n_533),
.B(n_535),
.Y(n_3450)
);

NAND2x1p5_ASAP7_75t_L g3451 ( 
.A(n_3084),
.B(n_536),
.Y(n_3451)
);

OAI22xp5_ASAP7_75t_L g3452 ( 
.A1(n_2865),
.A2(n_539),
.B1(n_537),
.B2(n_538),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_2965),
.Y(n_3453)
);

AND2x4_ASAP7_75t_L g3454 ( 
.A(n_3144),
.B(n_2964),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_2810),
.Y(n_3455)
);

OA21x2_ASAP7_75t_L g3456 ( 
.A1(n_2923),
.A2(n_2879),
.B(n_2820),
.Y(n_3456)
);

OAI221xp5_ASAP7_75t_L g3457 ( 
.A1(n_3062),
.A2(n_805),
.B1(n_540),
.B2(n_537),
.C(n_539),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_2964),
.Y(n_3458)
);

OAI21x1_ASAP7_75t_L g3459 ( 
.A1(n_3127),
.A2(n_540),
.B(n_542),
.Y(n_3459)
);

AOI22xp33_ASAP7_75t_L g3460 ( 
.A1(n_3090),
.A2(n_544),
.B1(n_542),
.B2(n_543),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_2992),
.Y(n_3461)
);

INVx4_ASAP7_75t_L g3462 ( 
.A(n_2964),
.Y(n_3462)
);

OAI21xp33_ASAP7_75t_SL g3463 ( 
.A1(n_2943),
.A2(n_2979),
.B(n_3043),
.Y(n_3463)
);

AND2x2_ASAP7_75t_L g3464 ( 
.A(n_2933),
.B(n_544),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_2965),
.Y(n_3465)
);

OAI21x1_ASAP7_75t_L g3466 ( 
.A1(n_2948),
.A2(n_545),
.B(n_546),
.Y(n_3466)
);

HB1xp67_ASAP7_75t_L g3467 ( 
.A(n_2996),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3150),
.B(n_2837),
.Y(n_3468)
);

HB1xp67_ASAP7_75t_L g3469 ( 
.A(n_3152),
.Y(n_3469)
);

OAI221xp5_ASAP7_75t_L g3470 ( 
.A1(n_3187),
.A2(n_3006),
.B1(n_2793),
.B2(n_3073),
.C(n_3111),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3199),
.B(n_3102),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3160),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3176),
.Y(n_3473)
);

AND2x2_ASAP7_75t_L g3474 ( 
.A(n_3292),
.B(n_3153),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3185),
.Y(n_3475)
);

INVx2_ASAP7_75t_L g3476 ( 
.A(n_3235),
.Y(n_3476)
);

AOI21xp5_ASAP7_75t_L g3477 ( 
.A1(n_3209),
.A2(n_3017),
.B(n_2996),
.Y(n_3477)
);

AND2x2_ASAP7_75t_L g3478 ( 
.A(n_3226),
.B(n_3044),
.Y(n_3478)
);

AOI221xp5_ASAP7_75t_L g3479 ( 
.A1(n_3306),
.A2(n_3378),
.B1(n_3423),
.B2(n_3457),
.C(n_3388),
.Y(n_3479)
);

NAND2xp33_ASAP7_75t_SL g3480 ( 
.A(n_3340),
.B(n_2852),
.Y(n_3480)
);

NAND2x1_ASAP7_75t_L g3481 ( 
.A(n_3288),
.B(n_3101),
.Y(n_3481)
);

AOI221xp5_ASAP7_75t_SL g3482 ( 
.A1(n_3306),
.A2(n_2985),
.B1(n_2770),
.B2(n_2782),
.C(n_2940),
.Y(n_3482)
);

CKINVDCx5p33_ASAP7_75t_R g3483 ( 
.A(n_3196),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3170),
.B(n_3349),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3232),
.B(n_3055),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3218),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3224),
.B(n_2865),
.Y(n_3487)
);

INVx3_ASAP7_75t_L g3488 ( 
.A(n_3233),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_3229),
.B(n_3043),
.Y(n_3489)
);

AOI22xp33_ASAP7_75t_L g3490 ( 
.A1(n_3267),
.A2(n_3006),
.B1(n_2930),
.B2(n_2911),
.Y(n_3490)
);

BUFx6f_ASAP7_75t_L g3491 ( 
.A(n_3446),
.Y(n_3491)
);

OAI22xp5_ASAP7_75t_L g3492 ( 
.A1(n_3267),
.A2(n_2935),
.B1(n_2940),
.B2(n_2916),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3241),
.B(n_3056),
.Y(n_3493)
);

AOI22xp33_ASAP7_75t_L g3494 ( 
.A1(n_3175),
.A2(n_3149),
.B1(n_3288),
.B2(n_3188),
.Y(n_3494)
);

AO21x2_ASAP7_75t_L g3495 ( 
.A1(n_3387),
.A2(n_3429),
.B(n_3426),
.Y(n_3495)
);

AO21x2_ASAP7_75t_L g3496 ( 
.A1(n_3387),
.A2(n_3140),
.B(n_2979),
.Y(n_3496)
);

NAND2x1_ASAP7_75t_L g3497 ( 
.A(n_3186),
.B(n_3129),
.Y(n_3497)
);

CKINVDCx5p33_ASAP7_75t_R g3498 ( 
.A(n_3196),
.Y(n_3498)
);

HB1xp67_ASAP7_75t_L g3499 ( 
.A(n_3152),
.Y(n_3499)
);

BUFx3_ASAP7_75t_L g3500 ( 
.A(n_3194),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3243),
.B(n_3056),
.Y(n_3501)
);

NAND3x1_ASAP7_75t_L g3502 ( 
.A(n_3297),
.B(n_2943),
.C(n_2879),
.Y(n_3502)
);

AND2x4_ASAP7_75t_L g3503 ( 
.A(n_3314),
.B(n_3056),
.Y(n_3503)
);

INVx3_ASAP7_75t_L g3504 ( 
.A(n_3233),
.Y(n_3504)
);

INVx4_ASAP7_75t_SL g3505 ( 
.A(n_3340),
.Y(n_3505)
);

BUFx6f_ASAP7_75t_L g3506 ( 
.A(n_3446),
.Y(n_3506)
);

OAI22xp33_ASAP7_75t_L g3507 ( 
.A1(n_3158),
.A2(n_3146),
.B1(n_2822),
.B2(n_2877),
.Y(n_3507)
);

CKINVDCx5p33_ASAP7_75t_R g3508 ( 
.A(n_3225),
.Y(n_3508)
);

AOI22xp33_ASAP7_75t_L g3509 ( 
.A1(n_3175),
.A2(n_3195),
.B1(n_3189),
.B2(n_3432),
.Y(n_3509)
);

BUFx3_ASAP7_75t_L g3510 ( 
.A(n_3245),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3361),
.B(n_2820),
.Y(n_3511)
);

AO22x1_ASAP7_75t_L g3512 ( 
.A1(n_3319),
.A2(n_2923),
.B1(n_3089),
.B2(n_3088),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3266),
.Y(n_3513)
);

BUFx2_ASAP7_75t_L g3514 ( 
.A(n_3262),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3264),
.Y(n_3515)
);

OAI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_3214),
.A2(n_2864),
.B1(n_3076),
.B2(n_3088),
.Y(n_3516)
);

AND2x2_ASAP7_75t_L g3517 ( 
.A(n_3385),
.B(n_3027),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3422),
.B(n_3028),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3268),
.Y(n_3519)
);

AOI221xp5_ASAP7_75t_L g3520 ( 
.A1(n_3457),
.A2(n_2836),
.B1(n_3004),
.B2(n_3071),
.C(n_2867),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3278),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3322),
.Y(n_3522)
);

AOI221xp5_ASAP7_75t_L g3523 ( 
.A1(n_3427),
.A2(n_3132),
.B1(n_3135),
.B2(n_3121),
.C(n_3113),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3189),
.A2(n_3076),
.B1(n_3108),
.B2(n_3098),
.Y(n_3524)
);

OAI21x1_ASAP7_75t_SL g3525 ( 
.A1(n_3377),
.A2(n_3117),
.B(n_3112),
.Y(n_3525)
);

A2O1A1Ixp33_ASAP7_75t_L g3526 ( 
.A1(n_3436),
.A2(n_3124),
.B(n_2751),
.C(n_3050),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3287),
.Y(n_3527)
);

NAND3xp33_ASAP7_75t_SL g3528 ( 
.A(n_3228),
.B(n_3124),
.C(n_3012),
.Y(n_3528)
);

AOI22xp5_ASAP7_75t_L g3529 ( 
.A1(n_3371),
.A2(n_2955),
.B1(n_3065),
.B2(n_3001),
.Y(n_3529)
);

OAI22x1_ASAP7_75t_L g3530 ( 
.A1(n_3203),
.A2(n_3108),
.B1(n_2787),
.B2(n_2843),
.Y(n_3530)
);

AOI22xp33_ASAP7_75t_L g3531 ( 
.A1(n_3195),
.A2(n_3039),
.B1(n_3046),
.B2(n_3018),
.Y(n_3531)
);

INVx3_ASAP7_75t_L g3532 ( 
.A(n_3250),
.Y(n_3532)
);

AOI22xp33_ASAP7_75t_L g3533 ( 
.A1(n_3432),
.A2(n_3087),
.B1(n_3095),
.B2(n_3085),
.Y(n_3533)
);

CKINVDCx6p67_ASAP7_75t_R g3534 ( 
.A(n_3261),
.Y(n_3534)
);

OAI22xp33_ASAP7_75t_L g3535 ( 
.A1(n_3380),
.A2(n_3432),
.B1(n_3203),
.B2(n_3192),
.Y(n_3535)
);

NAND2xp5_ASAP7_75t_L g3536 ( 
.A(n_3289),
.B(n_2917),
.Y(n_3536)
);

AOI22xp33_ASAP7_75t_L g3537 ( 
.A1(n_3353),
.A2(n_3118),
.B1(n_3138),
.B2(n_3114),
.Y(n_3537)
);

AOI22xp33_ASAP7_75t_L g3538 ( 
.A1(n_3362),
.A2(n_3141),
.B1(n_3145),
.B2(n_2889),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3312),
.Y(n_3539)
);

CKINVDCx5p33_ASAP7_75t_R g3540 ( 
.A(n_3183),
.Y(n_3540)
);

OR2x2_ASAP7_75t_L g3541 ( 
.A(n_3438),
.B(n_2754),
.Y(n_3541)
);

OAI221xp5_ASAP7_75t_L g3542 ( 
.A1(n_3227),
.A2(n_3110),
.B1(n_2928),
.B2(n_2919),
.C(n_2883),
.Y(n_3542)
);

INVx2_ASAP7_75t_SL g3543 ( 
.A(n_3240),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3316),
.B(n_3321),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3344),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3298),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_3205),
.A2(n_3275),
.B(n_3210),
.Y(n_3547)
);

INVx4_ASAP7_75t_SL g3548 ( 
.A(n_3240),
.Y(n_3548)
);

CKINVDCx20_ASAP7_75t_R g3549 ( 
.A(n_3345),
.Y(n_3549)
);

OAI211xp5_ASAP7_75t_L g3550 ( 
.A1(n_3356),
.A2(n_3106),
.B(n_2886),
.C(n_2893),
.Y(n_3550)
);

A2O1A1Ixp33_ASAP7_75t_L g3551 ( 
.A1(n_3463),
.A2(n_2786),
.B(n_2789),
.C(n_2854),
.Y(n_3551)
);

AND2x2_ASAP7_75t_L g3552 ( 
.A(n_3464),
.B(n_2814),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_L g3553 ( 
.A(n_3284),
.B(n_3125),
.Y(n_3553)
);

AOI22xp33_ASAP7_75t_L g3554 ( 
.A1(n_3372),
.A2(n_3145),
.B1(n_2799),
.B2(n_2912),
.Y(n_3554)
);

AOI22xp33_ASAP7_75t_L g3555 ( 
.A1(n_3356),
.A2(n_2939),
.B1(n_2960),
.B2(n_2894),
.Y(n_3555)
);

AND2x4_ASAP7_75t_L g3556 ( 
.A(n_3318),
.B(n_3060),
.Y(n_3556)
);

INVxp33_ASAP7_75t_L g3557 ( 
.A(n_3334),
.Y(n_3557)
);

AOI211xp5_ASAP7_75t_L g3558 ( 
.A1(n_3342),
.A2(n_3305),
.B(n_3180),
.C(n_3445),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_L g3559 ( 
.A(n_3342),
.B(n_2871),
.Y(n_3559)
);

INVx2_ASAP7_75t_L g3560 ( 
.A(n_3206),
.Y(n_3560)
);

INVx1_ASAP7_75t_SL g3561 ( 
.A(n_3259),
.Y(n_3561)
);

AOI22xp33_ASAP7_75t_L g3562 ( 
.A1(n_3255),
.A2(n_3165),
.B1(n_3204),
.B2(n_3200),
.Y(n_3562)
);

OR2x2_ASAP7_75t_L g3563 ( 
.A(n_3438),
.B(n_2756),
.Y(n_3563)
);

AND2x2_ASAP7_75t_L g3564 ( 
.A(n_3324),
.B(n_2814),
.Y(n_3564)
);

HB1xp67_ASAP7_75t_L g3565 ( 
.A(n_3442),
.Y(n_3565)
);

OAI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_3370),
.A2(n_3091),
.B(n_3110),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3231),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3308),
.Y(n_3568)
);

INVx1_ASAP7_75t_L g3569 ( 
.A(n_3223),
.Y(n_3569)
);

OR2x2_ASAP7_75t_L g3570 ( 
.A(n_3442),
.B(n_3125),
.Y(n_3570)
);

INVx1_ASAP7_75t_SL g3571 ( 
.A(n_3291),
.Y(n_3571)
);

OAI22xp5_ASAP7_75t_L g3572 ( 
.A1(n_3214),
.A2(n_2841),
.B1(n_2868),
.B2(n_2790),
.Y(n_3572)
);

AOI22xp33_ASAP7_75t_L g3573 ( 
.A1(n_3204),
.A2(n_2968),
.B1(n_2881),
.B2(n_2860),
.Y(n_3573)
);

AOI22xp33_ASAP7_75t_L g3574 ( 
.A1(n_3200),
.A2(n_2851),
.B1(n_2848),
.B2(n_2875),
.Y(n_3574)
);

A2O1A1Ixp33_ASAP7_75t_L g3575 ( 
.A1(n_3463),
.A2(n_2794),
.B(n_2816),
.C(n_2802),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3223),
.Y(n_3576)
);

NOR2xp33_ASAP7_75t_R g3577 ( 
.A(n_3197),
.B(n_3072),
.Y(n_3577)
);

OAI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_3260),
.A2(n_2801),
.B1(n_2818),
.B2(n_2811),
.Y(n_3578)
);

OAI22xp5_ASAP7_75t_L g3579 ( 
.A1(n_3260),
.A2(n_2819),
.B1(n_2900),
.B2(n_2891),
.Y(n_3579)
);

INVx2_ASAP7_75t_L g3580 ( 
.A(n_3169),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_3172),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3310),
.Y(n_3582)
);

AND2x2_ASAP7_75t_L g3583 ( 
.A(n_3327),
.B(n_2814),
.Y(n_3583)
);

OAI22xp33_ASAP7_75t_L g3584 ( 
.A1(n_3275),
.A2(n_2910),
.B1(n_2905),
.B2(n_3074),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3279),
.Y(n_3585)
);

OAI22xp33_ASAP7_75t_L g3586 ( 
.A1(n_3246),
.A2(n_3105),
.B1(n_2840),
.B2(n_3020),
.Y(n_3586)
);

INVx3_ASAP7_75t_SL g3587 ( 
.A(n_3230),
.Y(n_3587)
);

AOI22xp33_ASAP7_75t_L g3588 ( 
.A1(n_3300),
.A2(n_3008),
.B1(n_3025),
.B2(n_3021),
.Y(n_3588)
);

OAI222xp33_ASAP7_75t_L g3589 ( 
.A1(n_3451),
.A2(n_3038),
.B1(n_2765),
.B2(n_2927),
.C1(n_2885),
.C2(n_2878),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_L g3590 ( 
.A(n_3207),
.B(n_3125),
.Y(n_3590)
);

AND2x4_ASAP7_75t_L g3591 ( 
.A(n_3325),
.B(n_3239),
.Y(n_3591)
);

NAND2x1p5_ASAP7_75t_L g3592 ( 
.A(n_3265),
.B(n_3096),
.Y(n_3592)
);

CKINVDCx16_ASAP7_75t_R g3593 ( 
.A(n_3213),
.Y(n_3593)
);

AND2x6_ASAP7_75t_L g3594 ( 
.A(n_3239),
.B(n_3096),
.Y(n_3594)
);

NOR2xp33_ASAP7_75t_L g3595 ( 
.A(n_3346),
.B(n_3283),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3446),
.Y(n_3596)
);

AOI221xp5_ASAP7_75t_L g3597 ( 
.A1(n_3433),
.A2(n_3048),
.B1(n_3143),
.B2(n_2983),
.C(n_2885),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3440),
.B(n_3143),
.Y(n_3598)
);

INVx3_ASAP7_75t_L g3599 ( 
.A(n_3285),
.Y(n_3599)
);

BUFx2_ASAP7_75t_L g3600 ( 
.A(n_3332),
.Y(n_3600)
);

BUFx12f_ASAP7_75t_L g3601 ( 
.A(n_3222),
.Y(n_3601)
);

INVx2_ASAP7_75t_L g3602 ( 
.A(n_3281),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_L g3603 ( 
.A1(n_3151),
.A2(n_3122),
.B1(n_3096),
.B2(n_3143),
.Y(n_3603)
);

CKINVDCx5p33_ASAP7_75t_R g3604 ( 
.A(n_3270),
.Y(n_3604)
);

NAND2xp5_ASAP7_75t_L g3605 ( 
.A(n_3448),
.B(n_3048),
.Y(n_3605)
);

OR2x2_ASAP7_75t_L g3606 ( 
.A(n_3198),
.B(n_2983),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3281),
.Y(n_3607)
);

AOI22xp33_ASAP7_75t_L g3608 ( 
.A1(n_3151),
.A2(n_3167),
.B1(n_3408),
.B2(n_3431),
.Y(n_3608)
);

INVxp67_ASAP7_75t_L g3609 ( 
.A(n_3237),
.Y(n_3609)
);

INVx6_ASAP7_75t_L g3610 ( 
.A(n_3238),
.Y(n_3610)
);

BUFx4f_ASAP7_75t_SL g3611 ( 
.A(n_3236),
.Y(n_3611)
);

INVx4_ASAP7_75t_L g3612 ( 
.A(n_3238),
.Y(n_3612)
);

OR2x6_ASAP7_75t_L g3613 ( 
.A(n_3154),
.B(n_2878),
.Y(n_3613)
);

AOI221xp5_ASAP7_75t_L g3614 ( 
.A1(n_3461),
.A2(n_3048),
.B1(n_2983),
.B2(n_2885),
.C(n_2927),
.Y(n_3614)
);

AND2x4_ASAP7_75t_L g3615 ( 
.A(n_3258),
.B(n_2878),
.Y(n_3615)
);

NAND2xp33_ASAP7_75t_SL g3616 ( 
.A(n_3263),
.B(n_3336),
.Y(n_3616)
);

AOI22xp5_ASAP7_75t_L g3617 ( 
.A1(n_3384),
.A2(n_2927),
.B1(n_2834),
.B2(n_547),
.Y(n_3617)
);

AOI22xp33_ASAP7_75t_L g3618 ( 
.A1(n_3167),
.A2(n_548),
.B1(n_545),
.B2(n_546),
.Y(n_3618)
);

OR2x6_ASAP7_75t_L g3619 ( 
.A(n_3263),
.B(n_548),
.Y(n_3619)
);

OAI22xp5_ASAP7_75t_SL g3620 ( 
.A1(n_3359),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.Y(n_3620)
);

BUFx2_ASAP7_75t_L g3621 ( 
.A(n_3326),
.Y(n_3621)
);

BUFx2_ASAP7_75t_L g3622 ( 
.A(n_3326),
.Y(n_3622)
);

NAND3x1_ASAP7_75t_L g3623 ( 
.A(n_3156),
.B(n_551),
.C(n_552),
.Y(n_3623)
);

INVx1_ASAP7_75t_L g3624 ( 
.A(n_3286),
.Y(n_3624)
);

OAI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3451),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.Y(n_3625)
);

BUFx12f_ASAP7_75t_L g3626 ( 
.A(n_3368),
.Y(n_3626)
);

CKINVDCx5p33_ASAP7_75t_R g3627 ( 
.A(n_3270),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3455),
.B(n_554),
.Y(n_3628)
);

INVx3_ASAP7_75t_L g3629 ( 
.A(n_3155),
.Y(n_3629)
);

NAND2x1_ASAP7_75t_L g3630 ( 
.A(n_3205),
.B(n_555),
.Y(n_3630)
);

OAI22xp5_ASAP7_75t_L g3631 ( 
.A1(n_3430),
.A2(n_558),
.B1(n_555),
.B2(n_557),
.Y(n_3631)
);

INVx1_ASAP7_75t_L g3632 ( 
.A(n_3286),
.Y(n_3632)
);

OAI22xp5_ASAP7_75t_L g3633 ( 
.A1(n_3430),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_3633)
);

OR2x2_ASAP7_75t_L g3634 ( 
.A(n_3257),
.B(n_559),
.Y(n_3634)
);

NAND2x1p5_ASAP7_75t_L g3635 ( 
.A(n_3339),
.B(n_560),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3392),
.B(n_561),
.Y(n_3636)
);

HB1xp67_ASAP7_75t_L g3637 ( 
.A(n_3220),
.Y(n_3637)
);

AO31x2_ASAP7_75t_L g3638 ( 
.A1(n_3382),
.A2(n_3434),
.A3(n_3404),
.B(n_3453),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3190),
.Y(n_3639)
);

NOR2xp33_ASAP7_75t_L g3640 ( 
.A(n_3368),
.B(n_564),
.Y(n_3640)
);

OA21x2_ASAP7_75t_L g3641 ( 
.A1(n_3331),
.A2(n_565),
.B(n_566),
.Y(n_3641)
);

AOI22xp33_ASAP7_75t_L g3642 ( 
.A1(n_3394),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_3642)
);

AND2x4_ASAP7_75t_L g3643 ( 
.A(n_3258),
.B(n_567),
.Y(n_3643)
);

AOI22xp33_ASAP7_75t_L g3644 ( 
.A1(n_3400),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3644)
);

AND2x2_ASAP7_75t_L g3645 ( 
.A(n_3409),
.B(n_570),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3220),
.Y(n_3646)
);

HB1xp67_ASAP7_75t_L g3647 ( 
.A(n_3313),
.Y(n_3647)
);

CKINVDCx5p33_ASAP7_75t_R g3648 ( 
.A(n_3269),
.Y(n_3648)
);

AND2x2_ASAP7_75t_L g3649 ( 
.A(n_3216),
.B(n_805),
.Y(n_3649)
);

OAI22xp33_ASAP7_75t_L g3650 ( 
.A1(n_3393),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_3650)
);

NAND3xp33_ASAP7_75t_L g3651 ( 
.A(n_3418),
.B(n_574),
.C(n_575),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3313),
.Y(n_3652)
);

AOI22xp33_ASAP7_75t_L g3653 ( 
.A1(n_3401),
.A2(n_579),
.B1(n_577),
.B2(n_578),
.Y(n_3653)
);

BUFx4f_ASAP7_75t_SL g3654 ( 
.A(n_3358),
.Y(n_3654)
);

OAI22xp33_ASAP7_75t_L g3655 ( 
.A1(n_3393),
.A2(n_581),
.B1(n_577),
.B2(n_580),
.Y(n_3655)
);

NAND3x1_ASAP7_75t_L g3656 ( 
.A(n_3210),
.B(n_3360),
.C(n_3304),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3190),
.Y(n_3657)
);

INVx3_ASAP7_75t_L g3658 ( 
.A(n_3166),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3405),
.A2(n_583),
.B1(n_581),
.B2(n_582),
.Y(n_3659)
);

OR2x6_ASAP7_75t_L g3660 ( 
.A(n_3330),
.B(n_582),
.Y(n_3660)
);

AOI22xp33_ASAP7_75t_L g3661 ( 
.A1(n_3406),
.A2(n_585),
.B1(n_583),
.B2(n_584),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3411),
.Y(n_3662)
);

AOI22xp33_ASAP7_75t_L g3663 ( 
.A1(n_3251),
.A2(n_3418),
.B1(n_3460),
.B2(n_3163),
.Y(n_3663)
);

OAI22xp5_ASAP7_75t_L g3664 ( 
.A1(n_3460),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3251),
.B(n_587),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3386),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3191),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3191),
.Y(n_3668)
);

CKINVDCx5p33_ASAP7_75t_R g3669 ( 
.A(n_3363),
.Y(n_3669)
);

INVx1_ASAP7_75t_L g3670 ( 
.A(n_3386),
.Y(n_3670)
);

NOR2xp33_ASAP7_75t_L g3671 ( 
.A(n_3216),
.B(n_589),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3295),
.B(n_590),
.Y(n_3672)
);

OR2x6_ASAP7_75t_L g3673 ( 
.A(n_3294),
.B(n_3417),
.Y(n_3673)
);

BUFx3_ASAP7_75t_L g3674 ( 
.A(n_3304),
.Y(n_3674)
);

AOI22xp33_ASAP7_75t_L g3675 ( 
.A1(n_3163),
.A2(n_593),
.B1(n_591),
.B2(n_592),
.Y(n_3675)
);

AOI22xp33_ASAP7_75t_L g3676 ( 
.A1(n_3456),
.A2(n_594),
.B1(n_591),
.B2(n_592),
.Y(n_3676)
);

NOR2xp33_ASAP7_75t_L g3677 ( 
.A(n_3360),
.B(n_595),
.Y(n_3677)
);

AOI22xp33_ASAP7_75t_L g3678 ( 
.A1(n_3456),
.A2(n_599),
.B1(n_596),
.B2(n_598),
.Y(n_3678)
);

AND2x2_ASAP7_75t_L g3679 ( 
.A(n_3257),
.B(n_803),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_SL g3680 ( 
.A1(n_3335),
.A2(n_3452),
.B1(n_3148),
.B2(n_3428),
.Y(n_3680)
);

AO21x2_ASAP7_75t_L g3681 ( 
.A1(n_3426),
.A2(n_600),
.B(n_601),
.Y(n_3681)
);

AOI22xp33_ASAP7_75t_L g3682 ( 
.A1(n_3335),
.A2(n_3452),
.B1(n_3421),
.B2(n_3217),
.Y(n_3682)
);

NAND3xp33_ASAP7_75t_SL g3683 ( 
.A(n_3299),
.B(n_602),
.C(n_603),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3217),
.A2(n_605),
.B1(n_602),
.B2(n_604),
.Y(n_3684)
);

AND2x2_ASAP7_75t_L g3685 ( 
.A(n_3290),
.B(n_803),
.Y(n_3685)
);

AOI22xp5_ASAP7_75t_L g3686 ( 
.A1(n_3412),
.A2(n_606),
.B1(n_604),
.B2(n_605),
.Y(n_3686)
);

AOI21xp33_ASAP7_75t_SL g3687 ( 
.A1(n_3412),
.A2(n_606),
.B(n_607),
.Y(n_3687)
);

INVx2_ASAP7_75t_SL g3688 ( 
.A(n_3364),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3211),
.Y(n_3689)
);

OAI221xp5_ASAP7_75t_L g3690 ( 
.A1(n_3273),
.A2(n_609),
.B1(n_610),
.B2(n_611),
.C(n_614),
.Y(n_3690)
);

HB1xp67_ASAP7_75t_L g3691 ( 
.A(n_3290),
.Y(n_3691)
);

AOI22xp33_ASAP7_75t_L g3692 ( 
.A1(n_3171),
.A2(n_615),
.B1(n_609),
.B2(n_610),
.Y(n_3692)
);

A2O1A1Ixp33_ASAP7_75t_L g3693 ( 
.A1(n_3274),
.A2(n_617),
.B(n_615),
.C(n_616),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3364),
.B(n_616),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3211),
.Y(n_3695)
);

OAI22xp5_ASAP7_75t_L g3696 ( 
.A1(n_3414),
.A2(n_621),
.B1(n_618),
.B2(n_620),
.Y(n_3696)
);

OR2x2_ASAP7_75t_L g3697 ( 
.A(n_3219),
.B(n_3168),
.Y(n_3697)
);

OR2x2_ASAP7_75t_L g3698 ( 
.A(n_3219),
.B(n_618),
.Y(n_3698)
);

AND2x6_ASAP7_75t_L g3699 ( 
.A(n_3166),
.B(n_620),
.Y(n_3699)
);

OR2x6_ASAP7_75t_L g3700 ( 
.A(n_3417),
.B(n_621),
.Y(n_3700)
);

OAI22xp5_ASAP7_75t_L g3701 ( 
.A1(n_3414),
.A2(n_624),
.B1(n_622),
.B2(n_623),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_SL g3702 ( 
.A(n_3399),
.B(n_622),
.Y(n_3702)
);

AOI22xp33_ASAP7_75t_L g3703 ( 
.A1(n_3171),
.A2(n_626),
.B1(n_623),
.B2(n_625),
.Y(n_3703)
);

AOI22xp33_ASAP7_75t_L g3704 ( 
.A1(n_3147),
.A2(n_625),
.B1(n_626),
.B2(n_628),
.Y(n_3704)
);

INVx2_ASAP7_75t_SL g3705 ( 
.A(n_3391),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3424),
.Y(n_3706)
);

AO21x2_ASAP7_75t_L g3707 ( 
.A1(n_3429),
.A2(n_630),
.B(n_631),
.Y(n_3707)
);

INVx6_ASAP7_75t_L g3708 ( 
.A(n_3339),
.Y(n_3708)
);

AOI22xp33_ASAP7_75t_SL g3709 ( 
.A1(n_3428),
.A2(n_631),
.B1(n_632),
.B2(n_635),
.Y(n_3709)
);

AOI22xp33_ASAP7_75t_L g3710 ( 
.A1(n_3528),
.A2(n_3492),
.B1(n_3535),
.B2(n_3559),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_L g3711 ( 
.A1(n_3479),
.A2(n_3147),
.B1(n_3347),
.B2(n_3271),
.Y(n_3711)
);

OAI21xp33_ASAP7_75t_L g3712 ( 
.A1(n_3509),
.A2(n_3352),
.B(n_3247),
.Y(n_3712)
);

AOI22xp33_ASAP7_75t_SL g3713 ( 
.A1(n_3699),
.A2(n_3369),
.B1(n_3256),
.B2(n_3271),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3476),
.Y(n_3714)
);

AOI22xp33_ASAP7_75t_SL g3715 ( 
.A1(n_3699),
.A2(n_3369),
.B1(n_3256),
.B2(n_3402),
.Y(n_3715)
);

AOI22xp33_ASAP7_75t_SL g3716 ( 
.A1(n_3699),
.A2(n_3435),
.B1(n_3402),
.B2(n_3338),
.Y(n_3716)
);

INVx8_ASAP7_75t_L g3717 ( 
.A(n_3626),
.Y(n_3717)
);

OAI33xp33_ASAP7_75t_L g3718 ( 
.A1(n_3620),
.A2(n_3247),
.A3(n_3420),
.B1(n_3419),
.B2(n_3416),
.B3(n_3374),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_L g3719 ( 
.A(n_3557),
.B(n_3282),
.Y(n_3719)
);

AOI221xp5_ASAP7_75t_L g3720 ( 
.A1(n_3586),
.A2(n_3370),
.B1(n_3253),
.B2(n_3415),
.C(n_3413),
.Y(n_3720)
);

AOI22xp33_ASAP7_75t_L g3721 ( 
.A1(n_3651),
.A2(n_3347),
.B1(n_3157),
.B2(n_3443),
.Y(n_3721)
);

AND2x2_ASAP7_75t_L g3722 ( 
.A(n_3474),
.B(n_3467),
.Y(n_3722)
);

OAI21xp33_ASAP7_75t_L g3723 ( 
.A1(n_3619),
.A2(n_3352),
.B(n_3443),
.Y(n_3723)
);

A2O1A1Ixp33_ASAP7_75t_L g3724 ( 
.A1(n_3480),
.A2(n_3253),
.B(n_3415),
.C(n_3413),
.Y(n_3724)
);

OAI22xp33_ASAP7_75t_L g3725 ( 
.A1(n_3619),
.A2(n_3168),
.B1(n_3435),
.B2(n_3273),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_3471),
.B(n_3467),
.Y(n_3726)
);

BUFx6f_ASAP7_75t_L g3727 ( 
.A(n_3491),
.Y(n_3727)
);

AOI221xp5_ASAP7_75t_L g3728 ( 
.A1(n_3523),
.A2(n_3164),
.B1(n_3383),
.B2(n_3375),
.C(n_3276),
.Y(n_3728)
);

OAI221xp5_ASAP7_75t_L g3729 ( 
.A1(n_3558),
.A2(n_3328),
.B1(n_3276),
.B2(n_3301),
.C(n_3296),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_R g3730 ( 
.A(n_3483),
.B(n_3202),
.Y(n_3730)
);

AOI22xp33_ASAP7_75t_SL g3731 ( 
.A1(n_3699),
.A2(n_3338),
.B1(n_3341),
.B2(n_3390),
.Y(n_3731)
);

AO222x2_ASAP7_75t_L g3732 ( 
.A1(n_3645),
.A2(n_632),
.B1(n_635),
.B2(n_636),
.C1(n_637),
.C2(n_639),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3472),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_3581),
.B(n_3317),
.Y(n_3734)
);

OAI221xp5_ASAP7_75t_L g3735 ( 
.A1(n_3482),
.A2(n_3301),
.B1(n_3296),
.B2(n_3221),
.C(n_3193),
.Y(n_3735)
);

OR2x2_ASAP7_75t_L g3736 ( 
.A(n_3469),
.B(n_3193),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3478),
.B(n_3249),
.Y(n_3737)
);

AOI22xp33_ASAP7_75t_L g3738 ( 
.A1(n_3507),
.A2(n_3157),
.B1(n_3398),
.B2(n_3390),
.Y(n_3738)
);

OR2x2_ASAP7_75t_L g3739 ( 
.A(n_3499),
.B(n_3514),
.Y(n_3739)
);

OAI211xp5_ASAP7_75t_L g3740 ( 
.A1(n_3494),
.A2(n_3410),
.B(n_3277),
.C(n_3441),
.Y(n_3740)
);

AND2x2_ASAP7_75t_L g3741 ( 
.A(n_3468),
.B(n_3249),
.Y(n_3741)
);

AND2x4_ASAP7_75t_L g3742 ( 
.A(n_3615),
.B(n_3173),
.Y(n_3742)
);

AOI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3547),
.A2(n_3337),
.B(n_3329),
.Y(n_3743)
);

INVx2_ASAP7_75t_SL g3744 ( 
.A(n_3611),
.Y(n_3744)
);

AOI221xp5_ASAP7_75t_L g3745 ( 
.A1(n_3608),
.A2(n_3465),
.B1(n_3398),
.B2(n_3277),
.C(n_3373),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_L g3746 ( 
.A(n_3582),
.B(n_3317),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3473),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3565),
.B(n_3600),
.Y(n_3748)
);

AOI22xp33_ASAP7_75t_SL g3749 ( 
.A1(n_3525),
.A2(n_3341),
.B1(n_3373),
.B2(n_3323),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3562),
.A2(n_3323),
.B1(n_3159),
.B2(n_3179),
.Y(n_3750)
);

OAI22xp5_ASAP7_75t_L g3751 ( 
.A1(n_3700),
.A2(n_3303),
.B1(n_3173),
.B2(n_3366),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3663),
.A2(n_3159),
.B1(n_3179),
.B2(n_3221),
.Y(n_3752)
);

NAND3xp33_ASAP7_75t_L g3753 ( 
.A(n_3597),
.B(n_3215),
.C(n_3252),
.Y(n_3753)
);

AOI22xp33_ASAP7_75t_SL g3754 ( 
.A1(n_3621),
.A2(n_3303),
.B1(n_3397),
.B2(n_3254),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3513),
.Y(n_3755)
);

AOI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3511),
.A2(n_3215),
.B1(n_3252),
.B2(n_3272),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3585),
.B(n_3317),
.Y(n_3757)
);

BUFx3_ASAP7_75t_L g3758 ( 
.A(n_3500),
.Y(n_3758)
);

OAI222xp33_ASAP7_75t_L g3759 ( 
.A1(n_3700),
.A2(n_3280),
.B1(n_3333),
.B2(n_3462),
.C1(n_3350),
.C2(n_3355),
.Y(n_3759)
);

AND2x4_ASAP7_75t_L g3760 ( 
.A(n_3615),
.B(n_3339),
.Y(n_3760)
);

AOI22xp33_ASAP7_75t_L g3761 ( 
.A1(n_3470),
.A2(n_3272),
.B1(n_3282),
.B2(n_3293),
.Y(n_3761)
);

OAI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3490),
.A2(n_3339),
.B1(n_3293),
.B2(n_3462),
.Y(n_3762)
);

AO31x2_ASAP7_75t_L g3763 ( 
.A1(n_3530),
.A2(n_3389),
.A3(n_3178),
.B(n_3181),
.Y(n_3763)
);

AOI22xp33_ASAP7_75t_L g3764 ( 
.A1(n_3680),
.A2(n_3407),
.B1(n_3444),
.B2(n_3212),
.Y(n_3764)
);

AOI22xp33_ASAP7_75t_L g3765 ( 
.A1(n_3690),
.A2(n_3212),
.B1(n_3254),
.B2(n_3459),
.Y(n_3765)
);

AOI221xp5_ASAP7_75t_L g3766 ( 
.A1(n_3588),
.A2(n_3454),
.B1(n_3439),
.B2(n_3425),
.C(n_3458),
.Y(n_3766)
);

A2O1A1Ixp33_ASAP7_75t_L g3767 ( 
.A1(n_3616),
.A2(n_3357),
.B(n_3376),
.C(n_3365),
.Y(n_3767)
);

OAI221xp5_ASAP7_75t_L g3768 ( 
.A1(n_3529),
.A2(n_3389),
.B1(n_3425),
.B2(n_3439),
.C(n_3458),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3571),
.B(n_636),
.Y(n_3769)
);

INVx2_ASAP7_75t_SL g3770 ( 
.A(n_3510),
.Y(n_3770)
);

OAI211xp5_ASAP7_75t_L g3771 ( 
.A1(n_3709),
.A2(n_3466),
.B(n_3396),
.C(n_3403),
.Y(n_3771)
);

AOI22xp33_ASAP7_75t_L g3772 ( 
.A1(n_3520),
.A2(n_3234),
.B1(n_3381),
.B2(n_3379),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3475),
.Y(n_3773)
);

INVx3_ASAP7_75t_L g3774 ( 
.A(n_3656),
.Y(n_3774)
);

AOI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3579),
.A2(n_3248),
.B1(n_3454),
.B2(n_3450),
.Y(n_3775)
);

AOI22xp33_ASAP7_75t_L g3776 ( 
.A1(n_3578),
.A2(n_3449),
.B1(n_3395),
.B2(n_3242),
.Y(n_3776)
);

BUFx12f_ASAP7_75t_L g3777 ( 
.A(n_3498),
.Y(n_3777)
);

INVx1_ASAP7_75t_L g3778 ( 
.A(n_3486),
.Y(n_3778)
);

INVx1_ASAP7_75t_L g3779 ( 
.A(n_3515),
.Y(n_3779)
);

OAI221xp5_ASAP7_75t_L g3780 ( 
.A1(n_3660),
.A2(n_3458),
.B1(n_3447),
.B2(n_3437),
.C(n_3424),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3519),
.Y(n_3781)
);

AOI22xp33_ASAP7_75t_L g3782 ( 
.A1(n_3503),
.A2(n_3208),
.B1(n_3174),
.B2(n_3177),
.Y(n_3782)
);

OAI211xp5_ASAP7_75t_L g3783 ( 
.A1(n_3640),
.A2(n_3367),
.B(n_3351),
.C(n_3201),
.Y(n_3783)
);

AOI222xp33_ASAP7_75t_L g3784 ( 
.A1(n_3512),
.A2(n_3437),
.B1(n_3315),
.B2(n_3244),
.C1(n_3184),
.C2(n_3162),
.Y(n_3784)
);

OAI21xp33_ASAP7_75t_L g3785 ( 
.A1(n_3613),
.A2(n_3354),
.B(n_3311),
.Y(n_3785)
);

NAND2x1_ASAP7_75t_L g3786 ( 
.A(n_3673),
.B(n_3660),
.Y(n_3786)
);

INVx2_ASAP7_75t_SL g3787 ( 
.A(n_3654),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3521),
.Y(n_3788)
);

AND2x2_ASAP7_75t_L g3789 ( 
.A(n_3564),
.B(n_3437),
.Y(n_3789)
);

AND2x2_ASAP7_75t_L g3790 ( 
.A(n_3583),
.B(n_3447),
.Y(n_3790)
);

OAI22xp5_ASAP7_75t_L g3791 ( 
.A1(n_3502),
.A2(n_3447),
.B1(n_3348),
.B2(n_3161),
.Y(n_3791)
);

AOI22xp33_ASAP7_75t_L g3792 ( 
.A1(n_3503),
.A2(n_3643),
.B1(n_3572),
.B2(n_3542),
.Y(n_3792)
);

OAI221xp5_ASAP7_75t_L g3793 ( 
.A1(n_3574),
.A2(n_637),
.B1(n_640),
.B2(n_641),
.C(n_642),
.Y(n_3793)
);

BUFx6f_ASAP7_75t_L g3794 ( 
.A(n_3491),
.Y(n_3794)
);

OAI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3693),
.A2(n_3623),
.B(n_3625),
.Y(n_3795)
);

AOI22xp33_ASAP7_75t_SL g3796 ( 
.A1(n_3622),
.A2(n_3343),
.B1(n_3309),
.B2(n_3307),
.Y(n_3796)
);

OAI22xp33_ASAP7_75t_L g3797 ( 
.A1(n_3673),
.A2(n_3686),
.B1(n_3481),
.B2(n_3687),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3561),
.B(n_641),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3546),
.B(n_642),
.Y(n_3799)
);

AOI21xp33_ASAP7_75t_L g3800 ( 
.A1(n_3497),
.A2(n_3320),
.B(n_3182),
.Y(n_3800)
);

AOI22xp33_ASAP7_75t_SL g3801 ( 
.A1(n_3488),
.A2(n_3302),
.B1(n_644),
.B2(n_645),
.Y(n_3801)
);

AOI22xp33_ASAP7_75t_L g3802 ( 
.A1(n_3643),
.A2(n_643),
.B1(n_644),
.B2(n_645),
.Y(n_3802)
);

AOI22xp33_ASAP7_75t_L g3803 ( 
.A1(n_3631),
.A2(n_643),
.B1(n_646),
.B2(n_647),
.Y(n_3803)
);

BUFx2_ASAP7_75t_L g3804 ( 
.A(n_3577),
.Y(n_3804)
);

INVx5_ASAP7_75t_SL g3805 ( 
.A(n_3534),
.Y(n_3805)
);

AOI22xp33_ASAP7_75t_L g3806 ( 
.A1(n_3633),
.A2(n_647),
.B1(n_648),
.B2(n_649),
.Y(n_3806)
);

OR2x2_ASAP7_75t_L g3807 ( 
.A(n_3602),
.B(n_648),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3527),
.Y(n_3808)
);

OR2x6_ASAP7_75t_L g3809 ( 
.A(n_3543),
.B(n_650),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3522),
.Y(n_3810)
);

AOI21xp5_ASAP7_75t_L g3811 ( 
.A1(n_3477),
.A2(n_650),
.B(n_651),
.Y(n_3811)
);

OAI21xp5_ASAP7_75t_SL g3812 ( 
.A1(n_3485),
.A2(n_651),
.B(n_652),
.Y(n_3812)
);

OAI221xp5_ASAP7_75t_L g3813 ( 
.A1(n_3533),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.C(n_656),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3560),
.Y(n_3814)
);

AND2x2_ASAP7_75t_L g3815 ( 
.A(n_3568),
.B(n_3539),
.Y(n_3815)
);

AOI22xp33_ASAP7_75t_SL g3816 ( 
.A1(n_3488),
.A2(n_653),
.B1(n_654),
.B2(n_655),
.Y(n_3816)
);

NAND3xp33_ASAP7_75t_L g3817 ( 
.A(n_3614),
.B(n_657),
.C(n_658),
.Y(n_3817)
);

AOI22xp33_ASAP7_75t_SL g3818 ( 
.A1(n_3504),
.A2(n_660),
.B1(n_661),
.B2(n_662),
.Y(n_3818)
);

AOI21xp5_ASAP7_75t_L g3819 ( 
.A1(n_3516),
.A2(n_661),
.B(n_662),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3567),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3545),
.Y(n_3821)
);

AOI22xp33_ASAP7_75t_SL g3822 ( 
.A1(n_3504),
.A2(n_663),
.B1(n_664),
.B2(n_665),
.Y(n_3822)
);

AOI22xp33_ASAP7_75t_SL g3823 ( 
.A1(n_3591),
.A2(n_663),
.B1(n_665),
.B2(n_666),
.Y(n_3823)
);

AOI221xp5_ASAP7_75t_L g3824 ( 
.A1(n_3650),
.A2(n_667),
.B1(n_668),
.B2(n_669),
.C(n_671),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3544),
.Y(n_3825)
);

AND2x4_ASAP7_75t_L g3826 ( 
.A(n_3548),
.B(n_668),
.Y(n_3826)
);

OAI221xp5_ASAP7_75t_L g3827 ( 
.A1(n_3555),
.A2(n_669),
.B1(n_672),
.B2(n_673),
.C(n_675),
.Y(n_3827)
);

HB1xp67_ASAP7_75t_L g3828 ( 
.A(n_3691),
.Y(n_3828)
);

OAI22xp5_ASAP7_75t_L g3829 ( 
.A1(n_3635),
.A2(n_672),
.B1(n_673),
.B2(n_675),
.Y(n_3829)
);

INVx3_ASAP7_75t_L g3830 ( 
.A(n_3708),
.Y(n_3830)
);

OAI22xp5_ASAP7_75t_L g3831 ( 
.A1(n_3682),
.A2(n_676),
.B1(n_677),
.B2(n_678),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3484),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_3551),
.A2(n_679),
.B(n_681),
.Y(n_3833)
);

AND2x4_ASAP7_75t_L g3834 ( 
.A(n_3548),
.B(n_3505),
.Y(n_3834)
);

INVx1_ASAP7_75t_L g3835 ( 
.A(n_3662),
.Y(n_3835)
);

AOI22xp33_ASAP7_75t_L g3836 ( 
.A1(n_3664),
.A2(n_682),
.B1(n_683),
.B2(n_684),
.Y(n_3836)
);

CKINVDCx20_ASAP7_75t_R g3837 ( 
.A(n_3549),
.Y(n_3837)
);

AOI222xp33_ASAP7_75t_L g3838 ( 
.A1(n_3505),
.A2(n_682),
.B1(n_683),
.B2(n_684),
.C1(n_685),
.C2(n_686),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_SL g3839 ( 
.A1(n_3591),
.A2(n_686),
.B1(n_687),
.B2(n_688),
.Y(n_3839)
);

OAI22xp5_ASAP7_75t_L g3840 ( 
.A1(n_3675),
.A2(n_687),
.B1(n_690),
.B2(n_691),
.Y(n_3840)
);

OAI22xp5_ASAP7_75t_L g3841 ( 
.A1(n_3609),
.A2(n_3526),
.B1(n_3703),
.B2(n_3692),
.Y(n_3841)
);

AOI22xp33_ASAP7_75t_L g3842 ( 
.A1(n_3696),
.A2(n_691),
.B1(n_692),
.B2(n_693),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_L g3843 ( 
.A1(n_3684),
.A2(n_3677),
.B1(n_3678),
.B2(n_3676),
.Y(n_3843)
);

AOI221xp5_ASAP7_75t_L g3844 ( 
.A1(n_3655),
.A2(n_692),
.B1(n_694),
.B2(n_695),
.C(n_696),
.Y(n_3844)
);

AOI22xp33_ASAP7_75t_L g3845 ( 
.A1(n_3701),
.A2(n_695),
.B1(n_696),
.B2(n_697),
.Y(n_3845)
);

AO221x1_ASAP7_75t_L g3846 ( 
.A1(n_3589),
.A2(n_698),
.B1(n_700),
.B2(n_701),
.C(n_704),
.Y(n_3846)
);

OAI322xp33_ASAP7_75t_L g3847 ( 
.A1(n_3590),
.A2(n_698),
.A3(n_704),
.B1(n_705),
.B2(n_706),
.C1(n_707),
.C2(n_708),
.Y(n_3847)
);

AOI22xp33_ASAP7_75t_SL g3848 ( 
.A1(n_3594),
.A2(n_705),
.B1(n_706),
.B2(n_707),
.Y(n_3848)
);

AO31x2_ASAP7_75t_L g3849 ( 
.A1(n_3706),
.A2(n_709),
.A3(n_710),
.B(n_711),
.Y(n_3849)
);

AOI22xp33_ASAP7_75t_L g3850 ( 
.A1(n_3517),
.A2(n_712),
.B1(n_713),
.B2(n_714),
.Y(n_3850)
);

OAI22xp5_ASAP7_75t_L g3851 ( 
.A1(n_3704),
.A2(n_712),
.B1(n_714),
.B2(n_715),
.Y(n_3851)
);

AND2x2_ASAP7_75t_L g3852 ( 
.A(n_3518),
.B(n_802),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3607),
.Y(n_3853)
);

OAI211xp5_ASAP7_75t_L g3854 ( 
.A1(n_3659),
.A2(n_715),
.B(n_716),
.C(n_717),
.Y(n_3854)
);

AND2x2_ASAP7_75t_L g3855 ( 
.A(n_3624),
.B(n_801),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3632),
.B(n_801),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3569),
.B(n_3576),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3584),
.A2(n_716),
.B1(n_717),
.B2(n_718),
.Y(n_3858)
);

AOI22xp33_ASAP7_75t_SL g3859 ( 
.A1(n_3594),
.A2(n_719),
.B1(n_720),
.B2(n_722),
.Y(n_3859)
);

OAI22xp5_ASAP7_75t_L g3860 ( 
.A1(n_3618),
.A2(n_720),
.B1(n_722),
.B2(n_723),
.Y(n_3860)
);

AOI22xp33_ASAP7_75t_L g3861 ( 
.A1(n_3606),
.A2(n_723),
.B1(n_724),
.B2(n_725),
.Y(n_3861)
);

AOI22xp33_ASAP7_75t_L g3862 ( 
.A1(n_3552),
.A2(n_725),
.B1(n_726),
.B2(n_728),
.Y(n_3862)
);

AOI221xp5_ASAP7_75t_L g3863 ( 
.A1(n_3536),
.A2(n_726),
.B1(n_728),
.B2(n_730),
.C(n_731),
.Y(n_3863)
);

INVxp67_ASAP7_75t_L g3864 ( 
.A(n_3599),
.Y(n_3864)
);

AOI22xp33_ASAP7_75t_L g3865 ( 
.A1(n_3595),
.A2(n_730),
.B1(n_731),
.B2(n_733),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3679),
.B(n_3685),
.Y(n_3866)
);

CKINVDCx20_ASAP7_75t_R g3867 ( 
.A(n_3540),
.Y(n_3867)
);

OAI22xp33_ASAP7_75t_L g3868 ( 
.A1(n_3630),
.A2(n_800),
.B1(n_736),
.B2(n_737),
.Y(n_3868)
);

AOI22xp33_ASAP7_75t_SL g3869 ( 
.A1(n_3594),
.A2(n_735),
.B1(n_738),
.B2(n_739),
.Y(n_3869)
);

AOI22xp33_ASAP7_75t_L g3870 ( 
.A1(n_3573),
.A2(n_738),
.B1(n_739),
.B2(n_740),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3646),
.Y(n_3871)
);

INVx2_ASAP7_75t_SL g3872 ( 
.A(n_3669),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_3575),
.A2(n_740),
.B(n_741),
.Y(n_3873)
);

AND2x4_ASAP7_75t_L g3874 ( 
.A(n_3652),
.B(n_741),
.Y(n_3874)
);

OAI22xp5_ASAP7_75t_L g3875 ( 
.A1(n_3665),
.A2(n_742),
.B1(n_743),
.B2(n_744),
.Y(n_3875)
);

AOI22xp33_ASAP7_75t_SL g3876 ( 
.A1(n_3594),
.A2(n_743),
.B1(n_744),
.B2(n_745),
.Y(n_3876)
);

INVx3_ASAP7_75t_L g3877 ( 
.A(n_3708),
.Y(n_3877)
);

AOI221xp5_ASAP7_75t_L g3878 ( 
.A1(n_3628),
.A2(n_745),
.B1(n_746),
.B2(n_747),
.C(n_748),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3828),
.B(n_3697),
.Y(n_3879)
);

NAND3xp33_ASAP7_75t_L g3880 ( 
.A(n_3812),
.B(n_3613),
.C(n_3598),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_3714),
.Y(n_3881)
);

AO21x2_ASAP7_75t_L g3882 ( 
.A1(n_3743),
.A2(n_3617),
.B(n_3683),
.Y(n_3882)
);

AND2x2_ASAP7_75t_L g3883 ( 
.A(n_3737),
.B(n_3741),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3789),
.B(n_3639),
.Y(n_3884)
);

AND2x4_ASAP7_75t_L g3885 ( 
.A(n_3742),
.B(n_3657),
.Y(n_3885)
);

OAI22xp5_ASAP7_75t_L g3886 ( 
.A1(n_3710),
.A2(n_3666),
.B1(n_3670),
.B2(n_3672),
.Y(n_3886)
);

INVx2_ASAP7_75t_L g3887 ( 
.A(n_3755),
.Y(n_3887)
);

AND2x2_ASAP7_75t_L g3888 ( 
.A(n_3790),
.B(n_3667),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_L g3889 ( 
.A(n_3832),
.B(n_3605),
.Y(n_3889)
);

INVx2_ASAP7_75t_L g3890 ( 
.A(n_3810),
.Y(n_3890)
);

OR2x2_ASAP7_75t_L g3891 ( 
.A(n_3739),
.B(n_3736),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3814),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_L g3893 ( 
.A1(n_3846),
.A2(n_3537),
.B1(n_3702),
.B2(n_3496),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3734),
.B(n_3668),
.Y(n_3894)
);

NOR2x1_ASAP7_75t_L g3895 ( 
.A(n_3786),
.B(n_3674),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3820),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3821),
.Y(n_3897)
);

INVx1_ASAP7_75t_L g3898 ( 
.A(n_3733),
.Y(n_3898)
);

INVx3_ASAP7_75t_L g3899 ( 
.A(n_3760),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3747),
.Y(n_3900)
);

HB1xp67_ASAP7_75t_L g3901 ( 
.A(n_3722),
.Y(n_3901)
);

AND2x2_ASAP7_75t_L g3902 ( 
.A(n_3746),
.B(n_3689),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3748),
.B(n_3757),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3871),
.B(n_3695),
.Y(n_3904)
);

INVx2_ASAP7_75t_SL g3905 ( 
.A(n_3834),
.Y(n_3905)
);

BUFx3_ASAP7_75t_L g3906 ( 
.A(n_3758),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3825),
.B(n_3637),
.Y(n_3907)
);

INVx3_ASAP7_75t_L g3908 ( 
.A(n_3760),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_3773),
.Y(n_3909)
);

AND2x2_ASAP7_75t_L g3910 ( 
.A(n_3726),
.B(n_3495),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3720),
.A2(n_3550),
.B1(n_3489),
.B2(n_3487),
.Y(n_3911)
);

INVxp67_ASAP7_75t_SL g3912 ( 
.A(n_3751),
.Y(n_3912)
);

AND2x2_ASAP7_75t_L g3913 ( 
.A(n_3815),
.B(n_3570),
.Y(n_3913)
);

OR2x2_ASAP7_75t_L g3914 ( 
.A(n_3857),
.B(n_3647),
.Y(n_3914)
);

BUFx2_ASAP7_75t_L g3915 ( 
.A(n_3774),
.Y(n_3915)
);

AOI22xp33_ASAP7_75t_L g3916 ( 
.A1(n_3723),
.A2(n_3531),
.B1(n_3707),
.B2(n_3681),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3778),
.Y(n_3917)
);

AND2x2_ASAP7_75t_L g3918 ( 
.A(n_3779),
.B(n_3493),
.Y(n_3918)
);

OR2x2_ASAP7_75t_L g3919 ( 
.A(n_3781),
.B(n_3501),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3788),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3808),
.B(n_3756),
.Y(n_3921)
);

HB1xp67_ASAP7_75t_L g3922 ( 
.A(n_3874),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_L g3923 ( 
.A(n_3853),
.B(n_3835),
.Y(n_3923)
);

AND2x2_ASAP7_75t_L g3924 ( 
.A(n_3866),
.B(n_3580),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3849),
.Y(n_3925)
);

BUFx2_ASAP7_75t_L g3926 ( 
.A(n_3774),
.Y(n_3926)
);

AND2x2_ASAP7_75t_L g3927 ( 
.A(n_3752),
.B(n_3553),
.Y(n_3927)
);

INVx3_ASAP7_75t_L g3928 ( 
.A(n_3763),
.Y(n_3928)
);

INVx1_ASAP7_75t_L g3929 ( 
.A(n_3849),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3849),
.Y(n_3930)
);

BUFx2_ASAP7_75t_L g3931 ( 
.A(n_3730),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3750),
.B(n_3638),
.Y(n_3932)
);

AND2x2_ASAP7_75t_L g3933 ( 
.A(n_3784),
.B(n_3638),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3792),
.B(n_3698),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3735),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3785),
.Y(n_3936)
);

AND2x2_ASAP7_75t_L g3937 ( 
.A(n_3731),
.B(n_3638),
.Y(n_3937)
);

HB1xp67_ASAP7_75t_L g3938 ( 
.A(n_3874),
.Y(n_3938)
);

HB1xp67_ASAP7_75t_L g3939 ( 
.A(n_3864),
.Y(n_3939)
);

INVx2_ASAP7_75t_SL g3940 ( 
.A(n_3834),
.Y(n_3940)
);

INVx2_ASAP7_75t_L g3941 ( 
.A(n_3753),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3723),
.A2(n_3566),
.B1(n_3671),
.B2(n_3538),
.Y(n_3942)
);

AND2x2_ASAP7_75t_L g3943 ( 
.A(n_3749),
.B(n_3603),
.Y(n_3943)
);

INVx1_ASAP7_75t_L g3944 ( 
.A(n_3791),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3799),
.Y(n_3945)
);

BUFx2_ASAP7_75t_L g3946 ( 
.A(n_3804),
.Y(n_3946)
);

HB1xp67_ASAP7_75t_L g3947 ( 
.A(n_3770),
.Y(n_3947)
);

AND2x2_ASAP7_75t_L g3948 ( 
.A(n_3712),
.B(n_3641),
.Y(n_3948)
);

AOI22xp33_ASAP7_75t_L g3949 ( 
.A1(n_3880),
.A2(n_3718),
.B1(n_3797),
.B2(n_3795),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3881),
.Y(n_3950)
);

AND2x4_ASAP7_75t_L g3951 ( 
.A(n_3899),
.B(n_3908),
.Y(n_3951)
);

AND2x4_ASAP7_75t_L g3952 ( 
.A(n_3899),
.B(n_3830),
.Y(n_3952)
);

OR2x6_ASAP7_75t_L g3953 ( 
.A(n_3895),
.B(n_3717),
.Y(n_3953)
);

INVx2_ASAP7_75t_L g3954 ( 
.A(n_3881),
.Y(n_3954)
);

AO21x2_ASAP7_75t_L g3955 ( 
.A1(n_3936),
.A2(n_3783),
.B(n_3725),
.Y(n_3955)
);

OAI33xp33_ASAP7_75t_L g3956 ( 
.A1(n_3935),
.A2(n_3841),
.A3(n_3732),
.B1(n_3875),
.B2(n_3831),
.B3(n_3843),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3891),
.B(n_3541),
.Y(n_3957)
);

AND2x2_ASAP7_75t_L g3958 ( 
.A(n_3903),
.B(n_3719),
.Y(n_3958)
);

BUFx3_ASAP7_75t_L g3959 ( 
.A(n_3906),
.Y(n_3959)
);

OAI211xp5_ASAP7_75t_L g3960 ( 
.A1(n_3931),
.A2(n_3838),
.B(n_3724),
.C(n_3848),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_3946),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3898),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_3898),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_3900),
.Y(n_3964)
);

NOR3xp33_ASAP7_75t_L g3965 ( 
.A(n_3935),
.B(n_3769),
.C(n_3817),
.Y(n_3965)
);

INVx2_ASAP7_75t_L g3966 ( 
.A(n_3887),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3900),
.Y(n_3967)
);

OA222x2_ASAP7_75t_L g3968 ( 
.A1(n_3906),
.A2(n_3809),
.B1(n_3532),
.B2(n_3807),
.C1(n_3830),
.C2(n_3877),
.Y(n_3968)
);

OAI31xp33_ASAP7_75t_L g3969 ( 
.A1(n_3880),
.A2(n_3826),
.A3(n_3829),
.B(n_3780),
.Y(n_3969)
);

A2O1A1Ixp33_ASAP7_75t_L g3970 ( 
.A1(n_3931),
.A2(n_3826),
.B(n_3717),
.C(n_3744),
.Y(n_3970)
);

AOI22xp5_ASAP7_75t_L g3971 ( 
.A1(n_3934),
.A2(n_3809),
.B1(n_3839),
.B2(n_3823),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_L g3972 ( 
.A(n_3918),
.B(n_3761),
.Y(n_3972)
);

OR2x2_ASAP7_75t_L g3973 ( 
.A(n_3891),
.B(n_3563),
.Y(n_3973)
);

OAI221xp5_ASAP7_75t_L g3974 ( 
.A1(n_3912),
.A2(n_3721),
.B1(n_3713),
.B2(n_3711),
.C(n_3859),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3909),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3909),
.Y(n_3976)
);

INVx1_ASAP7_75t_L g3977 ( 
.A(n_3917),
.Y(n_3977)
);

AO21x2_ASAP7_75t_L g3978 ( 
.A1(n_3936),
.A2(n_3800),
.B(n_3740),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3917),
.Y(n_3979)
);

NAND3xp33_ASAP7_75t_L g3980 ( 
.A(n_3941),
.B(n_3876),
.C(n_3869),
.Y(n_3980)
);

AOI211xp5_ASAP7_75t_L g3981 ( 
.A1(n_3946),
.A2(n_3587),
.B(n_3847),
.C(n_3762),
.Y(n_3981)
);

OA21x2_ASAP7_75t_L g3982 ( 
.A1(n_3941),
.A2(n_3759),
.B(n_3745),
.Y(n_3982)
);

OAI221xp5_ASAP7_75t_L g3983 ( 
.A1(n_3942),
.A2(n_3822),
.B1(n_3818),
.B2(n_3816),
.C(n_3738),
.Y(n_3983)
);

OAI221xp5_ASAP7_75t_L g3984 ( 
.A1(n_3916),
.A2(n_3715),
.B1(n_3802),
.B2(n_3850),
.C(n_3766),
.Y(n_3984)
);

NOR2x1_ASAP7_75t_L g3985 ( 
.A(n_3895),
.B(n_3837),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_3920),
.Y(n_3986)
);

BUFx3_ASAP7_75t_L g3987 ( 
.A(n_3947),
.Y(n_3987)
);

HB1xp67_ASAP7_75t_L g3988 ( 
.A(n_3901),
.Y(n_3988)
);

OAI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3905),
.A2(n_3729),
.B1(n_3768),
.B2(n_3658),
.Y(n_3989)
);

AOI22xp33_ASAP7_75t_SL g3990 ( 
.A1(n_3922),
.A2(n_3805),
.B1(n_3658),
.B2(n_3629),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_L g3991 ( 
.A(n_3918),
.B(n_3728),
.Y(n_3991)
);

OR2x2_ASAP7_75t_L g3992 ( 
.A(n_3879),
.B(n_3914),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3920),
.Y(n_3993)
);

INVx1_ASAP7_75t_L g3994 ( 
.A(n_3897),
.Y(n_3994)
);

INVx2_ASAP7_75t_L g3995 ( 
.A(n_3887),
.Y(n_3995)
);

NOR4xp25_ASAP7_75t_SL g3996 ( 
.A(n_3915),
.B(n_3604),
.C(n_3627),
.D(n_3648),
.Y(n_3996)
);

AOI221xp5_ASAP7_75t_SL g3997 ( 
.A1(n_3933),
.A2(n_3798),
.B1(n_3852),
.B2(n_3819),
.C(n_3793),
.Y(n_3997)
);

NOR2xp33_ASAP7_75t_L g3998 ( 
.A(n_3939),
.B(n_3872),
.Y(n_3998)
);

AOI22xp33_ASAP7_75t_L g3999 ( 
.A1(n_3903),
.A2(n_3813),
.B1(n_3827),
.B2(n_3844),
.Y(n_3999)
);

NOR2xp33_ASAP7_75t_R g4000 ( 
.A(n_3905),
.B(n_3867),
.Y(n_4000)
);

OAI211xp5_ASAP7_75t_SL g4001 ( 
.A1(n_3911),
.A2(n_3878),
.B(n_3865),
.C(n_3863),
.Y(n_4001)
);

INVx3_ASAP7_75t_L g4002 ( 
.A(n_3899),
.Y(n_4002)
);

OAI211xp5_ASAP7_75t_L g4003 ( 
.A1(n_3944),
.A2(n_3764),
.B(n_3862),
.C(n_3858),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3883),
.B(n_3877),
.Y(n_4004)
);

AOI211xp5_ASAP7_75t_L g4005 ( 
.A1(n_3938),
.A2(n_3868),
.B(n_3854),
.C(n_3771),
.Y(n_4005)
);

AOI21xp5_ASAP7_75t_L g4006 ( 
.A1(n_3933),
.A2(n_3767),
.B(n_3886),
.Y(n_4006)
);

INVx2_ASAP7_75t_L g4007 ( 
.A(n_3890),
.Y(n_4007)
);

INVx1_ASAP7_75t_L g4008 ( 
.A(n_3897),
.Y(n_4008)
);

AND2x2_ASAP7_75t_L g4009 ( 
.A(n_3883),
.B(n_3556),
.Y(n_4009)
);

AOI221xp5_ASAP7_75t_SL g4010 ( 
.A1(n_3907),
.A2(n_3833),
.B1(n_3873),
.B2(n_3824),
.C(n_3861),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3913),
.B(n_3556),
.Y(n_4011)
);

BUFx2_ASAP7_75t_L g4012 ( 
.A(n_3940),
.Y(n_4012)
);

OAI22xp5_ASAP7_75t_L g4013 ( 
.A1(n_3940),
.A2(n_3805),
.B1(n_3801),
.B2(n_3754),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_3902),
.B(n_3855),
.Y(n_4014)
);

OAI221xp5_ASAP7_75t_L g4015 ( 
.A1(n_3893),
.A2(n_3775),
.B1(n_3870),
.B2(n_3716),
.C(n_3806),
.Y(n_4015)
);

BUFx2_ASAP7_75t_L g4016 ( 
.A(n_3908),
.Y(n_4016)
);

NAND4xp25_ASAP7_75t_L g4017 ( 
.A(n_3949),
.B(n_3911),
.C(n_3943),
.D(n_3944),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_L g4018 ( 
.A(n_3991),
.B(n_3921),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_L g4019 ( 
.A(n_3988),
.B(n_3921),
.Y(n_4019)
);

AND2x2_ASAP7_75t_L g4020 ( 
.A(n_3958),
.B(n_3913),
.Y(n_4020)
);

HB1xp67_ASAP7_75t_L g4021 ( 
.A(n_3961),
.Y(n_4021)
);

OR2x2_ASAP7_75t_L g4022 ( 
.A(n_3992),
.B(n_3879),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3950),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3994),
.Y(n_4024)
);

AND2x2_ASAP7_75t_L g4025 ( 
.A(n_4004),
.B(n_4011),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_4008),
.Y(n_4026)
);

AND2x2_ASAP7_75t_L g4027 ( 
.A(n_4009),
.B(n_3910),
.Y(n_4027)
);

INVx1_ASAP7_75t_SL g4028 ( 
.A(n_4000),
.Y(n_4028)
);

HB1xp67_ASAP7_75t_L g4029 ( 
.A(n_3959),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3953),
.B(n_3787),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_4012),
.B(n_3910),
.Y(n_4031)
);

INVx1_ASAP7_75t_L g4032 ( 
.A(n_3986),
.Y(n_4032)
);

AND2x2_ASAP7_75t_L g4033 ( 
.A(n_4016),
.B(n_3957),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3973),
.B(n_3951),
.Y(n_4034)
);

AND2x2_ASAP7_75t_L g4035 ( 
.A(n_3951),
.B(n_3937),
.Y(n_4035)
);

NAND2x1_ASAP7_75t_SL g4036 ( 
.A(n_3985),
.B(n_3937),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3954),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_4002),
.B(n_3924),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_4006),
.B(n_3902),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_4002),
.B(n_3924),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3966),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3972),
.B(n_3888),
.Y(n_4042)
);

AND2x2_ASAP7_75t_L g4043 ( 
.A(n_3987),
.B(n_3888),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_4014),
.B(n_3943),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3993),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_3995),
.B(n_3884),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3962),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3963),
.B(n_3894),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_L g4049 ( 
.A(n_3964),
.B(n_3894),
.Y(n_4049)
);

INVx1_ASAP7_75t_SL g4050 ( 
.A(n_3953),
.Y(n_4050)
);

AND2x4_ASAP7_75t_SL g4051 ( 
.A(n_3953),
.B(n_3908),
.Y(n_4051)
);

BUFx12f_ASAP7_75t_L g4052 ( 
.A(n_3952),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_3967),
.B(n_3927),
.Y(n_4053)
);

NOR2xp67_ASAP7_75t_L g4054 ( 
.A(n_4013),
.B(n_3948),
.Y(n_4054)
);

BUFx2_ASAP7_75t_SL g4055 ( 
.A(n_3971),
.Y(n_4055)
);

INVx2_ASAP7_75t_L g4056 ( 
.A(n_4007),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3952),
.B(n_3884),
.Y(n_4057)
);

INVx1_ASAP7_75t_L g4058 ( 
.A(n_3975),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3976),
.B(n_3927),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_SL g4060 ( 
.A(n_3969),
.B(n_3915),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3955),
.B(n_3932),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3955),
.B(n_3932),
.Y(n_4062)
);

OR2x2_ASAP7_75t_L g4063 ( 
.A(n_3977),
.B(n_3914),
.Y(n_4063)
);

OR2x2_ASAP7_75t_L g4064 ( 
.A(n_3979),
.B(n_3919),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_3982),
.B(n_3926),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3982),
.Y(n_4066)
);

AND2x4_ASAP7_75t_SL g4067 ( 
.A(n_3998),
.B(n_3885),
.Y(n_4067)
);

INVx2_ASAP7_75t_SL g4068 ( 
.A(n_3978),
.Y(n_4068)
);

OR2x2_ASAP7_75t_L g4069 ( 
.A(n_3978),
.B(n_3919),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3970),
.Y(n_4070)
);

INVx2_ASAP7_75t_L g4071 ( 
.A(n_3974),
.Y(n_4071)
);

OR2x2_ASAP7_75t_L g4072 ( 
.A(n_3969),
.B(n_3889),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3968),
.B(n_3926),
.Y(n_4073)
);

OR2x2_ASAP7_75t_L g4074 ( 
.A(n_3989),
.B(n_3890),
.Y(n_4074)
);

OR2x2_ASAP7_75t_L g4075 ( 
.A(n_4022),
.B(n_4048),
.Y(n_4075)
);

NOR2xp33_ASAP7_75t_L g4076 ( 
.A(n_4028),
.B(n_3956),
.Y(n_4076)
);

INVx2_ASAP7_75t_L g4077 ( 
.A(n_4023),
.Y(n_4077)
);

OAI22xp5_ASAP7_75t_L g4078 ( 
.A1(n_4054),
.A2(n_3990),
.B1(n_3981),
.B2(n_3971),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_4044),
.B(n_4071),
.Y(n_4079)
);

INVx2_ASAP7_75t_L g4080 ( 
.A(n_4023),
.Y(n_4080)
);

INVx3_ASAP7_75t_SL g4081 ( 
.A(n_4051),
.Y(n_4081)
);

AOI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_4055),
.A2(n_3960),
.B1(n_3965),
.B2(n_3997),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_4044),
.B(n_3948),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_4050),
.B(n_3968),
.Y(n_4084)
);

INVx1_ASAP7_75t_L g4085 ( 
.A(n_4064),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_4071),
.B(n_3904),
.Y(n_4086)
);

NAND2xp33_ASAP7_75t_SL g4087 ( 
.A(n_4073),
.B(n_3996),
.Y(n_4087)
);

INVx2_ASAP7_75t_SL g4088 ( 
.A(n_4051),
.Y(n_4088)
);

OR2x2_ASAP7_75t_L g4089 ( 
.A(n_4022),
.B(n_3892),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_4072),
.B(n_3904),
.Y(n_4090)
);

INVx1_ASAP7_75t_L g4091 ( 
.A(n_4064),
.Y(n_4091)
);

AND2x4_ASAP7_75t_L g4092 ( 
.A(n_4073),
.B(n_3945),
.Y(n_4092)
);

OR2x2_ASAP7_75t_L g4093 ( 
.A(n_4049),
.B(n_3892),
.Y(n_4093)
);

OR2x6_ASAP7_75t_L g4094 ( 
.A(n_4055),
.B(n_3980),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_4072),
.B(n_3945),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_4039),
.B(n_3925),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_4063),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_4063),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_4035),
.B(n_3885),
.Y(n_4099)
);

NOR2xp33_ASAP7_75t_L g4100 ( 
.A(n_4070),
.B(n_3777),
.Y(n_4100)
);

HB1xp67_ASAP7_75t_L g4101 ( 
.A(n_4021),
.Y(n_4101)
);

INVx1_ASAP7_75t_L g4102 ( 
.A(n_4024),
.Y(n_4102)
);

AOI32xp33_ASAP7_75t_L g4103 ( 
.A1(n_4060),
.A2(n_3981),
.A3(n_4005),
.B1(n_3983),
.B2(n_3984),
.Y(n_4103)
);

AND2x2_ASAP7_75t_L g4104 ( 
.A(n_4035),
.B(n_4031),
.Y(n_4104)
);

NOR2x1_ASAP7_75t_SL g4105 ( 
.A(n_4052),
.B(n_3980),
.Y(n_4105)
);

NAND2x1p5_ASAP7_75t_L g4106 ( 
.A(n_4030),
.B(n_3727),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4026),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_4018),
.B(n_3925),
.Y(n_4108)
);

INVxp67_ASAP7_75t_L g4109 ( 
.A(n_4029),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4047),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_4031),
.B(n_3885),
.Y(n_4111)
);

OAI21xp33_ASAP7_75t_L g4112 ( 
.A1(n_4017),
.A2(n_4003),
.B(n_4005),
.Y(n_4112)
);

CKINVDCx5p33_ASAP7_75t_R g4113 ( 
.A(n_4100),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4081),
.B(n_4067),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_4101),
.Y(n_4115)
);

INVx5_ASAP7_75t_L g4116 ( 
.A(n_4094),
.Y(n_4116)
);

NOR2xp33_ASAP7_75t_L g4117 ( 
.A(n_4112),
.B(n_4076),
.Y(n_4117)
);

INVx4_ASAP7_75t_L g4118 ( 
.A(n_4094),
.Y(n_4118)
);

AND2x2_ASAP7_75t_L g4119 ( 
.A(n_4092),
.B(n_4065),
.Y(n_4119)
);

CKINVDCx5p33_ASAP7_75t_R g4120 ( 
.A(n_4094),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4092),
.B(n_4065),
.Y(n_4121)
);

INVx2_ASAP7_75t_L g4122 ( 
.A(n_4077),
.Y(n_4122)
);

NAND4xp25_ASAP7_75t_L g4123 ( 
.A(n_4103),
.B(n_3999),
.C(n_4015),
.D(n_4001),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_4080),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4095),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_4084),
.B(n_4066),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_4086),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4088),
.B(n_4067),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_4079),
.B(n_4061),
.Y(n_4129)
);

INVx2_ASAP7_75t_SL g4130 ( 
.A(n_4106),
.Y(n_4130)
);

INVx2_ASAP7_75t_L g4131 ( 
.A(n_4089),
.Y(n_4131)
);

OR2x2_ASAP7_75t_L g4132 ( 
.A(n_4090),
.B(n_4074),
.Y(n_4132)
);

OAI22xp5_ASAP7_75t_L g4133 ( 
.A1(n_4078),
.A2(n_4052),
.B1(n_4074),
.B2(n_4066),
.Y(n_4133)
);

AND2x4_ASAP7_75t_L g4134 ( 
.A(n_4105),
.B(n_4061),
.Y(n_4134)
);

OAI22xp5_ASAP7_75t_L g4135 ( 
.A1(n_4082),
.A2(n_4062),
.B1(n_4019),
.B2(n_4033),
.Y(n_4135)
);

OR2x2_ASAP7_75t_L g4136 ( 
.A(n_4108),
.B(n_4053),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4104),
.B(n_4062),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4085),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4091),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_4075),
.Y(n_4140)
);

NOR4xp75_ASAP7_75t_L g4141 ( 
.A(n_4112),
.B(n_4036),
.C(n_4068),
.D(n_4059),
.Y(n_4141)
);

INVx2_ASAP7_75t_L g4142 ( 
.A(n_4093),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_4111),
.B(n_4109),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4097),
.Y(n_4144)
);

CKINVDCx16_ASAP7_75t_R g4145 ( 
.A(n_4082),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_L g4146 ( 
.A(n_4103),
.B(n_4042),
.Y(n_4146)
);

HB1xp67_ASAP7_75t_L g4147 ( 
.A(n_4102),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_4098),
.Y(n_4148)
);

HB1xp67_ASAP7_75t_L g4149 ( 
.A(n_4107),
.Y(n_4149)
);

NOR2x1_ASAP7_75t_L g4150 ( 
.A(n_4096),
.B(n_4069),
.Y(n_4150)
);

HB1xp67_ASAP7_75t_L g4151 ( 
.A(n_4110),
.Y(n_4151)
);

INVx2_ASAP7_75t_SL g4152 ( 
.A(n_4114),
.Y(n_4152)
);

AOI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_4123),
.A2(n_4087),
.B(n_4069),
.Y(n_4153)
);

INVxp67_ASAP7_75t_SL g4154 ( 
.A(n_4117),
.Y(n_4154)
);

HB1xp67_ASAP7_75t_L g4155 ( 
.A(n_4115),
.Y(n_4155)
);

AOI21xp5_ASAP7_75t_L g4156 ( 
.A1(n_4116),
.A2(n_4068),
.B(n_4083),
.Y(n_4156)
);

OR2x2_ASAP7_75t_L g4157 ( 
.A(n_4140),
.B(n_4033),
.Y(n_4157)
);

OAI21xp5_ASAP7_75t_SL g4158 ( 
.A1(n_4117),
.A2(n_3836),
.B(n_3803),
.Y(n_4158)
);

OR2x2_ASAP7_75t_L g4159 ( 
.A(n_4127),
.B(n_4032),
.Y(n_4159)
);

NAND2xp5_ASAP7_75t_L g4160 ( 
.A(n_4145),
.B(n_4042),
.Y(n_4160)
);

INVxp67_ASAP7_75t_L g4161 ( 
.A(n_4120),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4147),
.Y(n_4162)
);

NOR2xp33_ASAP7_75t_L g4163 ( 
.A(n_4113),
.B(n_3593),
.Y(n_4163)
);

CKINVDCx20_ASAP7_75t_R g4164 ( 
.A(n_4113),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4149),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_4118),
.B(n_3601),
.Y(n_4166)
);

OR2x2_ASAP7_75t_L g4167 ( 
.A(n_4132),
.B(n_4032),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_4151),
.Y(n_4168)
);

INVxp67_ASAP7_75t_SL g4169 ( 
.A(n_4118),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4143),
.Y(n_4170)
);

OAI22xp5_ASAP7_75t_L g4171 ( 
.A1(n_4116),
.A2(n_4043),
.B1(n_4034),
.B2(n_4099),
.Y(n_4171)
);

OR2x2_ASAP7_75t_L g4172 ( 
.A(n_4125),
.B(n_4045),
.Y(n_4172)
);

OAI31xp33_ASAP7_75t_L g4173 ( 
.A1(n_4133),
.A2(n_4043),
.A3(n_4034),
.B(n_4040),
.Y(n_4173)
);

AOI21xp5_ASAP7_75t_L g4174 ( 
.A1(n_4116),
.A2(n_3508),
.B(n_4038),
.Y(n_4174)
);

AOI322xp5_ASAP7_75t_L g4175 ( 
.A1(n_4146),
.A2(n_4020),
.A3(n_4038),
.B1(n_4040),
.B2(n_4027),
.C1(n_4046),
.C2(n_4057),
.Y(n_4175)
);

AOI221xp5_ASAP7_75t_L g4176 ( 
.A1(n_4118),
.A2(n_4058),
.B1(n_4045),
.B2(n_3923),
.C(n_4010),
.Y(n_4176)
);

INVx1_ASAP7_75t_L g4177 ( 
.A(n_4143),
.Y(n_4177)
);

BUFx2_ASAP7_75t_SL g4178 ( 
.A(n_4116),
.Y(n_4178)
);

AND2x4_ASAP7_75t_L g4179 ( 
.A(n_4128),
.B(n_4130),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4138),
.Y(n_4180)
);

INVx2_ASAP7_75t_L g4181 ( 
.A(n_4179),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_4155),
.Y(n_4182)
);

OAI22xp33_ASAP7_75t_L g4183 ( 
.A1(n_4160),
.A2(n_4120),
.B1(n_4135),
.B2(n_4134),
.Y(n_4183)
);

AOI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_4161),
.A2(n_4134),
.B1(n_4126),
.B2(n_4129),
.Y(n_4184)
);

INVx2_ASAP7_75t_SL g4185 ( 
.A(n_4179),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_4154),
.B(n_4126),
.Y(n_4186)
);

AOI322xp5_ASAP7_75t_L g4187 ( 
.A1(n_4169),
.A2(n_4166),
.A3(n_4176),
.B1(n_4177),
.B2(n_4170),
.C1(n_4152),
.C2(n_4134),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4157),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_4153),
.B(n_4162),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4165),
.Y(n_4190)
);

INVx1_ASAP7_75t_L g4191 ( 
.A(n_4168),
.Y(n_4191)
);

INVx1_ASAP7_75t_SL g4192 ( 
.A(n_4164),
.Y(n_4192)
);

AOI22xp5_ASAP7_75t_L g4193 ( 
.A1(n_4178),
.A2(n_4130),
.B1(n_4119),
.B2(n_4121),
.Y(n_4193)
);

OAI32xp33_ASAP7_75t_L g4194 ( 
.A1(n_4171),
.A2(n_4141),
.A3(n_4148),
.B1(n_4144),
.B2(n_4139),
.Y(n_4194)
);

INVxp67_ASAP7_75t_L g4195 ( 
.A(n_4163),
.Y(n_4195)
);

OR2x2_ASAP7_75t_L g4196 ( 
.A(n_4167),
.B(n_4142),
.Y(n_4196)
);

NOR2xp33_ASAP7_75t_L g4197 ( 
.A(n_4174),
.B(n_4142),
.Y(n_4197)
);

OAI22xp33_ASAP7_75t_L g4198 ( 
.A1(n_4156),
.A2(n_4119),
.B1(n_4121),
.B2(n_4150),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_4158),
.B(n_4137),
.Y(n_4199)
);

NOR3xp33_ASAP7_75t_SL g4200 ( 
.A(n_4173),
.B(n_3851),
.C(n_3860),
.Y(n_4200)
);

OAI21xp33_ASAP7_75t_L g4201 ( 
.A1(n_4175),
.A2(n_4036),
.B(n_4137),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4159),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4172),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4186),
.Y(n_4204)
);

OAI21xp5_ASAP7_75t_SL g4205 ( 
.A1(n_4187),
.A2(n_4175),
.B(n_4180),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_4192),
.B(n_4131),
.Y(n_4206)
);

HB1xp67_ASAP7_75t_L g4207 ( 
.A(n_4182),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4196),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4181),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4185),
.B(n_4131),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_4195),
.B(n_4122),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_4183),
.B(n_4122),
.Y(n_4212)
);

AOI21xp5_ASAP7_75t_L g4213 ( 
.A1(n_4189),
.A2(n_4124),
.B(n_4136),
.Y(n_4213)
);

NOR4xp25_ASAP7_75t_SL g4214 ( 
.A(n_4190),
.B(n_3610),
.C(n_3930),
.D(n_3929),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4188),
.Y(n_4215)
);

AND2x2_ASAP7_75t_L g4216 ( 
.A(n_4197),
.B(n_4020),
.Y(n_4216)
);

INVx1_ASAP7_75t_SL g4217 ( 
.A(n_4191),
.Y(n_4217)
);

AOI22x1_ASAP7_75t_L g4218 ( 
.A1(n_4202),
.A2(n_4124),
.B1(n_3612),
.B2(n_3811),
.Y(n_4218)
);

AOI22xp5_ASAP7_75t_L g4219 ( 
.A1(n_4184),
.A2(n_4057),
.B1(n_3882),
.B2(n_4027),
.Y(n_4219)
);

OR2x2_ASAP7_75t_L g4220 ( 
.A(n_4203),
.B(n_4025),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_4187),
.B(n_4025),
.Y(n_4221)
);

NAND2xp5_ASAP7_75t_L g4222 ( 
.A(n_4199),
.B(n_4037),
.Y(n_4222)
);

XOR2xp5_ASAP7_75t_L g4223 ( 
.A(n_4193),
.B(n_3794),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4200),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4224),
.B(n_4216),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_SL g4226 ( 
.A(n_4209),
.B(n_4198),
.Y(n_4226)
);

NAND2xp5_ASAP7_75t_L g4227 ( 
.A(n_4205),
.B(n_4201),
.Y(n_4227)
);

NOR2x1_ASAP7_75t_L g4228 ( 
.A(n_4206),
.B(n_4194),
.Y(n_4228)
);

NAND3xp33_ASAP7_75t_SL g4229 ( 
.A(n_4217),
.B(n_3845),
.C(n_3842),
.Y(n_4229)
);

NOR3xp33_ASAP7_75t_L g4230 ( 
.A(n_4212),
.B(n_3612),
.C(n_3840),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4210),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_4221),
.B(n_4208),
.Y(n_4232)
);

NOR2xp67_ASAP7_75t_L g4233 ( 
.A(n_4207),
.B(n_746),
.Y(n_4233)
);

INVxp67_ASAP7_75t_L g4234 ( 
.A(n_4211),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_4204),
.B(n_4046),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_4223),
.B(n_4037),
.Y(n_4236)
);

XNOR2x1_ASAP7_75t_L g4237 ( 
.A(n_4217),
.B(n_3649),
.Y(n_4237)
);

OAI22xp5_ASAP7_75t_L g4238 ( 
.A1(n_4219),
.A2(n_4222),
.B1(n_4220),
.B2(n_4215),
.Y(n_4238)
);

CKINVDCx20_ASAP7_75t_R g4239 ( 
.A(n_4222),
.Y(n_4239)
);

INVxp67_ASAP7_75t_L g4240 ( 
.A(n_4225),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4231),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_4227),
.A2(n_4213),
.B(n_4214),
.Y(n_4242)
);

INVx1_ASAP7_75t_L g4243 ( 
.A(n_4235),
.Y(n_4243)
);

NAND2xp5_ASAP7_75t_SL g4244 ( 
.A(n_4228),
.B(n_4218),
.Y(n_4244)
);

INVx3_ASAP7_75t_L g4245 ( 
.A(n_4236),
.Y(n_4245)
);

OAI221xp5_ASAP7_75t_L g4246 ( 
.A1(n_4226),
.A2(n_3610),
.B1(n_3661),
.B2(n_3642),
.C(n_3653),
.Y(n_4246)
);

XOR2x2_ASAP7_75t_L g4247 ( 
.A(n_4232),
.B(n_3856),
.Y(n_4247)
);

OAI21xp5_ASAP7_75t_L g4248 ( 
.A1(n_4234),
.A2(n_4239),
.B(n_4233),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4237),
.A2(n_4056),
.B1(n_4041),
.B2(n_3928),
.Y(n_4249)
);

BUFx2_ASAP7_75t_L g4250 ( 
.A(n_4238),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_L g4251 ( 
.A(n_4250),
.B(n_4230),
.Y(n_4251)
);

AOI221xp5_ASAP7_75t_L g4252 ( 
.A1(n_4242),
.A2(n_4229),
.B1(n_3636),
.B2(n_3644),
.C(n_3694),
.Y(n_4252)
);

NOR2x1_ASAP7_75t_L g4253 ( 
.A(n_4244),
.B(n_3634),
.Y(n_4253)
);

AND2x4_ASAP7_75t_L g4254 ( 
.A(n_4245),
.B(n_4041),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4245),
.Y(n_4255)
);

INVx2_ASAP7_75t_L g4256 ( 
.A(n_4254),
.Y(n_4256)
);

AND2x2_ASAP7_75t_L g4257 ( 
.A(n_4255),
.B(n_4240),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_4251),
.A2(n_4248),
.B(n_4241),
.Y(n_4258)
);

NOR2x1_ASAP7_75t_L g4259 ( 
.A(n_4253),
.B(n_4243),
.Y(n_4259)
);

O2A1O1Ixp33_ASAP7_75t_L g4260 ( 
.A1(n_4252),
.A2(n_4246),
.B(n_4249),
.C(n_4247),
.Y(n_4260)
);

HB1xp67_ASAP7_75t_L g4261 ( 
.A(n_4256),
.Y(n_4261)
);

NAND5xp2_ASAP7_75t_L g4262 ( 
.A(n_4258),
.B(n_3592),
.C(n_3524),
.D(n_3765),
.E(n_3772),
.Y(n_4262)
);

AOI211x1_ASAP7_75t_L g4263 ( 
.A1(n_4257),
.A2(n_3930),
.B(n_3929),
.C(n_3896),
.Y(n_4263)
);

NAND5xp2_ASAP7_75t_L g4264 ( 
.A(n_4260),
.B(n_3554),
.C(n_3776),
.D(n_751),
.E(n_752),
.Y(n_4264)
);

XOR2xp5_ASAP7_75t_L g4265 ( 
.A(n_4261),
.B(n_4259),
.Y(n_4265)
);

AOI22xp5_ASAP7_75t_L g4266 ( 
.A1(n_4264),
.A2(n_3491),
.B1(n_3506),
.B2(n_3596),
.Y(n_4266)
);

NAND2x1_ASAP7_75t_L g4267 ( 
.A(n_4266),
.B(n_4263),
.Y(n_4267)
);

AND2x2_ASAP7_75t_L g4268 ( 
.A(n_4267),
.B(n_4265),
.Y(n_4268)
);

OAI22x1_ASAP7_75t_L g4269 ( 
.A1(n_4267),
.A2(n_4262),
.B1(n_3688),
.B2(n_3705),
.Y(n_4269)
);

CKINVDCx20_ASAP7_75t_R g4270 ( 
.A(n_4268),
.Y(n_4270)
);

AOI21xp33_ASAP7_75t_L g4271 ( 
.A1(n_4270),
.A2(n_4269),
.B(n_750),
.Y(n_4271)
);

O2A1O1Ixp33_ASAP7_75t_L g4272 ( 
.A1(n_4271),
.A2(n_749),
.B(n_750),
.C(n_751),
.Y(n_4272)
);

XOR2x2_ASAP7_75t_L g4273 ( 
.A(n_4272),
.B(n_749),
.Y(n_4273)
);

OAI221xp5_ASAP7_75t_R g4274 ( 
.A1(n_4273),
.A2(n_3796),
.B1(n_3782),
.B2(n_3794),
.C(n_754),
.Y(n_4274)
);

AOI211xp5_ASAP7_75t_L g4275 ( 
.A1(n_4274),
.A2(n_3506),
.B(n_3596),
.C(n_3794),
.Y(n_4275)
);


endmodule