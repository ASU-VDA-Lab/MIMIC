module real_aes_17434_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_1403, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_1403;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1145;
wire n_645;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_249;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_1085;
wire n_276;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_0), .A2(n_60), .B1(n_686), .B2(n_691), .Y(n_690) );
INVxp33_ASAP7_75t_SL g724 ( .A(n_0), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_1), .A2(n_179), .B1(n_1141), .B2(n_1145), .Y(n_1171) );
INVx1_ASAP7_75t_L g977 ( .A(n_2), .Y(n_977) );
INVx1_ASAP7_75t_L g1093 ( .A(n_3), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_3), .A2(n_128), .B1(n_650), .B2(n_1104), .C(n_1110), .Y(n_1109) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_4), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_5), .A2(n_51), .B1(n_1141), .B2(n_1145), .Y(n_1179) );
INVx1_ASAP7_75t_L g269 ( .A(n_6), .Y(n_269) );
OAI221xp5_ASAP7_75t_SL g363 ( .A1(n_6), .A2(n_77), .B1(n_364), .B2(n_365), .C(n_369), .Y(n_363) );
INVx1_ASAP7_75t_L g438 ( .A(n_7), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_7), .A2(n_99), .B1(n_267), .B2(n_488), .Y(n_487) );
AOI21xp33_ASAP7_75t_L g992 ( .A1(n_8), .A2(n_578), .B(n_584), .Y(n_992) );
INVx1_ASAP7_75t_L g1014 ( .A(n_8), .Y(n_1014) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_9), .A2(n_188), .B1(n_364), .B2(n_365), .C(n_386), .Y(n_427) );
OA222x2_ASAP7_75t_L g503 ( .A1(n_9), .A2(n_42), .B1(n_193), .B2(n_504), .C1(n_508), .C2(n_512), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g1351 ( .A1(n_10), .A2(n_212), .B1(n_296), .B2(n_1352), .C(n_1354), .Y(n_1351) );
INVx1_ASAP7_75t_L g1373 ( .A(n_10), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g824 ( .A1(n_11), .A2(n_171), .B1(n_414), .B2(n_825), .C(n_827), .Y(n_824) );
INVx1_ASAP7_75t_L g856 ( .A(n_11), .Y(n_856) );
AND2x2_ASAP7_75t_L g271 ( .A(n_12), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g283 ( .A(n_12), .B(n_198), .Y(n_283) );
INVx1_ASAP7_75t_L g307 ( .A(n_12), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_12), .B(n_306), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g869 ( .A(n_13), .Y(n_869) );
INVx1_ASAP7_75t_L g545 ( .A(n_14), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_14), .A2(n_222), .B1(n_563), .B2(n_566), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_15), .A2(n_105), .B1(n_609), .B2(n_611), .Y(n_608) );
INVxp67_ASAP7_75t_SL g660 ( .A(n_15), .Y(n_660) );
INVx2_ASAP7_75t_L g1144 ( .A(n_16), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1146 ( .A(n_16), .B(n_95), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_16), .B(n_1150), .Y(n_1152) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_17), .A2(n_202), .B1(n_609), .B2(n_611), .Y(n_1081) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_17), .Y(n_1113) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_18), .A2(n_30), .B1(n_1148), .B2(n_1151), .Y(n_1165) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_19), .Y(n_877) );
INVx1_ASAP7_75t_L g624 ( .A(n_20), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g902 ( .A1(n_21), .A2(n_226), .B1(n_903), .B2(n_905), .Y(n_902) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_21), .A2(n_226), .B1(n_937), .B2(n_940), .Y(n_936) );
INVx1_ASAP7_75t_L g985 ( .A(n_22), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1009 ( .A1(n_22), .A2(n_127), .B1(n_275), .B2(n_541), .Y(n_1009) );
INVx1_ASAP7_75t_L g1047 ( .A(n_23), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_24), .A2(n_107), .B1(n_1148), .B2(n_1151), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_25), .A2(n_66), .B1(n_576), .B2(n_580), .C(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g734 ( .A1(n_25), .A2(n_27), .B1(n_277), .B2(n_541), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_26), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g684 ( .A1(n_27), .A2(n_118), .B1(n_685), .B2(n_686), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g884 ( .A(n_28), .Y(n_884) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_29), .A2(n_158), .B1(n_187), .B2(n_415), .C1(n_448), .C2(n_584), .Y(n_636) );
INVx1_ASAP7_75t_L g671 ( .A(n_29), .Y(n_671) );
INVx1_ASAP7_75t_L g528 ( .A(n_31), .Y(n_528) );
INVx1_ASAP7_75t_L g698 ( .A(n_32), .Y(n_698) );
OA222x2_ASAP7_75t_L g714 ( .A1(n_32), .A2(n_150), .B1(n_230), .B2(n_504), .C1(n_512), .C2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_33), .A2(n_91), .B1(n_1141), .B2(n_1300), .Y(n_1299) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_34), .A2(n_181), .B1(n_578), .B2(n_688), .C(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g730 ( .A(n_34), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_35), .A2(n_82), .B1(n_1141), .B2(n_1159), .Y(n_1158) );
AOI211xp5_ASAP7_75t_L g816 ( .A1(n_36), .A2(n_576), .B(n_817), .C(n_819), .Y(n_816) );
INVx1_ASAP7_75t_L g850 ( .A(n_36), .Y(n_850) );
INVx1_ASAP7_75t_L g1358 ( .A(n_37), .Y(n_1358) );
OAI21xp33_ASAP7_75t_L g530 ( .A1(n_38), .A2(n_504), .B(n_531), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g586 ( .A1(n_38), .A2(n_46), .B1(n_587), .B2(n_588), .C(n_590), .Y(n_586) );
OAI211xp5_ASAP7_75t_SL g973 ( .A1(n_39), .A2(n_593), .B(n_974), .C(n_978), .Y(n_973) );
INVx1_ASAP7_75t_L g998 ( .A(n_39), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_40), .A2(n_102), .B1(n_1084), .B2(n_1085), .C(n_1086), .Y(n_1083) );
INVx1_ASAP7_75t_L g1106 ( .A(n_40), .Y(n_1106) );
INVx1_ASAP7_75t_L g332 ( .A(n_41), .Y(n_332) );
INVx1_ASAP7_75t_L g353 ( .A(n_41), .Y(n_353) );
INVx1_ASAP7_75t_L g425 ( .A(n_42), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_43), .A2(n_135), .B1(n_277), .B2(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g384 ( .A(n_43), .Y(n_384) );
OAI221xp5_ASAP7_75t_L g813 ( .A1(n_44), .A2(n_215), .B1(n_566), .B2(n_570), .C(n_607), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_44), .A2(n_109), .B1(n_498), .B2(n_547), .Y(n_839) );
INVx1_ASAP7_75t_L g548 ( .A(n_45), .Y(n_548) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_46), .Y(n_598) );
INVx1_ASAP7_75t_L g1039 ( .A(n_47), .Y(n_1039) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_48), .A2(n_87), .B1(n_456), .B2(n_1091), .C(n_1092), .Y(n_1090) );
INVx1_ASAP7_75t_L g1112 ( .A(n_48), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_49), .A2(n_113), .B1(n_1141), .B2(n_1159), .Y(n_1176) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_50), .A2(n_141), .B1(n_615), .B2(n_617), .C(n_619), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_50), .A2(n_192), .B1(n_665), .B2(n_667), .C(n_669), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g606 ( .A1(n_52), .A2(n_214), .B1(n_566), .B2(n_570), .C(n_607), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_52), .A2(n_490), .B(n_512), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_53), .A2(n_196), .B1(n_1148), .B2(n_1151), .Y(n_1301) );
INVx1_ASAP7_75t_L g1125 ( .A(n_54), .Y(n_1125) );
INVx2_ASAP7_75t_L g339 ( .A(n_55), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_56), .Y(n_878) );
INVxp67_ASAP7_75t_SL g1345 ( .A(n_57), .Y(n_1345) );
OAI211xp5_ASAP7_75t_L g1380 ( .A1(n_57), .A2(n_570), .B(n_593), .C(n_1381), .Y(n_1380) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_58), .A2(n_62), .B1(n_626), .B2(n_629), .Y(n_625) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_58), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g1043 ( .A1(n_59), .A2(n_390), .B(n_578), .Y(n_1043) );
INVxp67_ASAP7_75t_L g1062 ( .A(n_59), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g733 ( .A(n_60), .Y(n_733) );
INVx1_ASAP7_75t_L g968 ( .A(n_61), .Y(n_968) );
INVx1_ASAP7_75t_L g646 ( .A(n_62), .Y(n_646) );
INVx1_ASAP7_75t_L g1094 ( .A(n_63), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g311 ( .A1(n_64), .A2(n_160), .B1(n_296), .B2(n_302), .C(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g385 ( .A(n_64), .Y(n_385) );
INVx1_ASAP7_75t_L g605 ( .A(n_65), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_65), .A2(n_508), .B(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_66), .A2(n_181), .B1(n_302), .B2(n_721), .C(n_722), .Y(n_720) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_67), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g908 ( .A1(n_68), .A2(n_217), .B1(n_909), .B2(n_912), .Y(n_908) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_68), .A2(n_217), .B1(n_958), .B2(n_960), .Y(n_957) );
INVx1_ASAP7_75t_L g442 ( .A(n_69), .Y(n_442) );
AOI221x1_ASAP7_75t_SL g467 ( .A1(n_69), .A2(n_85), .B1(n_296), .B2(n_309), .C(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g1347 ( .A(n_70), .Y(n_1347) );
INVx1_ASAP7_75t_L g705 ( .A(n_71), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_71), .B(n_712), .Y(n_711) );
XOR2x2_ASAP7_75t_L g808 ( .A(n_72), .B(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g995 ( .A(n_73), .Y(n_995) );
AOI22xp33_ASAP7_75t_L g1140 ( .A1(n_74), .A2(n_97), .B1(n_1141), .B2(n_1145), .Y(n_1140) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_75), .A2(n_108), .B1(n_1148), .B2(n_1151), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_76), .A2(n_122), .B1(n_580), .B2(n_987), .C(n_988), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_76), .A2(n_169), .B1(n_275), .B2(n_317), .Y(n_1015) );
INVx1_ASAP7_75t_L g288 ( .A(n_77), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g1349 ( .A1(n_78), .A2(n_205), .B1(n_554), .B2(n_555), .Y(n_1349) );
AOI21xp33_ASAP7_75t_L g1376 ( .A1(n_78), .A2(n_456), .B(n_578), .Y(n_1376) );
INVx1_ASAP7_75t_L g420 ( .A(n_79), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_79), .A2(n_188), .B1(n_496), .B2(n_501), .Y(n_495) );
OAI22xp5_ASAP7_75t_L g1048 ( .A1(n_80), .A2(n_161), .B1(n_626), .B2(n_629), .Y(n_1048) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_80), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_81), .A2(n_109), .B1(n_626), .B2(n_629), .Y(n_823) );
OAI211xp5_ASAP7_75t_L g832 ( .A1(n_81), .A2(n_712), .B(n_833), .C(n_836), .Y(n_832) );
INVx1_ASAP7_75t_L g707 ( .A(n_83), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_83), .A2(n_163), .B1(n_498), .B2(n_547), .Y(n_737) );
OAI221xp5_ASAP7_75t_L g249 ( .A1(n_84), .A2(n_232), .B1(n_250), .B2(n_256), .C(n_261), .Y(n_249) );
INVx1_ASAP7_75t_L g323 ( .A(n_84), .Y(n_323) );
INVx1_ASAP7_75t_L g458 ( .A(n_85), .Y(n_458) );
INVx1_ASAP7_75t_L g822 ( .A(n_86), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g1103 ( .A1(n_87), .A2(n_167), .B1(n_650), .B2(n_1104), .C(n_1105), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_88), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_88), .B(n_1125), .Y(n_1142) );
INVx1_ASAP7_75t_L g829 ( .A(n_89), .Y(n_829) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_90), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_92), .A2(n_143), .B1(n_694), .B2(n_768), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_92), .A2(n_93), .B1(n_275), .B2(n_541), .Y(n_801) );
INVx1_ASAP7_75t_L g780 ( .A(n_93), .Y(n_780) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_94), .A2(n_162), .B1(n_298), .B2(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_94), .A2(n_152), .B1(n_576), .B2(n_577), .C(n_578), .Y(n_575) );
AND2x2_ASAP7_75t_L g1143 ( .A(n_95), .B(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1150 ( .A(n_95), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_96), .A2(n_741), .B1(n_742), .B2(n_807), .Y(n_740) );
INVx1_ASAP7_75t_L g807 ( .A(n_96), .Y(n_807) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_96), .A2(n_151), .B1(n_1148), .B2(n_1151), .Y(n_1175) );
INVx1_ASAP7_75t_L g828 ( .A(n_98), .Y(n_828) );
INVx1_ASAP7_75t_L g449 ( .A(n_99), .Y(n_449) );
INVx1_ASAP7_75t_L g280 ( .A(n_100), .Y(n_280) );
OAI21xp33_ASAP7_75t_L g356 ( .A1(n_100), .A2(n_357), .B(n_361), .Y(n_356) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_101), .A2(n_138), .B1(n_626), .B2(n_629), .Y(n_1089) );
INVxp67_ASAP7_75t_SL g1115 ( .A(n_101), .Y(n_1115) );
INVx1_ASAP7_75t_L g1111 ( .A(n_102), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_103), .B(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g376 ( .A(n_103), .Y(n_376) );
INVx1_ASAP7_75t_L g404 ( .A(n_103), .Y(n_404) );
INVx1_ASAP7_75t_L g1041 ( .A(n_104), .Y(n_1041) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_105), .Y(n_639) );
INVxp67_ASAP7_75t_SL g991 ( .A(n_106), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g1003 ( .A1(n_106), .A2(n_122), .B1(n_1004), .B2(n_1006), .Y(n_1003) );
XOR2xp5_ASAP7_75t_L g405 ( .A(n_107), .B(n_406), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_110), .A2(n_244), .B1(n_245), .B2(n_246), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_110), .Y(n_244) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_111), .A2(n_223), .B1(n_315), .B2(n_541), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_111), .A2(n_185), .B1(n_362), .B2(n_576), .C(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_112), .A2(n_210), .B1(n_1148), .B2(n_1151), .Y(n_1147) );
AOI22xp5_ASAP7_75t_L g1155 ( .A1(n_114), .A2(n_116), .B1(n_1141), .B2(n_1145), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_115), .Y(n_445) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_117), .A2(n_174), .B1(n_566), .B2(n_570), .C(n_607), .Y(n_1080) );
OAI21xp33_ASAP7_75t_L g1100 ( .A1(n_117), .A2(n_490), .B(n_512), .Y(n_1100) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_118), .Y(n_723) );
OAI22xp33_ASAP7_75t_L g421 ( .A1(n_119), .A2(n_126), .B1(n_422), .B2(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g521 ( .A(n_119), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g1178 ( .A1(n_120), .A2(n_124), .B1(n_1148), .B2(n_1151), .Y(n_1178) );
AOI22xp33_ASAP7_75t_L g314 ( .A1(n_121), .A2(n_165), .B1(n_315), .B2(n_316), .Y(n_314) );
INVx1_ASAP7_75t_L g398 ( .A(n_121), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_123), .A2(n_971), .B1(n_1019), .B2(n_1020), .Y(n_970) );
INVx1_ASAP7_75t_L g1020 ( .A(n_123), .Y(n_1020) );
XOR2x2_ASAP7_75t_L g1024 ( .A(n_124), .B(n_1025), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_125), .A2(n_133), .B1(n_609), .B2(n_611), .Y(n_814) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_125), .Y(n_837) );
INVx1_ASAP7_75t_L g517 ( .A(n_126), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_127), .A2(n_169), .B1(n_574), .B2(n_694), .Y(n_993) );
INVx1_ASAP7_75t_L g1087 ( .A(n_128), .Y(n_1087) );
INVx1_ASAP7_75t_L g979 ( .A(n_129), .Y(n_979) );
OAI221xp5_ASAP7_75t_L g1000 ( .A1(n_129), .A2(n_168), .B1(n_501), .B2(n_1001), .C(n_1002), .Y(n_1000) );
INVx1_ASAP7_75t_L g1355 ( .A(n_130), .Y(n_1355) );
AOI22xp33_ASAP7_75t_L g1377 ( .A1(n_130), .A2(n_191), .B1(n_574), .B2(n_1378), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_131), .A2(n_184), .B1(n_315), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_131), .A2(n_223), .B1(n_362), .B2(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_SL g295 ( .A1(n_132), .A2(n_153), .B1(n_296), .B2(n_302), .C(n_303), .Y(n_295) );
INVx1_ASAP7_75t_L g388 ( .A(n_132), .Y(n_388) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_133), .Y(n_834) );
BUFx3_ASAP7_75t_L g329 ( .A(n_134), .Y(n_329) );
INVx1_ASAP7_75t_L g400 ( .A(n_135), .Y(n_400) );
INVx1_ASAP7_75t_L g980 ( .A(n_136), .Y(n_980) );
INVx1_ASAP7_75t_L g1079 ( .A(n_137), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_138), .A2(n_174), .B1(n_501), .B2(n_1001), .Y(n_1101) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_139), .A2(n_142), .B1(n_1148), .B2(n_1151), .Y(n_1160) );
INVx1_ASAP7_75t_L g1028 ( .A(n_140), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_141), .B(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_143), .A2(n_208), .B1(n_316), .B2(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g818 ( .A(n_144), .Y(n_818) );
INVx1_ASAP7_75t_L g621 ( .A(n_145), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_146), .A2(n_200), .B1(n_1141), .B2(n_1145), .Y(n_1166) );
INVx1_ASAP7_75t_L g1360 ( .A(n_147), .Y(n_1360) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_148), .Y(n_255) );
INVx1_ASAP7_75t_L g532 ( .A(n_149), .Y(n_532) );
INVx1_ASAP7_75t_L g709 ( .A(n_150), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_152), .A2(n_185), .B1(n_554), .B2(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g397 ( .A(n_153), .Y(n_397) );
AOI21xp5_ASAP7_75t_L g1033 ( .A1(n_154), .A2(n_362), .B(n_580), .Y(n_1033) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_154), .Y(n_1059) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_155), .Y(n_293) );
INVx1_ASAP7_75t_L g1346 ( .A(n_156), .Y(n_1346) );
INVx1_ASAP7_75t_L g930 ( .A(n_157), .Y(n_930) );
OAI211xp5_ASAP7_75t_L g943 ( .A1(n_157), .A2(n_944), .B(n_946), .C(n_948), .Y(n_943) );
INVx1_ASAP7_75t_L g656 ( .A(n_158), .Y(n_656) );
INVx1_ASAP7_75t_L g758 ( .A(n_159), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g797 ( .A1(n_159), .A2(n_475), .B1(n_512), .B2(n_798), .C(n_802), .Y(n_797) );
INVx1_ASAP7_75t_L g401 ( .A(n_160), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_161), .A2(n_183), .B1(n_490), .B2(n_496), .C(n_501), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_162), .A2(n_184), .B1(n_574), .B2(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g697 ( .A(n_163), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g870 ( .A(n_164), .Y(n_870) );
INVx1_ASAP7_75t_L g394 ( .A(n_165), .Y(n_394) );
INVx1_ASAP7_75t_L g1046 ( .A(n_166), .Y(n_1046) );
INVx1_ASAP7_75t_L g1088 ( .A(n_167), .Y(n_1088) );
INVx1_ASAP7_75t_L g996 ( .A(n_168), .Y(n_996) );
CKINVDCx5p33_ASAP7_75t_R g749 ( .A(n_170), .Y(n_749) );
INVx1_ASAP7_75t_L g843 ( .A(n_171), .Y(n_843) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
INVx1_ASAP7_75t_L g1036 ( .A(n_173), .Y(n_1036) );
OAI211xp5_ASAP7_75t_L g918 ( .A1(n_175), .A2(n_919), .B(n_921), .C(n_924), .Y(n_918) );
INVx1_ASAP7_75t_L g956 ( .A(n_175), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_176), .Y(n_435) );
XNOR2x1_ASAP7_75t_L g1075 ( .A(n_177), .B(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g820 ( .A(n_178), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_180), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_182), .Y(n_875) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_183), .A2(n_206), .B1(n_566), .B2(n_570), .C(n_607), .Y(n_1029) );
OAI21xp5_ASAP7_75t_L g1363 ( .A1(n_186), .A2(n_1018), .B(n_1364), .Y(n_1363) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_186), .A2(n_204), .B1(n_609), .B2(n_611), .Y(n_1365) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_187), .A2(n_266), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g812 ( .A(n_189), .Y(n_812) );
INVx1_ASAP7_75t_L g1342 ( .A(n_190), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1350 ( .A1(n_191), .A2(n_219), .B1(n_309), .B2(n_488), .Y(n_1350) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_192), .A2(n_632), .B(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g416 ( .A(n_193), .Y(n_416) );
INVx1_ASAP7_75t_L g744 ( .A(n_194), .Y(n_744) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_195), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_195), .A2(n_570), .B1(n_609), .B2(n_770), .C(n_777), .Y(n_769) );
INVx1_ASAP7_75t_L g1382 ( .A(n_196), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_196), .A2(n_1389), .B1(n_1392), .B2(n_1396), .Y(n_1388) );
XOR2xp5_ASAP7_75t_L g1393 ( .A(n_197), .B(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g272 ( .A(n_198), .Y(n_272) );
BUFx3_ASAP7_75t_L g306 ( .A(n_198), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g872 ( .A(n_199), .Y(n_872) );
INVx1_ASAP7_75t_L g738 ( .A(n_201), .Y(n_738) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_202), .Y(n_1097) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_203), .A2(n_578), .B(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g793 ( .A(n_203), .Y(n_793) );
INVxp33_ASAP7_75t_L g1362 ( .A(n_204), .Y(n_1362) );
INVx1_ASAP7_75t_L g1369 ( .A(n_205), .Y(n_1369) );
INVxp67_ASAP7_75t_SL g1073 ( .A(n_206), .Y(n_1073) );
INVx1_ASAP7_75t_L g975 ( .A(n_207), .Y(n_975) );
INVx1_ASAP7_75t_L g776 ( .A(n_208), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g755 ( .A(n_209), .Y(n_755) );
INVx2_ASAP7_75t_L g320 ( .A(n_211), .Y(n_320) );
INVx1_ASAP7_75t_L g337 ( .A(n_211), .Y(n_337) );
INVx1_ASAP7_75t_L g372 ( .A(n_211), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g1370 ( .A1(n_212), .A2(n_219), .B1(n_325), .B2(n_580), .C(n_1371), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_213), .A2(n_221), .B1(n_415), .B2(n_695), .Y(n_1044) );
INVxp67_ASAP7_75t_SL g1069 ( .A(n_213), .Y(n_1069) );
INVx1_ASAP7_75t_L g645 ( .A(n_214), .Y(n_645) );
INVxp67_ASAP7_75t_SL g835 ( .A(n_215), .Y(n_835) );
XOR2x2_ASAP7_75t_L g601 ( .A(n_216), .B(n_602), .Y(n_601) );
CKINVDCx5p33_ASAP7_75t_R g760 ( .A(n_218), .Y(n_760) );
INVx1_ASAP7_75t_L g1032 ( .A(n_220), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_221), .Y(n_1057) );
INVx1_ASAP7_75t_L g533 ( .A(n_222), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_224), .B(n_804), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_225), .Y(n_453) );
INVx1_ASAP7_75t_L g983 ( .A(n_227), .Y(n_983) );
INVxp67_ASAP7_75t_SL g524 ( .A(n_228), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_229), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g702 ( .A1(n_230), .A2(n_233), .B1(n_450), .B2(n_703), .C(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g757 ( .A(n_231), .Y(n_757) );
INVx1_ASAP7_75t_L g341 ( .A(n_232), .Y(n_341) );
INVxp67_ASAP7_75t_SL g717 ( .A(n_233), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_1118), .B(n_1132), .Y(n_234) );
XNOR2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_674), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
XNOR2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_522), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
XNOR2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_405), .Y(n_242) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_321), .Y(n_246) );
AOI21xp5_ASAP7_75t_SL g247 ( .A1(n_248), .A2(n_294), .B(n_318), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_270), .B(n_273), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_250), .A2(n_482), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx6f_ASAP7_75t_L g846 ( .A(n_251), .Y(n_846) );
BUFx4f_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g470 ( .A(n_252), .Y(n_470) );
INVx2_ASAP7_75t_L g655 ( .A(n_252), .Y(n_655) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g260 ( .A(n_254), .Y(n_260) );
INVx2_ASAP7_75t_L g264 ( .A(n_254), .Y(n_264) );
AND2x2_ASAP7_75t_L g268 ( .A(n_254), .B(n_255), .Y(n_268) );
INVx1_ASAP7_75t_L g292 ( .A(n_254), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_254), .B(n_301), .Y(n_300) );
NAND2x1_ASAP7_75t_L g473 ( .A(n_254), .B(n_255), .Y(n_473) );
OR2x2_ASAP7_75t_L g259 ( .A(n_255), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g263 ( .A(n_255), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g279 ( .A(n_255), .Y(n_279) );
BUFx2_ASAP7_75t_L g287 ( .A(n_255), .Y(n_287) );
INVx2_ASAP7_75t_L g301 ( .A(n_255), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_255), .B(n_264), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_256), .A2(n_818), .B1(n_842), .B2(n_843), .Y(n_841) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_L g799 ( .A(n_257), .Y(n_799) );
INVx4_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g481 ( .A(n_259), .Y(n_481) );
BUFx3_ASAP7_75t_L g729 ( .A(n_259), .Y(n_729) );
INVx2_ASAP7_75t_L g792 ( .A(n_259), .Y(n_792) );
BUFx2_ASAP7_75t_L g1064 ( .A(n_259), .Y(n_1064) );
AND2x2_ASAP7_75t_L g278 ( .A(n_260), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_265), .B1(n_266), .B2(n_269), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g310 ( .A(n_263), .Y(n_310) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_263), .Y(n_317) );
BUFx3_ASAP7_75t_L g541 ( .A(n_263), .Y(n_541) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_265), .A2(n_362), .B(n_363), .C(n_370), .Y(n_361) );
A2O1A1Ixp33_ASAP7_75t_L g274 ( .A1(n_266), .A2(n_275), .B(n_280), .C(n_281), .Y(n_274) );
BUFx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
BUFx3_ASAP7_75t_L g302 ( .A(n_267), .Y(n_302) );
BUFx3_ASAP7_75t_L g539 ( .A(n_267), .Y(n_539) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_267), .Y(n_666) );
AND2x2_ASAP7_75t_L g922 ( .A(n_267), .B(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g1353 ( .A(n_267), .Y(n_1353) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g557 ( .A(n_268), .Y(n_557) );
BUFx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_271), .B(n_372), .Y(n_511) );
AND2x2_ASAP7_75t_L g516 ( .A(n_271), .B(n_278), .Y(n_516) );
AND2x2_ASAP7_75t_L g519 ( .A(n_271), .B(n_520), .Y(n_519) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_272), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_284), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_277), .Y(n_315) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx3_ASAP7_75t_L g489 ( .A(n_278), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_278), .B(n_283), .Y(n_507) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g285 ( .A(n_283), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_283), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_283), .B(n_320), .Y(n_494) );
AOI22xp33_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B1(n_289), .B2(n_293), .Y(n_284) );
BUFx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g500 ( .A(n_287), .Y(n_500) );
AND2x2_ASAP7_75t_L g925 ( .A(n_287), .B(n_917), .Y(n_925) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g501 ( .A(n_290), .B(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g547 ( .A(n_290), .B(n_502), .Y(n_547) );
AND2x4_ASAP7_75t_L g929 ( .A(n_291), .B(n_306), .Y(n_929) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_293), .A2(n_341), .B1(n_342), .B2(n_348), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_308), .B1(n_311), .B2(n_314), .Y(n_294) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g554 ( .A(n_297), .Y(n_554) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g721 ( .A(n_299), .Y(n_721) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_300), .Y(n_520) );
BUFx3_ASAP7_75t_L g668 ( .A(n_300), .Y(n_668) );
AND2x4_ASAP7_75t_L g906 ( .A(n_300), .B(n_907), .Y(n_906) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVxp67_ASAP7_75t_L g904 ( .A(n_305), .Y(n_904) );
INVx1_ASAP7_75t_L g923 ( .A(n_305), .Y(n_923) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g313 ( .A(n_306), .B(n_307), .Y(n_313) );
BUFx2_ASAP7_75t_L g917 ( .A(n_306), .Y(n_917) );
INVx1_ASAP7_75t_L g933 ( .A(n_307), .Y(n_933) );
AND2x4_ASAP7_75t_L g509 ( .A(n_309), .B(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx4_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g476 ( .A(n_313), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_SL g853 ( .A(n_313), .B(n_335), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_313), .B(n_477), .Y(n_1008) );
BUFx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g552 ( .A(n_317), .Y(n_552) );
INVx1_ASAP7_75t_L g462 ( .A(n_318), .Y(n_462) );
BUFx2_ASAP7_75t_L g710 ( .A(n_318), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_318), .B(n_612), .Y(n_806) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g402 ( .A(n_319), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_L g465 ( .A(n_319), .B(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g559 ( .A(n_320), .Y(n_559) );
NAND3xp33_ASAP7_75t_SL g321 ( .A(n_322), .B(n_340), .C(n_355), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_333), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx8_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
INVx3_ASAP7_75t_L g426 ( .A(n_326), .Y(n_426) );
INVx2_ASAP7_75t_L g706 ( .A(n_326), .Y(n_706) );
INVx8_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_327), .B(n_373), .Y(n_595) );
BUFx3_ASAP7_75t_L g623 ( .A(n_327), .Y(n_623) );
AND2x2_ASAP7_75t_L g627 ( .A(n_327), .B(n_628), .Y(n_627) );
BUFx3_ASAP7_75t_L g695 ( .A(n_327), .Y(n_695) );
AND2x4_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
AND2x4_ASAP7_75t_L g345 ( .A(n_328), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_329), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_329), .B(n_353), .Y(n_360) );
OR2x2_ASAP7_75t_L g383 ( .A(n_329), .B(n_331), .Y(n_383) );
AND2x4_ASAP7_75t_L g419 ( .A(n_329), .B(n_368), .Y(n_419) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g346 ( .A(n_332), .Y(n_346) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g347 ( .A(n_334), .Y(n_347) );
OR2x2_ASAP7_75t_L g349 ( .A(n_334), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g357 ( .A(n_334), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_338), .Y(n_334) );
OR2x2_ASAP7_75t_L g379 ( .A(n_335), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g478 ( .A(n_335), .Y(n_478) );
HB1xp67_ASAP7_75t_L g967 ( .A(n_335), .Y(n_967) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g502 ( .A(n_336), .Y(n_502) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g412 ( .A(n_338), .Y(n_412) );
INVx1_ASAP7_75t_L g628 ( .A(n_338), .Y(n_628) );
INVx3_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_339), .B(n_376), .Y(n_380) );
BUFx3_ASAP7_75t_L g460 ( .A(n_339), .Y(n_460) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_347), .Y(n_342) );
INVx2_ASAP7_75t_L g396 ( .A(n_343), .Y(n_396) );
INVx2_ASAP7_75t_L g1368 ( .A(n_343), .Y(n_1368) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OR2x6_ASAP7_75t_SL g609 ( .A(n_344), .B(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_345), .Y(n_390) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_345), .Y(n_457) );
BUFx8_ASAP7_75t_L g584 ( .A(n_345), .Y(n_584) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
INVx4_ASAP7_75t_L g440 ( .A(n_350), .Y(n_440) );
INVx3_ASAP7_75t_L g763 ( .A(n_350), .Y(n_763) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_350), .Y(n_885) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g369 ( .A(n_351), .Y(n_369) );
BUFx2_ASAP7_75t_L g571 ( .A(n_351), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
BUFx2_ASAP7_75t_L g955 ( .A(n_352), .Y(n_955) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g368 ( .A(n_353), .Y(n_368) );
INVx2_ASAP7_75t_L g364 ( .A(n_354), .Y(n_364) );
AND2x4_ASAP7_75t_L g415 ( .A(n_354), .B(n_367), .Y(n_415) );
BUFx2_ASAP7_75t_L g952 ( .A(n_354), .Y(n_952) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_377), .Y(n_355) );
INVx1_ASAP7_75t_L g1038 ( .A(n_358), .Y(n_1038) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_359), .Y(n_589) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g393 ( .A(n_360), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_362), .A2(n_688), .B1(n_749), .B2(n_755), .Y(n_754) );
INVx3_ASAP7_75t_L g568 ( .A(n_364), .Y(n_568) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g565 ( .A(n_366), .B(n_373), .Y(n_565) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_369), .A2(n_382), .B1(n_400), .B2(n_401), .Y(n_399) );
INVx2_ASAP7_75t_L g772 ( .A(n_369), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_369), .A2(n_422), .B1(n_443), .B2(n_828), .C(n_829), .Y(n_827) );
AND2x4_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
OR2x2_ASAP7_75t_L g506 ( .A(n_371), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g662 ( .A(n_371), .Y(n_662) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g882 ( .A(n_372), .Y(n_882) );
INVx1_ASAP7_75t_L g429 ( .A(n_373), .Y(n_429) );
AND2x6_ASAP7_75t_L g567 ( .A(n_373), .B(n_568), .Y(n_567) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_374), .B(n_404), .Y(n_403) );
NAND3x1_ASAP7_75t_L g881 ( .A(n_374), .B(n_404), .C(n_882), .Y(n_881) );
OR2x4_ASAP7_75t_L g939 ( .A(n_374), .B(n_383), .Y(n_939) );
INVx1_ASAP7_75t_L g942 ( .A(n_374), .Y(n_942) );
AND2x4_ASAP7_75t_L g947 ( .A(n_374), .B(n_419), .Y(n_947) );
OR2x6_ASAP7_75t_L g962 ( .A(n_374), .B(n_393), .Y(n_962) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g459 ( .A(n_376), .B(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g965 ( .A(n_376), .Y(n_965) );
OAI33xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .A3(n_387), .B1(n_395), .B2(n_399), .B3(n_402), .Y(n_377) );
BUFx4f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx8_ASAP7_75t_L g867 ( .A(n_379), .Y(n_867) );
BUFx2_ASAP7_75t_L g578 ( .A(n_380), .Y(n_578) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B1(n_385), .B2(n_386), .Y(n_381) );
INVx1_ASAP7_75t_L g775 ( .A(n_382), .Y(n_775) );
BUFx4f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
BUFx3_ASAP7_75t_L g441 ( .A(n_383), .Y(n_441) );
INVx2_ASAP7_75t_L g448 ( .A(n_383), .Y(n_448) );
OR2x4_ASAP7_75t_L g959 ( .A(n_383), .B(n_942), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_391), .B2(n_394), .Y(n_387) );
INVx8_ASAP7_75t_L g577 ( .A(n_389), .Y(n_577) );
OAI221xp5_ASAP7_75t_L g982 ( .A1(n_389), .A2(n_983), .B1(n_984), .B2(n_985), .C(n_986), .Y(n_982) );
INVx5_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_SL g423 ( .A(n_390), .Y(n_423) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
INVx2_ASAP7_75t_SL g692 ( .A(n_390), .Y(n_692) );
INVx3_ASAP7_75t_L g703 ( .A(n_390), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_391), .A2(n_396), .B1(n_397), .B2(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g451 ( .A(n_392), .Y(n_451) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g436 ( .A(n_393), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g876 ( .A1(n_396), .A2(n_436), .B1(n_877), .B2(n_878), .Y(n_876) );
INVx3_ASAP7_75t_L g443 ( .A(n_403), .Y(n_443) );
NAND4xp75_ASAP7_75t_L g406 ( .A(n_407), .B(n_463), .C(n_503), .D(n_513), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_430), .B(n_461), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B(n_424), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_410), .A2(n_532), .B1(n_586), .B2(n_592), .Y(n_585) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g701 ( .A(n_411), .Y(n_701) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g610 ( .A(n_412), .Y(n_610) );
AND2x4_ASAP7_75t_L g612 ( .A(n_412), .B(n_415), .Y(n_612) );
AOI221xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_416), .B1(n_417), .B2(n_420), .C(n_421), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx12f_ASAP7_75t_L g574 ( .A(n_415), .Y(n_574) );
INVx5_ASAP7_75t_L g620 ( .A(n_415), .Y(n_620) );
BUFx2_ASAP7_75t_L g686 ( .A(n_415), .Y(n_686) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g1371 ( .A(n_418), .Y(n_1371) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g576 ( .A(n_419), .Y(n_576) );
BUFx2_ASAP7_75t_L g591 ( .A(n_419), .Y(n_591) );
AND2x2_ASAP7_75t_L g630 ( .A(n_419), .B(n_628), .Y(n_630) );
BUFx2_ASAP7_75t_L g688 ( .A(n_419), .Y(n_688) );
BUFx2_ASAP7_75t_L g708 ( .A(n_419), .Y(n_708) );
BUFx2_ASAP7_75t_L g987 ( .A(n_419), .Y(n_987) );
INVx2_ASAP7_75t_L g689 ( .A(n_423), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B(n_427), .C(n_428), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_426), .A2(n_528), .B1(n_548), .B2(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
OR2x6_ASAP7_75t_L g570 ( .A(n_429), .B(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_437), .B1(n_444), .B2(n_452), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_432), .A2(n_445), .B1(n_469), .B2(n_471), .Y(n_468) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_435), .A2(n_453), .B1(n_480), .B2(n_482), .C(n_487), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g454 ( .A(n_440), .Y(n_454) );
INVx2_ASAP7_75t_L g618 ( .A(n_440), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_441), .A2(n_820), .B1(n_821), .B2(n_822), .Y(n_819) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_441), .A2(n_771), .B1(n_869), .B2(n_870), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g883 ( .A1(n_441), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_883) );
OAI221xp5_ASAP7_75t_L g1092 ( .A1(n_441), .A2(n_443), .B1(n_1042), .B2(n_1093), .C(n_1094), .Y(n_1092) );
INVx3_ASAP7_75t_L g580 ( .A(n_443), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_443), .B(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_443), .A2(n_771), .B1(n_773), .B2(n_774), .C(n_776), .Y(n_770) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_449), .B2(n_450), .Y(n_444) );
BUFx4f_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_455), .B2(n_458), .C(n_459), .Y(n_452) );
OAI21xp33_ASAP7_75t_L g1031 ( .A1(n_454), .A2(n_1032), .B(n_1033), .Y(n_1031) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g587 ( .A(n_457), .Y(n_587) );
INVx1_ASAP7_75t_L g616 ( .A(n_457), .Y(n_616) );
INVx2_ASAP7_75t_L g826 ( .A(n_457), .Y(n_826) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_457), .Y(n_874) );
AND2x4_ASAP7_75t_L g941 ( .A(n_457), .B(n_942), .Y(n_941) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_459), .A2(n_620), .B1(n_621), .B2(n_622), .C(n_624), .Y(n_619) );
OAI21xp33_ASAP7_75t_L g817 ( .A1(n_459), .A2(n_583), .B(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g1086 ( .A1(n_459), .A2(n_778), .B1(n_1042), .B2(n_1087), .C(n_1088), .Y(n_1086) );
INVx3_ASAP7_75t_L g951 ( .A(n_460), .Y(n_951) );
OAI31xp33_ASAP7_75t_L g1364 ( .A1(n_461), .A2(n_1365), .A3(n_1366), .B(n_1380), .Y(n_1364) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AOI211x1_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_467), .B(n_474), .C(n_495), .Y(n_463) );
AOI222xp33_ASAP7_75t_L g1102 ( .A1(n_464), .A2(n_476), .B1(n_661), .B2(n_1103), .C1(n_1109), .C2(n_1113), .Y(n_1102) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI31xp33_ASAP7_75t_L g537 ( .A1(n_465), .A2(n_538), .A3(n_540), .B(n_542), .Y(n_537) );
INVx2_ASAP7_75t_L g659 ( .A(n_465), .Y(n_659) );
INVx2_ASAP7_75t_L g736 ( .A(n_465), .Y(n_736) );
INVx4_ASAP7_75t_L g789 ( .A(n_465), .Y(n_789) );
INVx1_ASAP7_75t_L g888 ( .A(n_465), .Y(n_888) );
INVx2_ASAP7_75t_L g1055 ( .A(n_465), .Y(n_1055) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g670 ( .A(n_470), .Y(n_670) );
BUFx6f_ASAP7_75t_L g1058 ( .A(n_470), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1068 ( .A(n_470), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_471), .A2(n_480), .B1(n_1036), .B2(n_1062), .Y(n_1061) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OR2x2_ASAP7_75t_L g512 ( .A(n_472), .B(n_511), .Y(n_512) );
OR2x2_ASAP7_75t_L g535 ( .A(n_472), .B(n_511), .Y(n_535) );
INVx2_ASAP7_75t_SL g896 ( .A(n_472), .Y(n_896) );
BUFx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_473), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_479), .B(n_490), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g549 ( .A(n_476), .B(n_550), .C(n_553), .Y(n_549) );
AOI322xp5_ASAP7_75t_L g648 ( .A1(n_476), .A2(n_649), .A3(n_652), .B1(n_658), .B2(n_660), .C1(n_661), .C2(n_664), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_476), .A2(n_720), .B(n_725), .C(n_737), .Y(n_719) );
INVx2_ASAP7_75t_L g897 ( .A(n_476), .Y(n_897) );
AOI322xp5_ASAP7_75t_L g1348 ( .A1(n_476), .A2(n_534), .A3(n_1012), .B1(n_1349), .B2(n_1350), .C1(n_1351), .C2(n_1360), .Y(n_1348) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g889 ( .A1(n_482), .A2(n_869), .B1(n_884), .B2(n_890), .Y(n_889) );
INVx6_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx5_ASAP7_75t_L g657 ( .A(n_483), .Y(n_657) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g672 ( .A(n_484), .Y(n_672) );
INVx2_ASAP7_75t_SL g855 ( .A(n_484), .Y(n_855) );
INVx1_ASAP7_75t_L g900 ( .A(n_484), .Y(n_900) );
INVx4_ASAP7_75t_L g1359 ( .A(n_484), .Y(n_1359) );
INVx8_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g916 ( .A(n_485), .B(n_917), .Y(n_916) );
BUFx2_ASAP7_75t_L g1060 ( .A(n_485), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g796 ( .A(n_489), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_490), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_490), .A2(n_726), .B(n_735), .Y(n_725) );
OAI21xp5_ASAP7_75t_SL g785 ( .A1(n_490), .A2(n_786), .B(n_790), .Y(n_785) );
OAI21xp5_ASAP7_75t_L g1010 ( .A1(n_490), .A2(n_1011), .B(n_1013), .Y(n_1010) );
OR2x6_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx4_ASAP7_75t_L g732 ( .A(n_491), .Y(n_732) );
BUFx4f_ASAP7_75t_L g794 ( .A(n_491), .Y(n_794) );
BUFx4f_ASAP7_75t_L g800 ( .A(n_491), .Y(n_800) );
BUFx4f_ASAP7_75t_L g842 ( .A(n_491), .Y(n_842) );
BUFx6f_ASAP7_75t_L g1065 ( .A(n_491), .Y(n_1065) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2x2_ASAP7_75t_L g498 ( .A(n_493), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g544 ( .A(n_498), .Y(n_544) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_498), .Y(n_1001) );
INVx2_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g515 ( .A(n_502), .Y(n_515) );
INVxp67_ASAP7_75t_L g747 ( .A(n_502), .Y(n_747) );
INVx1_ASAP7_75t_L g934 ( .A(n_502), .Y(n_934) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_506), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g663 ( .A(n_507), .Y(n_663) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_509), .A2(n_532), .B1(n_533), .B2(n_534), .Y(n_531) );
INVxp67_ASAP7_75t_L g715 ( .A(n_509), .Y(n_715) );
INVx1_ASAP7_75t_L g748 ( .A(n_509), .Y(n_748) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_509), .A2(n_534), .B1(n_661), .B2(n_812), .C1(n_834), .C2(n_835), .Y(n_833) );
AOI222xp33_ASAP7_75t_L g997 ( .A1(n_509), .A2(n_534), .B1(n_661), .B2(n_977), .C1(n_980), .C2(n_998), .Y(n_997) );
AOI222xp33_ASAP7_75t_L g1072 ( .A1(n_509), .A2(n_534), .B1(n_661), .B2(n_1028), .C1(n_1047), .C2(n_1073), .Y(n_1072) );
AOI211xp5_ASAP7_75t_L g1099 ( .A1(n_509), .A2(n_1079), .B(n_1100), .C(n_1101), .Y(n_1099) );
AOI222xp33_ASAP7_75t_L g1344 ( .A1(n_509), .A2(n_544), .B1(n_546), .B2(n_1345), .C1(n_1346), .C2(n_1347), .Y(n_1344) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_517), .B1(n_518), .B2(n_521), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_514), .B(n_528), .Y(n_527) );
AOI211xp5_ASAP7_75t_L g641 ( .A1(n_514), .A2(n_642), .B(n_643), .C(n_647), .Y(n_641) );
INVx3_ASAP7_75t_L g712 ( .A(n_514), .Y(n_712) );
AOI222xp33_ASAP7_75t_L g743 ( .A1(n_514), .A2(n_518), .B1(n_744), .B2(n_745), .C1(n_749), .C2(n_750), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_514), .A2(n_975), .B1(n_995), .B2(n_1017), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_514), .B(n_1115), .Y(n_1114) );
AOI211x1_ASAP7_75t_L g1341 ( .A1(n_514), .A2(n_1342), .B(n_1343), .C(n_1363), .Y(n_1341) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AND2x4_ASAP7_75t_L g518 ( .A(n_515), .B(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g597 ( .A(n_518), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_518), .B(n_639), .Y(n_638) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_518), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_518), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1018 ( .A(n_518), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_518), .B(n_1046), .Y(n_1074) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_520), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_600), .B1(n_601), .B2(n_673), .Y(n_522) );
INVx1_ASAP7_75t_L g673 ( .A(n_523), .Y(n_673) );
OAI21x1_ASAP7_75t_SL g523 ( .A1(n_524), .A2(n_525), .B(n_599), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g599 ( .A(n_524), .B(n_527), .C(n_529), .D(n_558), .Y(n_599) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND3xp33_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .C(n_558), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_536), .Y(n_529) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND3xp33_ASAP7_75t_SL g536 ( .A(n_537), .B(n_543), .C(n_549), .Y(n_536) );
OR3x1_ASAP7_75t_L g838 ( .A(n_542), .B(n_839), .C(n_840), .Y(n_838) );
AOI21xp33_ASAP7_75t_L g1361 ( .A1(n_542), .A2(n_661), .B(n_1362), .Y(n_1361) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_545), .B1(n_546), .B2(n_548), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_544), .A2(n_546), .B1(n_645), .B2(n_646), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_544), .A2(n_546), .B1(n_755), .B2(n_757), .Y(n_802) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g1006 ( .A(n_556), .Y(n_1006) );
INVx2_ASAP7_75t_L g1104 ( .A(n_556), .Y(n_1104) );
BUFx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_560), .B1(n_596), .B2(n_598), .Y(n_558) );
INVx2_ASAP7_75t_SL g637 ( .A(n_559), .Y(n_637) );
INVx1_ASAP7_75t_L g783 ( .A(n_559), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_572), .C(n_585), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_562), .B(n_569), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g607 ( .A(n_565), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_565), .A2(n_567), .B1(n_569), .B2(n_697), .C(n_698), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_565), .A2(n_567), .B1(n_757), .B2(n_758), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_565), .A2(n_567), .B1(n_569), .B2(n_979), .C(n_980), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_565), .A2(n_567), .B1(n_1346), .B2(n_1360), .Y(n_1381) );
INVx4_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g634 ( .A(n_571), .Y(n_634) );
INVx1_ASAP7_75t_L g945 ( .A(n_571), .Y(n_945) );
INVx1_ASAP7_75t_L g1375 ( .A(n_571), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B1(n_579), .B2(n_581), .Y(n_572) );
BUFx2_ASAP7_75t_L g1085 ( .A(n_574), .Y(n_1085) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g766 ( .A(n_584), .Y(n_766) );
INVx2_ASAP7_75t_SL g778 ( .A(n_584), .Y(n_778) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_584), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_588), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_588), .A2(n_872), .B1(n_873), .B2(n_875), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g1367 ( .A1(n_588), .A2(n_1358), .B1(n_1368), .B2(n_1369), .C(n_1370), .Y(n_1367) );
CKINVDCx8_ASAP7_75t_R g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g821 ( .A(n_589), .Y(n_821) );
INVx3_ASAP7_75t_L g984 ( .A(n_589), .Y(n_984) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI211xp5_ASAP7_75t_SL g604 ( .A1(n_594), .A2(n_605), .B(n_606), .C(n_608), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_594), .A2(n_700), .B1(n_702), .B2(n_709), .Y(n_699) );
AOI211xp5_ASAP7_75t_L g811 ( .A1(n_594), .A2(n_812), .B(n_813), .C(n_814), .Y(n_811) );
AOI211xp5_ASAP7_75t_L g1027 ( .A1(n_594), .A2(n_1028), .B(n_1029), .C(n_1030), .Y(n_1027) );
AOI211xp5_ASAP7_75t_L g1078 ( .A1(n_594), .A2(n_1079), .B(n_1080), .C(n_1081), .Y(n_1078) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g746 ( .A(n_595), .B(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_603), .B(n_640), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_613), .B(n_637), .C(n_638), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g976 ( .A(n_609), .Y(n_976) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_612), .A2(n_975), .B1(n_976), .B2(n_977), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g1045 ( .A1(n_612), .A2(n_976), .B1(n_1046), .B2(n_1047), .C(n_1048), .Y(n_1045) );
NOR3xp33_ASAP7_75t_SL g613 ( .A(n_614), .B(n_625), .C(n_631), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g768 ( .A(n_620), .Y(n_768) );
INVx2_ASAP7_75t_R g1091 ( .A(n_620), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_621), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g685 ( .A(n_622), .Y(n_685) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
BUFx3_ASAP7_75t_L g1378 ( .A(n_623), .Y(n_1378) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_624), .A2(n_654), .B1(n_656), .B2(n_657), .Y(n_653) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_627), .A2(n_630), .B1(n_995), .B2(n_996), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_627), .A2(n_630), .B1(n_1342), .B2(n_1347), .Y(n_1379) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_648), .Y(n_640) );
BUFx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g1110 ( .A1(n_654), .A2(n_1060), .B1(n_1111), .B2(n_1112), .Y(n_1110) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x6_ASAP7_75t_L g903 ( .A(n_655), .B(n_904), .Y(n_903) );
OR2x6_ASAP7_75t_L g911 ( .A(n_655), .B(n_907), .Y(n_911) );
INVxp67_ASAP7_75t_L g1108 ( .A(n_655), .Y(n_1108) );
INVx1_ASAP7_75t_L g1357 ( .A(n_655), .Y(n_1357) );
OAI33xp33_ASAP7_75t_L g840 ( .A1(n_659), .A2(n_841), .A3(n_844), .B1(n_847), .B2(n_852), .B3(n_854), .Y(n_840) );
AND2x4_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g1005 ( .A(n_668), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_670), .A2(n_822), .B1(n_855), .B2(n_856), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g844 ( .A1(n_672), .A2(n_820), .B1(n_829), .B2(n_845), .Y(n_844) );
XNOR2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_858), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_808), .B2(n_857), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
XNOR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_740), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_738), .B(n_739), .Y(n_679) );
AND3x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_713), .C(n_719), .Y(n_680) );
AOI31xp33_ASAP7_75t_L g739 ( .A1(n_681), .A2(n_713), .A3(n_719), .B(n_738), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_710), .B(n_711), .Y(n_681) );
NAND3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_696), .C(n_699), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B1(n_690), .B2(n_693), .Y(n_683) );
BUFx2_ASAP7_75t_SL g1084 ( .A(n_685), .Y(n_1084) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g989 ( .A(n_695), .Y(n_989) );
INVxp67_ASAP7_75t_L g753 ( .A(n_700), .Y(n_753) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_704) );
INVx2_ASAP7_75t_L g831 ( .A(n_710), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g972 ( .A1(n_710), .A2(n_973), .B(n_981), .Y(n_972) );
INVx1_ASAP7_75t_L g1095 ( .A(n_710), .Y(n_1095) );
INVx1_ASAP7_75t_L g1051 ( .A(n_712), .Y(n_1051) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B1(n_731), .B2(n_733), .C(n_734), .Y(n_726) );
INVx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g1013 ( .A1(n_731), .A2(n_799), .B1(n_983), .B2(n_1014), .C(n_1015), .Y(n_1013) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g851 ( .A(n_732), .Y(n_851) );
INVx1_ASAP7_75t_L g1012 ( .A(n_735), .Y(n_1012) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_751), .C(n_784), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_748), .Y(n_745) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_769), .B(n_781), .Y(n_751) );
OAI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_756), .C(n_759), .Y(n_752) );
OAI211xp5_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_761), .B(n_764), .C(n_767), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g798 ( .A1(n_760), .A2(n_773), .B1(n_799), .B2(n_800), .C(n_801), .Y(n_798) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
OAI211xp5_ASAP7_75t_L g990 ( .A1(n_762), .A2(n_991), .B(n_992), .C(n_993), .Y(n_990) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx3_ASAP7_75t_L g1042 ( .A(n_763), .Y(n_1042) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g790 ( .A1(n_779), .A2(n_791), .B1(n_793), .B2(n_794), .C(n_795), .Y(n_790) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
A2O1A1Ixp33_ASAP7_75t_SL g1026 ( .A1(n_782), .A2(n_1027), .B(n_1045), .C(n_1049), .Y(n_1026) );
BUFx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_797), .C(n_803), .Y(n_784) );
INVxp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_791), .A2(n_794), .B1(n_872), .B2(n_877), .Y(n_891) );
INVx1_ASAP7_75t_L g894 ( .A(n_791), .Y(n_894) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
BUFx2_ASAP7_75t_L g849 ( .A(n_792), .Y(n_849) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g857 ( .A(n_808), .Y(n_857) );
AOI211x1_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_830), .B(n_832), .C(n_838), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_815), .Y(n_810) );
NOR3xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_823), .C(n_824), .Y(n_815) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g847 ( .A1(n_828), .A2(n_848), .B1(n_850), .B2(n_851), .Y(n_847) );
INVx1_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g920 ( .A(n_842), .Y(n_920) );
INVx3_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g890 ( .A(n_846), .Y(n_890) );
INVx4_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx2_ASAP7_75t_L g1070 ( .A(n_853), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_859), .A2(n_860), .B1(n_1021), .B2(n_1022), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_969), .B2(n_970), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
XOR2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_968), .Y(n_863) );
AND3x1_ASAP7_75t_L g864 ( .A(n_865), .B(n_901), .C(n_935), .Y(n_864) );
NOR2xp33_ASAP7_75t_SL g865 ( .A(n_866), .B(n_887), .Y(n_865) );
OAI33xp33_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .A3(n_871), .B1(n_876), .B2(n_879), .B3(n_883), .Y(n_866) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_870), .A2(n_886), .B1(n_893), .B2(n_895), .Y(n_892) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g898 ( .A1(n_875), .A2(n_878), .B1(n_890), .B2(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx3_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
OAI33xp33_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_889), .A3(n_891), .B1(n_892), .B2(n_897), .B3(n_898), .Y(n_887) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx5_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
OAI31xp33_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_908), .A3(n_918), .B(n_931), .Y(n_901) );
INVx3_ASAP7_75t_L g1131 ( .A(n_903), .Y(n_1131) );
INVx4_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx3_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B1(n_927), .B2(n_930), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_926), .A2(n_949), .B1(n_953), .B2(n_956), .Y(n_948) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
BUFx3_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
AND2x4_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g1130 ( .A(n_933), .Y(n_1130) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_933), .B(n_1122), .Y(n_1387) );
OAI31xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_943), .A3(n_957), .B(n_963), .Y(n_935) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx2_ASAP7_75t_SL g938 ( .A(n_939), .Y(n_938) );
INVx2_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVxp67_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
CKINVDCx8_ASAP7_75t_R g946 ( .A(n_947), .Y(n_946) );
BUFx3_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
AND2x2_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
AND2x4_ASAP7_75t_L g954 ( .A(n_951), .B(n_955), .Y(n_954) );
BUFx6f_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
BUFx2_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx2_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
AND2x2_ASAP7_75t_SL g963 ( .A(n_964), .B(n_966), .Y(n_963) );
INVx1_ASAP7_75t_SL g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g966 ( .A(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
INVx1_ASAP7_75t_L g1019 ( .A(n_971), .Y(n_1019) );
NAND4xp25_ASAP7_75t_L g971 ( .A(n_972), .B(n_997), .C(n_999), .D(n_1016), .Y(n_971) );
NAND3xp33_ASAP7_75t_L g981 ( .A(n_982), .B(n_990), .C(n_994), .Y(n_981) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1010), .Y(n_999) );
NAND3xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1007), .C(n_1009), .Y(n_1002) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1017), .B(n_1097), .Y(n_1096) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
OA22x2_ASAP7_75t_L g1022 ( .A1(n_1023), .A2(n_1075), .B1(n_1116), .B2(n_1117), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
BUFx2_ASAP7_75t_SL g1117 ( .A(n_1024), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1052), .Y(n_1025) );
OAI21xp33_ASAP7_75t_L g1030 ( .A1(n_1031), .A2(n_1034), .B(n_1040), .Y(n_1030) );
OAI22xp5_ASAP7_75t_L g1063 ( .A1(n_1032), .A2(n_1041), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1036), .B1(n_1037), .B2(n_1039), .Y(n_1034) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1066 ( .A1(n_1039), .A2(n_1060), .B1(n_1067), .B2(n_1069), .Y(n_1066) );
OAI211xp5_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .B(n_1043), .C(n_1044), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1051), .Y(n_1049) );
NAND3xp33_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1072), .C(n_1074), .Y(n_1052) );
NOR2xp33_ASAP7_75t_SL g1053 ( .A(n_1054), .B(n_1071), .Y(n_1053) );
OAI33xp33_ASAP7_75t_L g1054 ( .A1(n_1055), .A2(n_1056), .A3(n_1061), .B1(n_1063), .B2(n_1066), .B3(n_1070), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1056 ( .A1(n_1057), .A2(n_1058), .B1(n_1059), .B2(n_1060), .Y(n_1056) );
OAI22xp33_ASAP7_75t_L g1105 ( .A1(n_1060), .A2(n_1094), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
INVx2_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1075), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1098), .Y(n_1076) );
A2O1A1Ixp33_ASAP7_75t_SL g1077 ( .A1(n_1078), .A2(n_1082), .B(n_1095), .C(n_1096), .Y(n_1077) );
NOR3xp33_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1089), .C(n_1090), .Y(n_1082) );
NAND3xp33_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1102), .C(n_1114), .Y(n_1098) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1108), .Y(n_1107) );
INVx2_ASAP7_75t_SL g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx3_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1128), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
NOR2xp33_ASAP7_75t_L g1123 ( .A(n_1124), .B(n_1126), .Y(n_1123) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_1124), .B(n_1127), .Y(n_1391) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1124), .Y(n_1399) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1127), .B(n_1399), .Y(n_1401) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1131), .Y(n_1129) );
AND2x4_ASAP7_75t_SL g1386 ( .A(n_1131), .B(n_1387), .Y(n_1386) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1337), .B1(n_1340), .B2(n_1383), .C(n_1388), .Y(n_1132) );
AND4x1_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1266), .C(n_1302), .D(n_1326), .Y(n_1133) );
NOR4xp25_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1207), .C(n_1229), .D(n_1243), .Y(n_1134) );
OAI211xp5_ASAP7_75t_L g1135 ( .A1(n_1136), .A2(n_1161), .B(n_1180), .C(n_1200), .Y(n_1135) );
OAI211xp5_ASAP7_75t_SL g1303 ( .A1(n_1136), .A2(n_1304), .B(n_1305), .C(n_1315), .Y(n_1303) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1153), .Y(n_1137) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1138), .B(n_1157), .Y(n_1248) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1138), .Y(n_1261) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1139), .B(n_1189), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1193 ( .A(n_1139), .B(n_1157), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1139), .B(n_1163), .Y(n_1236) );
INVx2_ASAP7_75t_SL g1242 ( .A(n_1139), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1147), .Y(n_1139) );
AND2x6_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1143), .Y(n_1141) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1142), .B(n_1146), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_1142), .B(n_1149), .Y(n_1148) );
AND2x6_ASAP7_75t_L g1151 ( .A(n_1142), .B(n_1152), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1142), .B(n_1146), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1142), .B(n_1146), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1144), .B(n_1150), .Y(n_1149) );
INVx2_ASAP7_75t_L g1339 ( .A(n_1151), .Y(n_1339) );
HB1xp67_ASAP7_75t_L g1398 ( .A(n_1152), .Y(n_1398) );
A2O1A1Ixp33_ASAP7_75t_L g1235 ( .A1(n_1153), .A2(n_1236), .B(n_1237), .C(n_1238), .Y(n_1235) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1153), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1157), .Y(n_1153) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1154), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1154), .B(n_1189), .Y(n_1211) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1154), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1154), .B(n_1236), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1154), .B(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1154), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1156), .Y(n_1154) );
CKINVDCx5p33_ASAP7_75t_R g1189 ( .A(n_1157), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1157), .B(n_1191), .Y(n_1234) );
HB1xp67_ASAP7_75t_SL g1277 ( .A(n_1157), .Y(n_1277) );
OAI322xp33_ASAP7_75t_L g1331 ( .A1(n_1157), .A2(n_1162), .A3(n_1173), .B1(n_1193), .B2(n_1304), .C1(n_1318), .C2(n_1332), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1167), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1162), .B(n_1215), .Y(n_1282) );
NOR2xp33_ASAP7_75t_L g1306 ( .A(n_1162), .B(n_1307), .Y(n_1306) );
CKINVDCx14_ASAP7_75t_R g1162 ( .A(n_1163), .Y(n_1162) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1163), .B(n_1193), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1163), .B(n_1215), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1163), .B(n_1185), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1163), .B(n_1242), .Y(n_1293) );
NOR2xp33_ASAP7_75t_L g1319 ( .A(n_1163), .B(n_1311), .Y(n_1319) );
NOR2xp33_ASAP7_75t_L g1323 ( .A(n_1163), .B(n_1241), .Y(n_1323) );
INVx3_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_1164), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1164), .B(n_1228), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1164), .B(n_1241), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_1164), .B(n_1258), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1164), .B(n_1169), .Y(n_1265) );
NOR2xp33_ASAP7_75t_L g1330 ( .A(n_1164), .B(n_1217), .Y(n_1330) );
AND2x4_ASAP7_75t_SL g1164 ( .A(n_1165), .B(n_1166), .Y(n_1164) );
INVx1_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1172), .Y(n_1168) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1169), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1169), .B(n_1195), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1198 ( .A(n_1169), .B(n_1174), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1169), .B(n_1173), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1258 ( .A(n_1169), .B(n_1174), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1169), .B(n_1276), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
OR2x2_ASAP7_75t_L g1213 ( .A(n_1172), .B(n_1185), .Y(n_1213) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1172), .Y(n_1245) );
OAI322xp33_ASAP7_75t_L g1271 ( .A1(n_1172), .A2(n_1222), .A3(n_1260), .B1(n_1272), .B2(n_1273), .C1(n_1274), .C2(n_1277), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1177), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1173), .B(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1174), .B(n_1177), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1174), .B(n_1218), .Y(n_1217) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1174), .B(n_1185), .Y(n_1224) );
NOR3xp33_ASAP7_75t_SL g1324 ( .A(n_1174), .B(n_1182), .C(n_1298), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1176), .Y(n_1174) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1177), .Y(n_1196) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1177), .Y(n_1218) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1177), .Y(n_1297) );
NAND2x1_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1179), .Y(n_1177) );
AOI221xp5_ASAP7_75t_L g1180 ( .A1(n_1181), .A2(n_1187), .B1(n_1190), .B2(n_1194), .C(n_1197), .Y(n_1180) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1181), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1184), .Y(n_1181) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1182), .B(n_1213), .Y(n_1212) );
A2O1A1Ixp33_ASAP7_75t_L g1295 ( .A1(n_1182), .A2(n_1211), .B(n_1219), .C(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1183), .B(n_1187), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1183), .B(n_1253), .Y(n_1252) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1183), .B(n_1195), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1290 ( .A(n_1183), .B(n_1248), .Y(n_1290) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1184), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1205 ( .A(n_1185), .B(n_1206), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1185), .B(n_1216), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1222 ( .A(n_1185), .B(n_1217), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1185), .B(n_1195), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g1283 ( .A(n_1185), .B(n_1284), .C(n_1286), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1185), .B(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1186), .Y(n_1206) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1187), .Y(n_1225) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
OR2x2_ASAP7_75t_L g1202 ( .A(n_1188), .B(n_1203), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1189), .B(n_1255), .Y(n_1254) );
HB1xp67_ASAP7_75t_SL g1273 ( .A(n_1189), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_1189), .B(n_1242), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1192), .Y(n_1190) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1191), .Y(n_1203) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1191), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1191), .B(n_1270), .Y(n_1269) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
OAI221xp5_ASAP7_75t_SL g1243 ( .A1(n_1193), .A2(n_1244), .B1(n_1248), .B2(n_1249), .C(n_1251), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1195), .B(n_1246), .Y(n_1250) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1195), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1199), .Y(n_1197) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1198), .Y(n_1294) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_1198), .A2(n_1210), .B1(n_1318), .B2(n_1320), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1204), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1202), .Y(n_1201) );
NOR2xp33_ASAP7_75t_L g1336 ( .A(n_1203), .B(n_1298), .Y(n_1336) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
AOI21xp33_ASAP7_75t_L g1238 ( .A1(n_1205), .A2(n_1239), .B(n_1240), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1214), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g1209 ( .A(n_1210), .B(n_1212), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1287 ( .A(n_1211), .B(n_1241), .Y(n_1287) );
INVxp67_ASAP7_75t_L g1335 ( .A(n_1212), .Y(n_1335) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1213), .Y(n_1219) );
O2A1O1Ixp33_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1219), .B(n_1220), .C(n_1221), .Y(n_1214) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1215), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1264 ( .A(n_1216), .B(n_1265), .Y(n_1264) );
NOR2xp33_ASAP7_75t_L g1285 ( .A(n_1216), .B(n_1245), .Y(n_1285) );
OAI21xp5_ASAP7_75t_SL g1312 ( .A1(n_1216), .A2(n_1293), .B(n_1296), .Y(n_1312) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
AOI211xp5_ASAP7_75t_L g1221 ( .A1(n_1222), .A2(n_1223), .B(n_1225), .C(n_1226), .Y(n_1221) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1222), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_1222), .B(n_1314), .Y(n_1313) );
CKINVDCx14_ASAP7_75t_R g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1228), .B(n_1261), .Y(n_1260) );
A2O1A1Ixp33_ASAP7_75t_L g1279 ( .A1(n_1228), .A2(n_1280), .B(n_1281), .C(n_1282), .Y(n_1279) );
A2O1A1Ixp33_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1232), .B(n_1233), .C(n_1235), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
NAND3xp33_ASAP7_75t_L g1263 ( .A(n_1234), .B(n_1261), .C(n_1264), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1237), .B(n_1261), .Y(n_1315) );
OAI221xp5_ASAP7_75t_L g1327 ( .A1(n_1239), .A2(n_1241), .B1(n_1297), .B2(n_1328), .C(n_1329), .Y(n_1327) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1240), .Y(n_1280) );
INVx2_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1246), .Y(n_1244) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1248), .Y(n_1270) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1248), .Y(n_1325) );
CKINVDCx14_ASAP7_75t_R g1249 ( .A(n_1250), .Y(n_1249) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_1252), .A2(n_1254), .B1(n_1256), .B2(n_1259), .C(n_1262), .Y(n_1251) );
OAI31xp33_ASAP7_75t_L g1309 ( .A1(n_1255), .A2(n_1310), .A3(n_1311), .B(n_1312), .Y(n_1309) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1258), .Y(n_1281) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1261), .B(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
OAI31xp33_ASAP7_75t_SL g1266 ( .A1(n_1267), .A2(n_1271), .A3(n_1278), .B(n_1298), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1269), .Y(n_1267) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1268), .Y(n_1308) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
NAND4xp25_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1283), .C(n_1288), .D(n_1295), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_1285), .Y(n_1284) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
OAI21xp5_ASAP7_75t_L g1288 ( .A1(n_1289), .A2(n_1291), .B(n_1294), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
INVxp67_ASAP7_75t_SL g1291 ( .A(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1293), .Y(n_1328) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1296), .Y(n_1304) );
NOR2xp33_ASAP7_75t_L g1321 ( .A(n_1297), .B(n_1322), .Y(n_1321) );
INVx3_ASAP7_75t_L g1316 ( .A(n_1298), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1301), .Y(n_1298) );
AOI222xp33_ASAP7_75t_L g1302 ( .A1(n_1303), .A2(n_1316), .B1(n_1317), .B2(n_1324), .C1(n_1325), .C2(n_1403), .Y(n_1302) );
AOI211xp5_ASAP7_75t_L g1305 ( .A1(n_1306), .A2(n_1308), .B(n_1309), .C(n_1313), .Y(n_1305) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVxp67_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
OAI31xp33_ASAP7_75t_L g1326 ( .A1(n_1327), .A2(n_1331), .A3(n_1333), .B(n_1336), .Y(n_1326) );
INVxp67_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVxp67_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
CKINVDCx20_ASAP7_75t_R g1337 ( .A(n_1338), .Y(n_1337) );
CKINVDCx20_ASAP7_75t_R g1338 ( .A(n_1339), .Y(n_1338) );
XOR2x2_ASAP7_75t_L g1340 ( .A(n_1341), .B(n_1382), .Y(n_1340) );
HB1xp67_ASAP7_75t_L g1395 ( .A(n_1341), .Y(n_1395) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1348), .C(n_1361), .Y(n_1343) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
OAI22xp5_ASAP7_75t_L g1354 ( .A1(n_1355), .A2(n_1356), .B1(n_1358), .B2(n_1359), .Y(n_1354) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
NAND3xp33_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1372), .C(n_1379), .Y(n_1366) );
OAI211xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B(n_1376), .C(n_1377), .Y(n_1372) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
CKINVDCx20_ASAP7_75t_R g1383 ( .A(n_1384), .Y(n_1383) );
CKINVDCx20_ASAP7_75t_R g1384 ( .A(n_1385), .Y(n_1384) );
INVx3_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
BUFx3_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVxp33_ASAP7_75t_SL g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
HB1xp67_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
OAI21xp5_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1399), .B(n_1400), .Y(n_1397) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1401), .Y(n_1400) );
endmodule