module real_aes_15983_n_361 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_361);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_361;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1760;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_1499;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_1612;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_1171;
wire n_569;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_1403;
wire n_643;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_1772;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1761;
wire n_1015;
wire n_1375;
wire n_863;
wire n_525;
wire n_1790;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_0), .A2(n_63), .B1(n_544), .B2(n_690), .Y(n_689) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_0), .Y(n_720) );
XNOR2xp5_ASAP7_75t_L g1379 ( .A(n_1), .B(n_1380), .Y(n_1379) );
OAI22xp33_ASAP7_75t_L g1766 ( .A1(n_2), .A2(n_329), .B1(n_550), .B2(n_552), .Y(n_1766) );
OAI22xp33_ASAP7_75t_SL g1776 ( .A1(n_2), .A2(n_329), .B1(n_510), .B2(n_1204), .Y(n_1776) );
INVx1_ASAP7_75t_L g929 ( .A(n_3), .Y(n_929) );
INVx1_ASAP7_75t_L g375 ( .A(n_4), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_4), .B(n_385), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_5), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_6), .A2(n_265), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_6), .A2(n_205), .B1(n_902), .B2(n_905), .Y(n_901) );
INVx1_ASAP7_75t_L g1436 ( .A(n_7), .Y(n_1436) );
OAI22xp33_ASAP7_75t_L g1329 ( .A1(n_8), .A2(n_62), .B1(n_377), .B2(n_552), .Y(n_1329) );
OAI22xp33_ASAP7_75t_L g1370 ( .A1(n_8), .A2(n_62), .B1(n_591), .B2(n_1134), .Y(n_1370) );
OAI22xp5_ASAP7_75t_SL g1454 ( .A1(n_9), .A2(n_232), .B1(n_527), .B2(n_573), .Y(n_1454) );
OAI22xp5_ASAP7_75t_L g1457 ( .A1(n_9), .A2(n_232), .B1(n_1417), .B2(n_1458), .Y(n_1457) );
INVx1_ASAP7_75t_L g1266 ( .A(n_10), .Y(n_1266) );
OAI22xp33_ASAP7_75t_SL g780 ( .A1(n_11), .A2(n_346), .B1(n_550), .B2(n_699), .Y(n_780) );
OAI22xp33_ASAP7_75t_L g794 ( .A1(n_11), .A2(n_189), .B1(n_510), .B2(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g1221 ( .A(n_12), .Y(n_1221) );
INVx1_ASAP7_75t_L g1427 ( .A(n_13), .Y(n_1427) );
INVx1_ASAP7_75t_L g870 ( .A(n_14), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_14), .A2(n_265), .B1(n_905), .B2(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1267 ( .A1(n_15), .A2(n_163), .B1(n_377), .B2(n_552), .Y(n_1267) );
OAI22xp5_ASAP7_75t_L g1269 ( .A1(n_15), .A2(n_163), .B1(n_795), .B2(n_1270), .Y(n_1269) );
AOI22xp5_ASAP7_75t_L g1529 ( .A1(n_16), .A2(n_217), .B1(n_1516), .B2(n_1530), .Y(n_1529) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_17), .Y(n_621) );
INVx1_ASAP7_75t_L g662 ( .A(n_18), .Y(n_662) );
OAI22xp33_ASAP7_75t_L g1455 ( .A1(n_19), .A2(n_161), .B1(n_377), .B2(n_552), .Y(n_1455) );
OAI22xp33_ASAP7_75t_L g1464 ( .A1(n_19), .A2(n_161), .B1(n_589), .B2(n_591), .Y(n_1464) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_20), .A2(n_47), .B1(n_591), .B2(n_1134), .Y(n_1133) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_20), .A2(n_47), .B1(n_377), .B2(n_552), .Y(n_1155) );
AOI22xp33_ASAP7_75t_L g1550 ( .A1(n_21), .A2(n_99), .B1(n_1516), .B2(n_1520), .Y(n_1550) );
INVx1_ASAP7_75t_L g971 ( .A(n_22), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g981 ( .A1(n_22), .A2(n_301), .B1(n_678), .B2(n_982), .C(n_983), .Y(n_981) );
CKINVDCx5p33_ASAP7_75t_R g803 ( .A(n_23), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_24), .A2(n_341), .B1(n_1523), .B2(n_1526), .Y(n_1613) );
OAI22xp33_ASAP7_75t_L g1773 ( .A1(n_25), .A2(n_303), .B1(n_837), .B2(n_1774), .Y(n_1773) );
OAI22xp33_ASAP7_75t_L g1780 ( .A1(n_25), .A2(n_303), .B1(n_505), .B2(n_513), .Y(n_1780) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_26), .A2(n_324), .B1(n_573), .B2(n_574), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_26), .A2(n_324), .B1(n_579), .B2(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g404 ( .A(n_27), .Y(n_404) );
XNOR2xp5_ASAP7_75t_L g650 ( .A(n_28), .B(n_651), .Y(n_650) );
OAI22xp33_ASAP7_75t_SL g1039 ( .A1(n_29), .A2(n_274), .B1(n_510), .B2(n_795), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g1046 ( .A1(n_29), .A2(n_274), .B1(n_550), .B2(n_838), .Y(n_1046) );
INVx1_ASAP7_75t_L g1497 ( .A(n_30), .Y(n_1497) );
INVx1_ASAP7_75t_L g1217 ( .A(n_31), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_32), .A2(n_289), .B1(n_994), .B2(n_996), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1002 ( .A1(n_32), .A2(n_166), .B1(n_1003), .B2(n_1004), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g1243 ( .A1(n_33), .A2(n_174), .B1(n_717), .B2(n_882), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_33), .A2(n_212), .B1(n_664), .B2(n_1004), .Y(n_1255) );
AOI22xp5_ASAP7_75t_L g1522 ( .A1(n_34), .A2(n_225), .B1(n_1523), .B2(n_1526), .Y(n_1522) );
INVx1_ASAP7_75t_L g437 ( .A(n_35), .Y(n_437) );
INVx1_ASAP7_75t_L g1054 ( .A(n_36), .Y(n_1054) );
OAI221xp5_ASAP7_75t_L g941 ( .A1(n_37), .A2(n_94), .B1(n_513), .B2(n_795), .C(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g955 ( .A(n_37), .Y(n_955) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_38), .A2(n_327), .B1(n_830), .B2(n_837), .Y(n_1200) );
OAI22xp33_ASAP7_75t_L g1210 ( .A1(n_38), .A2(n_327), .B1(n_505), .B2(n_513), .Y(n_1210) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_39), .Y(n_370) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_39), .B(n_368), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1611 ( .A1(n_40), .A2(n_200), .B1(n_1516), .B2(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1391 ( .A(n_41), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1564 ( .A1(n_42), .A2(n_213), .B1(n_1516), .B2(n_1520), .Y(n_1564) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_43), .Y(n_1105) );
INVx1_ASAP7_75t_L g1452 ( .A(n_44), .Y(n_1452) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_45), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_45), .A2(n_63), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g1486 ( .A(n_46), .Y(n_1486) );
INVx1_ASAP7_75t_L g1284 ( .A(n_48), .Y(n_1284) );
OAI22xp33_ASAP7_75t_L g1201 ( .A1(n_49), .A2(n_280), .B1(n_550), .B2(n_838), .Y(n_1201) );
OAI22xp33_ASAP7_75t_SL g1203 ( .A1(n_49), .A2(n_280), .B1(n_510), .B2(n_1204), .Y(n_1203) );
INVx1_ASAP7_75t_L g1351 ( .A(n_50), .Y(n_1351) );
INVx1_ASAP7_75t_L g503 ( .A(n_51), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g522 ( .A1(n_51), .A2(n_352), .B1(n_523), .B2(n_527), .Y(n_522) );
INVx1_ASAP7_75t_L g1160 ( .A(n_52), .Y(n_1160) );
XNOR2x1_ASAP7_75t_L g1016 ( .A(n_53), .B(n_1017), .Y(n_1016) );
AOI22xp5_ASAP7_75t_L g1537 ( .A1(n_54), .A2(n_177), .B1(n_1516), .B2(n_1520), .Y(n_1537) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_55), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g867 ( .A(n_56), .Y(n_867) );
INVx1_ASAP7_75t_L g1394 ( .A(n_57), .Y(n_1394) );
INVx1_ASAP7_75t_L g1754 ( .A(n_58), .Y(n_1754) );
AOI22xp33_ASAP7_75t_SL g1235 ( .A1(n_59), .A2(n_212), .B1(n_854), .B2(n_1236), .Y(n_1235) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_59), .A2(n_174), .B1(n_1247), .B2(n_1248), .Y(n_1246) );
INVx1_ASAP7_75t_L g932 ( .A(n_60), .Y(n_932) );
INVx1_ASAP7_75t_L g420 ( .A(n_61), .Y(n_420) );
INVx1_ASAP7_75t_L g1435 ( .A(n_64), .Y(n_1435) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_65), .B(n_488), .Y(n_944) );
INVxp67_ASAP7_75t_SL g952 ( .A(n_65), .Y(n_952) );
OAI211xp5_ASAP7_75t_SL g1136 ( .A1(n_66), .A2(n_645), .B(n_793), .C(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1151 ( .A(n_66), .Y(n_1151) );
OAI211xp5_ASAP7_75t_L g1470 ( .A1(n_67), .A2(n_582), .B(n_584), .C(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1479 ( .A(n_67), .Y(n_1479) );
OAI211xp5_ASAP7_75t_L g769 ( .A1(n_68), .A2(n_770), .B(n_771), .C(n_775), .Y(n_769) );
INVx1_ASAP7_75t_L g792 ( .A(n_68), .Y(n_792) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_69), .A2(n_183), .B1(n_579), .B2(n_580), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1152 ( .A1(n_69), .A2(n_183), .B1(n_573), .B2(n_1153), .Y(n_1152) );
INVx1_ASAP7_75t_L g1433 ( .A(n_70), .Y(n_1433) );
CKINVDCx5p33_ASAP7_75t_R g742 ( .A(n_71), .Y(n_742) );
INVx1_ASAP7_75t_L g692 ( .A(n_72), .Y(n_692) );
OAI222xp33_ASAP7_75t_L g855 ( .A1(n_73), .A2(n_191), .B1(n_551), .B2(n_779), .C1(n_856), .C2(n_858), .Y(n_855) );
OAI222xp33_ASAP7_75t_L g888 ( .A1(n_73), .A2(n_191), .B1(n_233), .B2(n_889), .C1(n_890), .C2(n_891), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_74), .A2(n_132), .B1(n_830), .B2(n_837), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_74), .A2(n_132), .B1(n_505), .B2(n_513), .Y(n_984) );
OAI211xp5_ASAP7_75t_L g1296 ( .A1(n_75), .A2(n_1147), .B(n_1149), .C(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1306 ( .A(n_75), .Y(n_1306) );
INVx1_ASAP7_75t_L g1220 ( .A(n_76), .Y(n_1220) );
OAI22xp33_ASAP7_75t_L g947 ( .A1(n_77), .A2(n_194), .B1(n_510), .B2(n_948), .Y(n_947) );
INVxp67_ASAP7_75t_SL g954 ( .A(n_77), .Y(n_954) );
INVx1_ASAP7_75t_L g1753 ( .A(n_78), .Y(n_1753) );
INVx1_ASAP7_75t_L g1261 ( .A(n_79), .Y(n_1261) );
INVx1_ASAP7_75t_L g1496 ( .A(n_80), .Y(n_1496) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_81), .Y(n_816) );
INVx1_ASAP7_75t_L g697 ( .A(n_82), .Y(n_697) );
INVx1_ASAP7_75t_L g1492 ( .A(n_83), .Y(n_1492) );
INVx1_ASAP7_75t_L g1173 ( .A(n_84), .Y(n_1173) );
CKINVDCx5p33_ASAP7_75t_R g1067 ( .A(n_85), .Y(n_1067) );
INVx1_ASAP7_75t_L g1031 ( .A(n_86), .Y(n_1031) );
OAI211xp5_ASAP7_75t_L g1195 ( .A1(n_87), .A2(n_771), .B(n_1196), .C(n_1197), .Y(n_1195) );
INVx1_ASAP7_75t_L g1207 ( .A(n_87), .Y(n_1207) );
INVx1_ASAP7_75t_L g683 ( .A(n_88), .Y(n_683) );
XNOR2xp5_ASAP7_75t_L g960 ( .A(n_89), .B(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g931 ( .A(n_90), .Y(n_931) );
INVx1_ASAP7_75t_L g1389 ( .A(n_91), .Y(n_1389) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_92), .A2(n_125), .B1(n_505), .B2(n_513), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1050 ( .A1(n_92), .A2(n_125), .B1(n_830), .B2(n_837), .Y(n_1050) );
XNOR2xp5_ASAP7_75t_L g1094 ( .A(n_93), .B(n_1095), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g957 ( .A1(n_94), .A2(n_194), .B1(n_550), .B2(n_838), .Y(n_957) );
INVx1_ASAP7_75t_L g1081 ( .A(n_95), .Y(n_1081) );
OAI211xp5_ASAP7_75t_L g1087 ( .A1(n_95), .A2(n_584), .B(n_1088), .C(n_1091), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_96), .A2(n_279), .B1(n_550), .B2(n_830), .Y(n_829) );
OAI22xp5_ASAP7_75t_SL g841 ( .A1(n_96), .A2(n_141), .B1(n_505), .B2(n_510), .Y(n_841) );
INVx1_ASAP7_75t_L g946 ( .A(n_97), .Y(n_946) );
INVx1_ASAP7_75t_L g1171 ( .A(n_98), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_100), .Y(n_833) );
INVx1_ASAP7_75t_L g1473 ( .A(n_101), .Y(n_1473) );
OAI211xp5_ASAP7_75t_L g1477 ( .A1(n_101), .A2(n_466), .B(n_535), .C(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1224 ( .A(n_102), .Y(n_1224) );
CKINVDCx5p33_ASAP7_75t_R g802 ( .A(n_103), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_104), .Y(n_740) );
AOI22xp33_ASAP7_75t_SL g1244 ( .A1(n_105), .A2(n_358), .B1(n_854), .B2(n_1236), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g1257 ( .A1(n_105), .A2(n_107), .B1(n_1250), .B2(n_1253), .Y(n_1257) );
OAI22xp33_ASAP7_75t_SL g1337 ( .A1(n_106), .A2(n_278), .B1(n_523), .B2(n_1338), .Y(n_1337) );
OAI22xp33_ASAP7_75t_L g1374 ( .A1(n_106), .A2(n_278), .B1(n_580), .B2(n_1310), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1239 ( .A1(n_107), .A2(n_330), .B1(n_882), .B2(n_1240), .Y(n_1239) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_108), .A2(n_256), .B1(n_994), .B2(n_998), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_108), .A2(n_178), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
XOR2xp5_ASAP7_75t_L g735 ( .A(n_109), .B(n_736), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g1541 ( .A1(n_109), .A2(n_224), .B1(n_1523), .B2(n_1526), .Y(n_1541) );
INVx1_ASAP7_75t_L g1747 ( .A(n_110), .Y(n_1747) );
INVx1_ASAP7_75t_L g1392 ( .A(n_111), .Y(n_1392) );
INVx1_ASAP7_75t_L g665 ( .A(n_112), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_112), .A2(n_294), .B1(n_709), .B2(n_717), .Y(n_716) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_113), .Y(n_1108) );
INVx1_ASAP7_75t_L g1491 ( .A(n_114), .Y(n_1491) );
CKINVDCx5p33_ASAP7_75t_R g812 ( .A(n_115), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g1409 ( .A1(n_116), .A2(n_152), .B1(n_550), .B2(n_552), .Y(n_1409) );
OAI22xp5_ASAP7_75t_L g1411 ( .A1(n_116), .A2(n_139), .B1(n_510), .B2(n_579), .Y(n_1411) );
INVx1_ASAP7_75t_L g1385 ( .A(n_117), .Y(n_1385) );
INVx1_ASAP7_75t_L g1199 ( .A(n_118), .Y(n_1199) );
INVx1_ASAP7_75t_L g1396 ( .A(n_119), .Y(n_1396) );
OAI211xp5_ASAP7_75t_L g1078 ( .A1(n_120), .A2(n_609), .B(n_771), .C(n_1079), .Y(n_1078) );
INVx1_ASAP7_75t_L g1092 ( .A(n_120), .Y(n_1092) );
INVx1_ASAP7_75t_L g368 ( .A(n_121), .Y(n_368) );
INVx1_ASAP7_75t_L g1358 ( .A(n_122), .Y(n_1358) );
INVx1_ASAP7_75t_L g1430 ( .A(n_123), .Y(n_1430) );
INVx1_ASAP7_75t_L g679 ( .A(n_124), .Y(n_679) );
XNOR2xp5_ASAP7_75t_L g1791 ( .A(n_126), .B(n_1792), .Y(n_1791) );
OAI22xp33_ASAP7_75t_L g1084 ( .A1(n_127), .A2(n_299), .B1(n_524), .B2(n_552), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1093 ( .A1(n_127), .A2(n_168), .B1(n_505), .B2(n_513), .Y(n_1093) );
XOR2xp5_ASAP7_75t_L g847 ( .A(n_128), .B(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g1024 ( .A(n_129), .Y(n_1024) );
INVx1_ASAP7_75t_L g1021 ( .A(n_130), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g1405 ( .A(n_131), .Y(n_1405) );
INVx1_ASAP7_75t_L g1335 ( .A(n_133), .Y(n_1335) );
AOI22xp5_ASAP7_75t_L g1546 ( .A1(n_134), .A2(n_325), .B1(n_1523), .B2(n_1526), .Y(n_1546) );
INVx1_ASAP7_75t_L g660 ( .A(n_135), .Y(n_660) );
INVx1_ASAP7_75t_L g1757 ( .A(n_136), .Y(n_1757) );
AOI22xp33_ASAP7_75t_L g1291 ( .A1(n_137), .A2(n_199), .B1(n_1292), .B2(n_1293), .Y(n_1291) );
INVx1_ASAP7_75t_L g1315 ( .A(n_137), .Y(n_1315) );
INVx1_ASAP7_75t_L g1472 ( .A(n_138), .Y(n_1472) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_139), .A2(n_226), .B1(n_523), .B2(n_1408), .Y(n_1407) );
OAI22xp33_ASAP7_75t_SL g836 ( .A1(n_140), .A2(n_141), .B1(n_837), .B2(n_838), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_140), .A2(n_146), .B1(n_789), .B2(n_790), .Y(n_845) );
INVx1_ASAP7_75t_L g1176 ( .A(n_142), .Y(n_1176) );
INVx1_ASAP7_75t_L g1769 ( .A(n_143), .Y(n_1769) );
AOI22xp5_ASAP7_75t_L g1515 ( .A1(n_144), .A2(n_227), .B1(n_1516), .B2(n_1520), .Y(n_1515) );
CKINVDCx5p33_ASAP7_75t_R g612 ( .A(n_145), .Y(n_612) );
INVx1_ASAP7_75t_L g834 ( .A(n_146), .Y(n_834) );
INVx1_ASAP7_75t_L g1489 ( .A(n_147), .Y(n_1489) );
INVx1_ASAP7_75t_L g964 ( .A(n_148), .Y(n_964) );
INVx1_ASAP7_75t_L g1043 ( .A(n_149), .Y(n_1043) );
OAI211xp5_ASAP7_75t_L g1047 ( .A1(n_149), .A2(n_771), .B(n_937), .C(n_1048), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1531 ( .A1(n_150), .A2(n_240), .B1(n_1523), .B2(n_1526), .Y(n_1531) );
CKINVDCx5p33_ASAP7_75t_R g1042 ( .A(n_151), .Y(n_1042) );
OAI22xp5_ASAP7_75t_L g1416 ( .A1(n_152), .A2(n_226), .B1(n_591), .B2(n_1417), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g620 ( .A(n_153), .Y(n_620) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_154), .Y(n_1106) );
OAI22xp33_ASAP7_75t_L g1121 ( .A1(n_155), .A2(n_196), .B1(n_552), .B2(n_837), .Y(n_1121) );
OAI22xp33_ASAP7_75t_L g1127 ( .A1(n_155), .A2(n_186), .B1(n_505), .B2(n_513), .Y(n_1127) );
OAI22xp33_ASAP7_75t_L g1474 ( .A1(n_156), .A2(n_171), .B1(n_589), .B2(n_1475), .Y(n_1474) );
OAI22xp33_ASAP7_75t_L g1481 ( .A1(n_156), .A2(n_171), .B1(n_550), .B2(n_552), .Y(n_1481) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_157), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g1099 ( .A(n_158), .Y(n_1099) );
INVx1_ASAP7_75t_L g1164 ( .A(n_159), .Y(n_1164) );
INVx1_ASAP7_75t_L g1749 ( .A(n_160), .Y(n_1749) );
INVx1_ASAP7_75t_L g1140 ( .A(n_162), .Y(n_1140) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_164), .Y(n_744) );
INVx1_ASAP7_75t_L g1387 ( .A(n_165), .Y(n_1387) );
AOI22xp33_ASAP7_75t_SL g999 ( .A1(n_166), .A2(n_215), .B1(n_710), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1265 ( .A(n_167), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g1082 ( .A1(n_168), .A2(n_283), .B1(n_550), .B2(n_1083), .Y(n_1082) );
INVx1_ASAP7_75t_L g1119 ( .A(n_169), .Y(n_1119) );
OAI211xp5_ASAP7_75t_L g1124 ( .A1(n_169), .A2(n_584), .B(n_1088), .C(n_1125), .Y(n_1124) );
CKINVDCx5p33_ASAP7_75t_R g1059 ( .A(n_170), .Y(n_1059) );
INVx1_ASAP7_75t_L g928 ( .A(n_172), .Y(n_928) );
OAI211xp5_ASAP7_75t_SL g1448 ( .A1(n_173), .A2(n_1149), .B(n_1449), .C(n_1451), .Y(n_1448) );
INVx1_ASAP7_75t_L g1463 ( .A(n_173), .Y(n_1463) );
INVx1_ASAP7_75t_L g1336 ( .A(n_175), .Y(n_1336) );
OAI211xp5_ASAP7_75t_L g1371 ( .A1(n_175), .A2(n_645), .B(n_793), .C(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g966 ( .A(n_176), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_178), .A2(n_271), .B1(n_990), .B2(n_991), .Y(n_989) );
OAI211xp5_ASAP7_75t_L g1116 ( .A1(n_179), .A2(n_609), .B(n_771), .C(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1126 ( .A(n_179), .Y(n_1126) );
INVx1_ASAP7_75t_L g1488 ( .A(n_180), .Y(n_1488) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_181), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g970 ( .A(n_182), .Y(n_970) );
OAI22xp33_ASAP7_75t_L g1120 ( .A1(n_184), .A2(n_186), .B1(n_550), .B2(n_1083), .Y(n_1120) );
OAI22xp33_ASAP7_75t_L g1123 ( .A1(n_184), .A2(n_196), .B1(n_510), .B2(n_795), .Y(n_1123) );
INVx1_ASAP7_75t_L g1142 ( .A(n_185), .Y(n_1142) );
OAI211xp5_ASAP7_75t_L g1146 ( .A1(n_185), .A2(n_1147), .B(n_1149), .C(n_1150), .Y(n_1146) );
OAI211xp5_ASAP7_75t_L g1040 ( .A1(n_187), .A2(n_584), .B(n_677), .C(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1049 ( .A(n_187), .Y(n_1049) );
INVx1_ASAP7_75t_L g1349 ( .A(n_188), .Y(n_1349) );
OAI22xp33_ASAP7_75t_SL g781 ( .A1(n_189), .A2(n_308), .B1(n_524), .B2(n_552), .Y(n_781) );
INVx1_ASAP7_75t_L g1345 ( .A(n_190), .Y(n_1345) );
INVx2_ASAP7_75t_L g1519 ( .A(n_192), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_192), .B(n_302), .Y(n_1521) );
AND2x2_ASAP7_75t_L g1527 ( .A(n_192), .B(n_1525), .Y(n_1527) );
AOI22xp5_ASAP7_75t_L g1536 ( .A1(n_193), .A2(n_282), .B1(n_1523), .B2(n_1526), .Y(n_1536) );
AO22x2_ASAP7_75t_L g1741 ( .A1(n_193), .A2(n_1742), .B1(n_1781), .B2(n_1782), .Y(n_1741) );
INVx1_ASAP7_75t_L g1781 ( .A(n_193), .Y(n_1781) );
AOI22xp33_ASAP7_75t_L g1786 ( .A1(n_193), .A2(n_1787), .B1(n_1790), .B2(n_1793), .Y(n_1786) );
INVx1_ASAP7_75t_L g1357 ( .A(n_195), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_197), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_198), .Y(n_810) );
INVx1_ASAP7_75t_L g1323 ( .A(n_199), .Y(n_1323) );
INVx1_ASAP7_75t_L g1161 ( .A(n_201), .Y(n_1161) );
XNOR2xp5_ASAP7_75t_L g1421 ( .A(n_202), .B(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g1406 ( .A(n_203), .Y(n_1406) );
OAI211xp5_ASAP7_75t_L g1412 ( .A1(n_203), .A2(n_584), .B(n_1413), .C(n_1414), .Y(n_1412) );
AOI22xp5_ASAP7_75t_L g1547 ( .A1(n_204), .A2(n_311), .B1(n_1516), .B2(n_1530), .Y(n_1547) );
INVx1_ASAP7_75t_L g871 ( .A(n_205), .Y(n_871) );
XOR2xp5_ASAP7_75t_L g916 ( .A(n_206), .B(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g508 ( .A(n_207), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g549 ( .A1(n_207), .A2(n_242), .B1(n_550), .B2(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g922 ( .A(n_208), .Y(n_922) );
CKINVDCx5p33_ASAP7_75t_R g1065 ( .A(n_209), .Y(n_1065) );
INVx1_ASAP7_75t_L g1298 ( .A(n_210), .Y(n_1298) );
INVx1_ASAP7_75t_L g1198 ( .A(n_211), .Y(n_1198) );
XOR2x2_ASAP7_75t_L g1192 ( .A(n_214), .B(n_1193), .Y(n_1192) );
AOI22xp33_ASAP7_75t_SL g1010 ( .A1(n_215), .A2(n_289), .B1(n_1004), .B2(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1432 ( .A(n_216), .Y(n_1432) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_218), .Y(n_569) );
OAI211xp5_ASAP7_75t_L g850 ( .A1(n_219), .A2(n_851), .B(n_852), .C(n_862), .Y(n_850) );
INVx1_ASAP7_75t_L g894 ( .A(n_219), .Y(n_894) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_220), .A2(n_244), .B1(n_579), .B2(n_1417), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1480 ( .A1(n_220), .A2(n_244), .B1(n_523), .B2(n_527), .Y(n_1480) );
INVx1_ASAP7_75t_L g925 ( .A(n_221), .Y(n_925) );
INVx2_ASAP7_75t_L g403 ( .A(n_222), .Y(n_403) );
INVx1_ASAP7_75t_L g442 ( .A(n_222), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_223), .Y(n_1060) );
XNOR2xp5_ASAP7_75t_L g1326 ( .A(n_225), .B(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g446 ( .A(n_228), .Y(n_446) );
INVx1_ASAP7_75t_L g1028 ( .A(n_229), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g1549 ( .A1(n_230), .A2(n_315), .B1(n_1523), .B2(n_1526), .Y(n_1549) );
INVx1_ASAP7_75t_L g861 ( .A(n_231), .Y(n_861) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_231), .A2(n_262), .B1(n_505), .B2(n_513), .Y(n_892) );
INVx1_ASAP7_75t_L g853 ( .A(n_233), .Y(n_853) );
INVx1_ASAP7_75t_L g490 ( .A(n_234), .Y(n_490) );
OA211x2_ASAP7_75t_L g531 ( .A1(n_234), .A2(n_532), .B(n_535), .C(n_540), .Y(n_531) );
BUFx3_ASAP7_75t_L g409 ( .A(n_235), .Y(n_409) );
INVx1_ASAP7_75t_L g1022 ( .A(n_236), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g1069 ( .A(n_237), .Y(n_1069) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_238), .Y(n_613) );
CKINVDCx5p33_ASAP7_75t_R g1109 ( .A(n_239), .Y(n_1109) );
OAI22xp5_ASAP7_75t_SL g393 ( .A1(n_240), .A2(n_394), .B1(n_520), .B2(n_561), .Y(n_393) );
NAND4xp25_ASAP7_75t_L g394 ( .A(n_240), .B(n_395), .C(n_449), .D(n_480), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g1295 ( .A1(n_241), .A2(n_349), .B1(n_377), .B2(n_552), .Y(n_1295) );
OAI22xp33_ASAP7_75t_L g1302 ( .A1(n_241), .A2(n_349), .B1(n_591), .B2(n_1270), .Y(n_1302) );
INVx1_ASAP7_75t_L g499 ( .A(n_242), .Y(n_499) );
INVx1_ASAP7_75t_L g1299 ( .A(n_243), .Y(n_1299) );
OAI211xp5_ASAP7_75t_L g1303 ( .A1(n_243), .A2(n_793), .B(n_1304), .C(n_1305), .Y(n_1303) );
OA22x2_ASAP7_75t_L g1466 ( .A1(n_245), .A2(n_1467), .B1(n_1504), .B2(n_1505), .Y(n_1466) );
INVxp67_ASAP7_75t_L g1505 ( .A(n_245), .Y(n_1505) );
INVx1_ASAP7_75t_L g670 ( .A(n_246), .Y(n_670) );
INVx1_ASAP7_75t_L g571 ( .A(n_247), .Y(n_571) );
OAI211xp5_ASAP7_75t_L g581 ( .A1(n_247), .A2(n_582), .B(n_584), .C(n_585), .Y(n_581) );
INVx1_ASAP7_75t_L g1264 ( .A(n_248), .Y(n_1264) );
INVx1_ASAP7_75t_L g866 ( .A(n_249), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_249), .B(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g1770 ( .A(n_250), .Y(n_1770) );
INVx1_ASAP7_75t_L g427 ( .A(n_251), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_252), .Y(n_1102) );
CKINVDCx5p33_ASAP7_75t_R g1062 ( .A(n_253), .Y(n_1062) );
AOI22xp5_ASAP7_75t_L g1542 ( .A1(n_254), .A2(n_275), .B1(n_1516), .B2(n_1520), .Y(n_1542) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_255), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g1012 ( .A1(n_256), .A2(n_271), .B1(n_721), .B2(n_1006), .C(n_1013), .Y(n_1012) );
INVx1_ASAP7_75t_L g676 ( .A(n_257), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_257), .A2(n_304), .B1(n_707), .B2(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g1746 ( .A(n_258), .Y(n_1746) );
INVx1_ASAP7_75t_L g1027 ( .A(n_259), .Y(n_1027) );
XOR2xp5_ASAP7_75t_L g797 ( .A(n_260), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1218 ( .A(n_261), .Y(n_1218) );
INVx1_ASAP7_75t_L g863 ( .A(n_262), .Y(n_863) );
BUFx3_ASAP7_75t_L g385 ( .A(n_263), .Y(n_385) );
INVx1_ASAP7_75t_L g526 ( .A(n_263), .Y(n_526) );
XOR2x2_ASAP7_75t_L g1130 ( .A(n_264), .B(n_1131), .Y(n_1130) );
INVx1_ASAP7_75t_L g485 ( .A(n_266), .Y(n_485) );
INVx1_ASAP7_75t_L g921 ( .A(n_267), .Y(n_921) );
INVx1_ASAP7_75t_L g448 ( .A(n_268), .Y(n_448) );
INVx1_ASAP7_75t_L g1214 ( .A(n_269), .Y(n_1214) );
XNOR2x1_ASAP7_75t_L g1278 ( .A(n_270), .B(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1285 ( .A(n_272), .Y(n_1285) );
OAI211xp5_ASAP7_75t_L g1330 ( .A1(n_273), .A2(n_1331), .B(n_1332), .C(n_1333), .Y(n_1330) );
INVx1_ASAP7_75t_L g1373 ( .A(n_273), .Y(n_1373) );
AOI22xp33_ASAP7_75t_L g1286 ( .A1(n_276), .A2(n_353), .B1(n_943), .B2(n_1287), .Y(n_1286) );
INVxp33_ASAP7_75t_SL g1314 ( .A(n_276), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g747 ( .A(n_277), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_279), .B(n_513), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g815 ( .A(n_281), .Y(n_815) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_283), .A2(n_299), .B1(n_510), .B2(n_795), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_284), .Y(n_751) );
INVx1_ASAP7_75t_L g436 ( .A(n_285), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_286), .Y(n_1100) );
XOR2x2_ASAP7_75t_L g1231 ( .A(n_287), .B(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1262 ( .A(n_288), .Y(n_1262) );
INVx1_ASAP7_75t_L g411 ( .A(n_290), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_290), .Y(n_418) );
OAI22xp33_ASAP7_75t_L g1300 ( .A1(n_291), .A2(n_340), .B1(n_573), .B2(n_574), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g1307 ( .A1(n_291), .A2(n_340), .B1(n_1308), .B2(n_1310), .Y(n_1307) );
INVx1_ASAP7_75t_L g432 ( .A(n_292), .Y(n_432) );
INVx1_ASAP7_75t_L g1289 ( .A(n_293), .Y(n_1289) );
INVx1_ASAP7_75t_L g671 ( .A(n_294), .Y(n_671) );
INVx1_ASAP7_75t_L g776 ( .A(n_295), .Y(n_776) );
OAI211xp5_ASAP7_75t_SL g784 ( .A1(n_295), .A2(n_723), .B(n_785), .C(n_793), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g575 ( .A1(n_296), .A2(n_297), .B1(n_377), .B2(n_552), .Y(n_575) );
OAI22xp33_ASAP7_75t_L g588 ( .A1(n_296), .A2(n_297), .B1(n_589), .B2(n_591), .Y(n_588) );
INVx1_ASAP7_75t_L g1167 ( .A(n_298), .Y(n_1167) );
INVx1_ASAP7_75t_L g924 ( .A(n_300), .Y(n_924) );
INVx1_ASAP7_75t_L g976 ( .A(n_301), .Y(n_976) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_302), .B(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1525 ( .A(n_302), .Y(n_1525) );
INVx1_ASAP7_75t_L g656 ( .A(n_304), .Y(n_656) );
INVx1_ASAP7_75t_L g1030 ( .A(n_305), .Y(n_1030) );
INVx1_ASAP7_75t_L g1215 ( .A(n_306), .Y(n_1215) );
CKINVDCx5p33_ASAP7_75t_R g1063 ( .A(n_307), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_308), .A2(n_346), .B1(n_505), .B2(n_513), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g597 ( .A(n_309), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_310), .A2(n_345), .B1(n_1523), .B2(n_1526), .Y(n_1565) );
INVx1_ASAP7_75t_L g1223 ( .A(n_312), .Y(n_1223) );
INVx1_ASAP7_75t_L g682 ( .A(n_313), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g1118 ( .A(n_314), .Y(n_1118) );
INVx1_ASAP7_75t_L g1756 ( .A(n_316), .Y(n_1756) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_317), .Y(n_873) );
OAI211xp5_ASAP7_75t_SL g831 ( .A1(n_318), .A2(n_770), .B(n_771), .C(n_832), .Y(n_831) );
OAI211xp5_ASAP7_75t_SL g842 ( .A1(n_318), .A2(n_793), .B(n_843), .C(n_844), .Y(n_842) );
INVx1_ASAP7_75t_L g1025 ( .A(n_319), .Y(n_1025) );
INVx1_ASAP7_75t_L g1453 ( .A(n_320), .Y(n_1453) );
OAI211xp5_ASAP7_75t_SL g1459 ( .A1(n_320), .A2(n_793), .B(n_1460), .C(n_1462), .Y(n_1459) );
INVx1_ASAP7_75t_L g945 ( .A(n_321), .Y(n_945) );
INVx1_ASAP7_75t_L g1290 ( .A(n_322), .Y(n_1290) );
INVx1_ASAP7_75t_L g1354 ( .A(n_323), .Y(n_1354) );
OAI211xp5_ASAP7_75t_L g565 ( .A1(n_326), .A2(n_535), .B(n_566), .C(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g587 ( .A(n_326), .Y(n_587) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_328), .A2(n_535), .B(n_826), .C(n_1404), .Y(n_1403) );
INVx1_ASAP7_75t_L g1415 ( .A(n_328), .Y(n_1415) );
AOI22xp33_ASAP7_75t_SL g1249 ( .A1(n_330), .A2(n_358), .B1(n_1250), .B2(n_1253), .Y(n_1249) );
INVx1_ASAP7_75t_L g1342 ( .A(n_331), .Y(n_1342) );
INVx1_ASAP7_75t_L g1485 ( .A(n_332), .Y(n_1485) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_333), .Y(n_754) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_334), .Y(n_601) );
INVx1_ASAP7_75t_L g412 ( .A(n_335), .Y(n_412) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_336), .Y(n_381) );
INVx1_ASAP7_75t_L g1750 ( .A(n_337), .Y(n_1750) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_338), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g1080 ( .A(n_339), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g777 ( .A(n_342), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g805 ( .A(n_343), .Y(n_805) );
INVx1_ASAP7_75t_L g1772 ( .A(n_344), .Y(n_1772) );
XOR2x2_ASAP7_75t_L g562 ( .A(n_345), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g401 ( .A(n_347), .Y(n_401) );
INVx2_ASAP7_75t_L g440 ( .A(n_347), .Y(n_440) );
INVx1_ASAP7_75t_L g641 ( .A(n_347), .Y(n_641) );
INVx1_ASAP7_75t_L g1384 ( .A(n_348), .Y(n_1384) );
INVx1_ASAP7_75t_L g1348 ( .A(n_350), .Y(n_1348) );
INVx1_ASAP7_75t_L g1426 ( .A(n_351), .Y(n_1426) );
INVx1_ASAP7_75t_L g511 ( .A(n_352), .Y(n_511) );
INVxp67_ASAP7_75t_SL g1322 ( .A(n_353), .Y(n_1322) );
INVx1_ASAP7_75t_L g1429 ( .A(n_354), .Y(n_1429) );
AOI21xp33_ASAP7_75t_L g875 ( .A1(n_355), .A2(n_876), .B(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g898 ( .A(n_355), .Y(n_898) );
INVx1_ASAP7_75t_L g1175 ( .A(n_356), .Y(n_1175) );
INVx1_ASAP7_75t_L g493 ( .A(n_357), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g1070 ( .A(n_359), .Y(n_1070) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_360), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_386), .B(n_1507), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_371), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g1785 ( .A(n_365), .B(n_374), .Y(n_1785) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g1789 ( .A(n_367), .B(n_370), .Y(n_1789) );
INVx1_ASAP7_75t_L g1796 ( .A(n_367), .Y(n_1796) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g1799 ( .A(n_370), .B(n_1796), .Y(n_1799) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g558 ( .A(n_374), .B(n_559), .Y(n_558) );
AOI21xp5_ASAP7_75t_SL g849 ( .A1(n_374), .A2(n_850), .B(n_864), .Y(n_849) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g476 ( .A(n_375), .B(n_385), .Y(n_476) );
AND2x4_ASAP7_75t_L g879 ( .A(n_375), .B(n_384), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_376), .A2(n_553), .B1(n_682), .B2(n_683), .Y(n_681) );
AND2x4_ASAP7_75t_SL g1784 ( .A(n_376), .B(n_1785), .Y(n_1784) );
INVx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_378), .B(n_383), .Y(n_377) );
BUFx4f_ASAP7_75t_L g457 ( .A(n_378), .Y(n_457) );
OR2x6_ASAP7_75t_L g524 ( .A(n_378), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g766 ( .A(n_378), .Y(n_766) );
OR2x2_ASAP7_75t_L g837 ( .A(n_378), .B(n_525), .Y(n_837) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g551 ( .A(n_379), .Y(n_551) );
BUFx4f_ASAP7_75t_L g600 ( .A(n_379), .Y(n_600) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx2_ASAP7_75t_L g461 ( .A(n_381), .Y(n_461) );
INVx2_ASAP7_75t_L g465 ( .A(n_381), .Y(n_465) );
NAND2x1_ASAP7_75t_L g469 ( .A(n_381), .B(n_382), .Y(n_469) );
AND2x2_ASAP7_75t_L g539 ( .A(n_381), .B(n_382), .Y(n_539) );
INVx1_ASAP7_75t_L g547 ( .A(n_381), .Y(n_547) );
AND2x2_ASAP7_75t_L g554 ( .A(n_381), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_382), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g464 ( .A(n_382), .B(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g542 ( .A(n_382), .Y(n_542) );
INVx2_ASAP7_75t_L g555 ( .A(n_382), .Y(n_555) );
INVx1_ASAP7_75t_L g696 ( .A(n_382), .Y(n_696) );
AND2x2_ASAP7_75t_L g711 ( .A(n_382), .B(n_461), .Y(n_711) );
OR2x6_ASAP7_75t_L g550 ( .A(n_383), .B(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_383), .A2(n_859), .B1(n_860), .B2(n_861), .Y(n_858) );
INVxp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g537 ( .A(n_384), .Y(n_537) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g530 ( .A(n_385), .Y(n_530) );
AND2x4_ASAP7_75t_L g545 ( .A(n_385), .B(n_546), .Y(n_545) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B1(n_1188), .B2(n_1506), .Y(n_386) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
XNOR2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_730), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_649), .B2(n_729), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_562), .B1(n_647), .B2(n_648), .Y(n_391) );
INVx1_ASAP7_75t_L g647 ( .A(n_392), .Y(n_647) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR4xp25_ASAP7_75t_L g561 ( .A(n_396), .B(n_450), .C(n_481), .D(n_520), .Y(n_561) );
OAI33xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_405), .A3(n_421), .B1(n_433), .B2(n_438), .B3(n_444), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_397), .A2(n_897), .B1(n_909), .B2(n_910), .Y(n_896) );
OAI33xp33_ASAP7_75t_L g919 ( .A1(n_397), .A2(n_438), .A3(n_920), .B1(n_923), .B2(n_926), .B3(n_930), .Y(n_919) );
OAI33xp33_ASAP7_75t_L g1158 ( .A1(n_397), .A2(n_909), .A3(n_1159), .B1(n_1163), .B2(n_1168), .B3(n_1174), .Y(n_1158) );
OAI33xp33_ASAP7_75t_L g1437 ( .A1(n_397), .A2(n_909), .A3(n_1438), .B1(n_1440), .B2(n_1442), .B3(n_1444), .Y(n_1437) );
OAI33xp33_ASAP7_75t_L g1498 ( .A1(n_397), .A2(n_637), .A3(n_1499), .B1(n_1501), .B2(n_1502), .B3(n_1503), .Y(n_1498) );
OAI33xp33_ASAP7_75t_L g1758 ( .A1(n_397), .A2(n_438), .A3(n_1759), .B1(n_1760), .B2(n_1761), .B3(n_1764), .Y(n_1758) );
BUFx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx8_ASAP7_75t_L g623 ( .A(n_398), .Y(n_623) );
BUFx4f_ASAP7_75t_L g654 ( .A(n_398), .Y(n_654) );
OR2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_402), .Y(n_398) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_399), .B(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_399), .Y(n_519) );
INVx1_ASAP7_75t_L g618 ( .A(n_399), .Y(n_618) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g560 ( .A(n_400), .Y(n_560) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_404), .Y(n_402) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_403), .Y(n_517) );
AND3x4_ASAP7_75t_L g1014 ( .A(n_403), .B(n_488), .C(n_1015), .Y(n_1014) );
INVx3_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
BUFx3_ASAP7_75t_L g488 ( .A(n_404), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_412), .B1(n_413), .B2(n_420), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_SL g659 ( .A(n_407), .Y(n_659) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx3_ASAP7_75t_L g445 ( .A(n_408), .Y(n_445) );
OR2x4_ASAP7_75t_L g510 ( .A(n_408), .B(n_443), .Y(n_510) );
OR2x4_ASAP7_75t_L g513 ( .A(n_408), .B(n_501), .Y(n_513) );
BUFx3_ASAP7_75t_L g627 ( .A(n_408), .Y(n_627) );
BUFx4f_ASAP7_75t_L g741 ( .A(n_408), .Y(n_741) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_409), .Y(n_419) );
INVx2_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_409), .B(n_418), .Y(n_431) );
AND2x4_ASAP7_75t_L g495 ( .A(n_409), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g904 ( .A(n_410), .Y(n_904) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_412), .A2(n_446), .B1(n_457), .B2(n_458), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_413), .A2(n_741), .B1(n_802), .B2(n_803), .Y(n_801) );
OAI22xp5_ASAP7_75t_SL g1023 ( .A1(n_413), .A2(n_741), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1058 ( .A1(n_413), .A2(n_741), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
OAI22xp33_ASAP7_75t_L g1759 ( .A1(n_413), .A2(n_741), .B1(n_1749), .B2(n_1756), .Y(n_1759) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g628 ( .A(n_414), .Y(n_628) );
INVx2_ASAP7_75t_L g1162 ( .A(n_414), .Y(n_1162) );
INVx3_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
INVx4_ASAP7_75t_L g646 ( .A(n_415), .Y(n_646) );
HB1xp67_ASAP7_75t_L g1439 ( .A(n_415), .Y(n_1439) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx3_ASAP7_75t_L g678 ( .A(n_416), .Y(n_678) );
BUFx2_ASAP7_75t_L g1090 ( .A(n_416), .Y(n_1090) );
NAND2x1p5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
BUFx2_ASAP7_75t_L g492 ( .A(n_417), .Y(n_492) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g496 ( .A(n_418), .Y(n_496) );
BUFx2_ASAP7_75t_L g489 ( .A(n_419), .Y(n_489) );
INVx2_ASAP7_75t_L g790 ( .A(n_419), .Y(n_790) );
AND2x4_ASAP7_75t_L g908 ( .A(n_419), .B(n_788), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_420), .A2(n_448), .B1(n_466), .B2(n_471), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_427), .B1(n_428), .B2(n_432), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g911 ( .A(n_423), .Y(n_911) );
INVx3_ASAP7_75t_L g1011 ( .A(n_423), .Y(n_1011) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx8_ASAP7_75t_L g435 ( .A(n_424), .Y(n_435) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_424), .Y(n_502) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_424), .Y(n_664) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AND2x4_ASAP7_75t_L g903 ( .A(n_426), .B(n_904), .Y(n_903) );
OAI22xp5_ASAP7_75t_SL g462 ( .A1(n_427), .A2(n_436), .B1(n_463), .B2(n_466), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g433 ( .A1(n_428), .A2(n_434), .B1(n_436), .B2(n_437), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_428), .A2(n_669), .B1(n_670), .B2(n_671), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_428), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
OAI22xp5_ASAP7_75t_L g923 ( .A1(n_428), .A2(n_911), .B1(n_924), .B2(n_925), .Y(n_923) );
OAI22xp5_ASAP7_75t_L g1219 ( .A1(n_428), .A2(n_745), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
BUFx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g1763 ( .A(n_429), .Y(n_1763) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_430), .Y(n_667) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g506 ( .A(n_431), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_432), .A2(n_437), .B1(n_457), .B2(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_SL g669 ( .A(n_435), .Y(n_669) );
INVx2_ASAP7_75t_SL g745 ( .A(n_435), .Y(n_745) );
INVx3_ASAP7_75t_L g927 ( .A(n_435), .Y(n_927) );
INVx1_ASAP7_75t_L g1009 ( .A(n_438), .Y(n_1009) );
OR2x6_ASAP7_75t_L g438 ( .A(n_439), .B(n_441), .Y(n_438) );
AND2x4_ASAP7_75t_L g454 ( .A(n_439), .B(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g755 ( .A(n_439), .B(n_441), .Y(n_755) );
INVx1_ASAP7_75t_L g884 ( .A(n_439), .Y(n_884) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g1015 ( .A(n_440), .Y(n_1015) );
NAND2x1p5_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
NAND3x1_ASAP7_75t_L g639 ( .A(n_442), .B(n_443), .C(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g497 ( .A(n_443), .B(n_495), .Y(n_497) );
INVx1_ASAP7_75t_L g501 ( .A(n_443), .Y(n_501) );
OR2x6_ASAP7_75t_L g505 ( .A(n_443), .B(n_506), .Y(n_505) );
OAI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_444) );
OAI22xp33_ASAP7_75t_L g1159 ( .A1(n_445), .A2(n_1160), .B1(n_1161), .B2(n_1162), .Y(n_1159) );
OAI22xp33_ASAP7_75t_L g1174 ( .A1(n_445), .A2(n_1088), .B1(n_1175), .B2(n_1176), .Y(n_1174) );
OAI22xp33_ASAP7_75t_L g1356 ( .A1(n_445), .A2(n_677), .B1(n_1357), .B2(n_1358), .Y(n_1356) );
OAI22xp33_ASAP7_75t_L g1438 ( .A1(n_445), .A2(n_1426), .B1(n_1432), .B2(n_1439), .Y(n_1438) );
OAI22xp33_ASAP7_75t_L g1444 ( .A1(n_445), .A2(n_1427), .B1(n_1433), .B2(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g583 ( .A(n_447), .Y(n_583) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_447), .A2(n_656), .B1(n_657), .B2(n_660), .Y(n_655) );
OAI22xp33_ASAP7_75t_L g739 ( .A1(n_447), .A2(n_740), .B1(n_741), .B2(n_742), .Y(n_739) );
OAI22xp33_ASAP7_75t_L g930 ( .A1(n_447), .A2(n_741), .B1(n_931), .B2(n_932), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g1111 ( .A1(n_447), .A2(n_659), .B1(n_1099), .B2(n_1105), .Y(n_1111) );
OAI22xp33_ASAP7_75t_L g1213 ( .A1(n_447), .A2(n_741), .B1(n_1214), .B2(n_1215), .Y(n_1213) );
OAI22xp33_ASAP7_75t_L g1503 ( .A1(n_447), .A2(n_625), .B1(n_1486), .B2(n_1492), .Y(n_1503) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI33xp33_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_456), .A3(n_462), .B1(n_470), .B2(n_474), .B3(n_477), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g988 ( .A(n_453), .Y(n_988) );
OAI33xp33_ASAP7_75t_L g1382 ( .A1(n_453), .A2(n_615), .A3(n_1383), .B1(n_1386), .B2(n_1390), .B3(n_1393), .Y(n_1382) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g604 ( .A(n_454), .Y(n_604) );
INVx2_ASAP7_75t_L g703 ( .A(n_454), .Y(n_703) );
INVx2_ASAP7_75t_L g818 ( .A(n_454), .Y(n_818) );
INVx2_ASAP7_75t_L g1178 ( .A(n_454), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g865 ( .A1(n_457), .A2(n_866), .B1(n_867), .B2(n_868), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g1313 ( .A1(n_457), .A2(n_868), .B1(n_1314), .B2(n_1315), .Y(n_1313) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx8_ASAP7_75t_L g479 ( .A(n_459), .Y(n_479) );
OR2x2_ASAP7_75t_L g529 ( .A(n_459), .B(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g830 ( .A(n_459), .B(n_537), .Y(n_830) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g1035 ( .A1(n_463), .A2(n_824), .B1(n_1021), .B2(n_1030), .Y(n_1035) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_463), .A2(n_534), .B1(n_1060), .B2(n_1070), .Y(n_1075) );
BUFx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g473 ( .A(n_464), .Y(n_473) );
INVx1_ASAP7_75t_L g608 ( .A(n_464), .Y(n_608) );
BUFx3_ASAP7_75t_L g715 ( .A(n_464), .Y(n_715) );
BUFx2_ASAP7_75t_L g1319 ( .A(n_464), .Y(n_1319) );
AND2x2_ASAP7_75t_L g695 ( .A(n_465), .B(n_696), .Y(n_695) );
OAI221xp5_ASAP7_75t_L g869 ( .A1(n_466), .A2(n_471), .B1(n_476), .B2(n_870), .C(n_871), .Y(n_869) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g609 ( .A(n_467), .Y(n_609) );
INVx2_ASAP7_75t_L g762 ( .A(n_467), .Y(n_762) );
INVx2_ASAP7_75t_L g826 ( .A(n_467), .Y(n_826) );
INVx2_ASAP7_75t_L g1184 ( .A(n_467), .Y(n_1184) );
INVx4_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx4f_ASAP7_75t_L g614 ( .A(n_468), .Y(n_614) );
BUFx4f_ASAP7_75t_L g770 ( .A(n_468), .Y(n_770) );
BUFx4f_ASAP7_75t_L g824 ( .A(n_468), .Y(n_824) );
BUFx4f_ASAP7_75t_L g874 ( .A(n_468), .Y(n_874) );
BUFx6f_ASAP7_75t_L g937 ( .A(n_468), .Y(n_937) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx3_ASAP7_75t_L g534 ( .A(n_469), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g1183 ( .A1(n_471), .A2(n_1164), .B1(n_1171), .B2(n_1184), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1185 ( .A1(n_471), .A2(n_609), .B1(n_1161), .B2(n_1176), .Y(n_1185) );
OAI22xp5_ASAP7_75t_L g1321 ( .A1(n_471), .A2(n_770), .B1(n_1322), .B2(n_1323), .Y(n_1321) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g705 ( .A(n_473), .Y(n_705) );
INVx2_ASAP7_75t_L g1074 ( .A(n_473), .Y(n_1074) );
OAI33xp33_ASAP7_75t_L g1071 ( .A1(n_474), .A2(n_703), .A3(n_1072), .B1(n_1073), .B2(n_1075), .B3(n_1076), .Y(n_1071) );
OAI33xp33_ASAP7_75t_L g1097 ( .A1(n_474), .A2(n_818), .A3(n_1098), .B1(n_1101), .B2(n_1104), .B3(n_1107), .Y(n_1097) );
OAI33xp33_ASAP7_75t_L g1744 ( .A1(n_474), .A2(n_1745), .A3(n_1748), .B1(n_1751), .B2(n_1752), .B3(n_1755), .Y(n_1744) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g767 ( .A(n_475), .Y(n_767) );
AOI33xp33_ASAP7_75t_L g987 ( .A1(n_475), .A2(n_988), .A3(n_989), .B1(n_993), .B2(n_997), .B3(n_999), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g1242 ( .A(n_475), .B(n_1243), .C(n_1244), .Y(n_1242) );
AND2x4_ASAP7_75t_L g616 ( .A(n_476), .B(n_617), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_478), .A2(n_758), .B1(n_1099), .B2(n_1100), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g1383 ( .A1(n_478), .A2(n_598), .B1(n_1384), .B2(n_1385), .Y(n_1383) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_479), .Y(n_603) );
INVx4_ASAP7_75t_L g759 ( .A(n_479), .Y(n_759) );
INVx2_ASAP7_75t_L g822 ( .A(n_479), .Y(n_822) );
INVx1_ASAP7_75t_L g1034 ( .A(n_479), .Y(n_1034) );
INVx1_ASAP7_75t_L g1227 ( .A(n_479), .Y(n_1227) );
INVx2_ASAP7_75t_L g1395 ( .A(n_479), .Y(n_1395) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AOI31xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_498), .A3(n_507), .B(n_514), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_497), .Y(n_482) );
INVxp67_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_486), .B1(n_490), .B2(n_491), .C1(n_493), .C2(n_494), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_485), .A2(n_493), .B1(n_541), .B2(n_543), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_486), .A2(n_786), .B1(n_833), .B2(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g890 ( .A(n_486), .Y(n_890) );
AOI222xp33_ASAP7_75t_L g942 ( .A1(n_486), .A2(n_791), .B1(n_943), .B2(n_944), .C1(n_945), .C2(n_946), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g983 ( .A(n_486), .B(n_970), .Y(n_983) );
AOI22xp33_ASAP7_75t_SL g1041 ( .A1(n_486), .A2(n_791), .B1(n_1042), .B2(n_1043), .Y(n_1041) );
AOI22xp33_ASAP7_75t_SL g1091 ( .A1(n_486), .A2(n_791), .B1(n_1080), .B2(n_1092), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g1125 ( .A1(n_486), .A2(n_791), .B1(n_1118), .B2(n_1126), .Y(n_1125) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_489), .Y(n_486) );
AND2x4_ASAP7_75t_L g491 ( .A(n_487), .B(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g586 ( .A(n_487), .B(n_489), .Y(n_586) );
AND2x2_ASAP7_75t_L g791 ( .A(n_487), .B(n_492), .Y(n_791) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_487), .B(n_489), .Y(n_1139) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g786 ( .A(n_488), .B(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_491), .A2(n_569), .B1(n_586), .B2(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g724 ( .A(n_491), .Y(n_724) );
BUFx6f_ASAP7_75t_L g1141 ( .A(n_491), .Y(n_1141) );
AOI222xp33_ASAP7_75t_L g1272 ( .A1(n_491), .A2(n_494), .B1(n_1264), .B2(n_1265), .C1(n_1266), .C2(n_1273), .Y(n_1272) );
AOI22xp33_ASAP7_75t_L g1414 ( .A1(n_491), .A2(n_586), .B1(n_1405), .B2(n_1415), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_491), .A2(n_586), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g1778 ( .A1(n_491), .A2(n_586), .B1(n_1769), .B2(n_1772), .Y(n_1778) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx3_ASAP7_75t_L g721 ( .A(n_495), .Y(n_721) );
BUFx2_ASAP7_75t_L g905 ( .A(n_495), .Y(n_905) );
BUFx2_ASAP7_75t_L g943 ( .A(n_495), .Y(n_943) );
INVx2_ASAP7_75t_L g1008 ( .A(n_495), .Y(n_1008) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_495), .Y(n_1293) );
INVx1_ASAP7_75t_L g788 ( .A(n_496), .Y(n_788) );
CKINVDCx8_ASAP7_75t_R g584 ( .A(n_497), .Y(n_584) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_497), .A2(n_720), .B(n_721), .C(n_722), .Y(n_719) );
CKINVDCx8_ASAP7_75t_R g793 ( .A(n_497), .Y(n_793) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_497), .B(n_888), .C(n_892), .Y(n_887) );
NOR3xp33_ASAP7_75t_L g980 ( .A(n_497), .B(n_981), .C(n_984), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_500), .B1(n_503), .B2(n_504), .Y(n_498) );
INVx2_ASAP7_75t_L g795 ( .A(n_500), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_500), .A2(n_590), .B1(n_859), .B2(n_894), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g979 ( .A1(n_500), .A2(n_726), .B1(n_964), .B2(n_966), .Y(n_979) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
AND2x4_ASAP7_75t_L g592 ( .A(n_501), .B(n_502), .Y(n_592) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_502), .Y(n_631) );
INVx2_ASAP7_75t_L g636 ( .A(n_502), .Y(n_636) );
INVx2_ASAP7_75t_L g806 ( .A(n_502), .Y(n_806) );
BUFx6f_ASAP7_75t_L g900 ( .A(n_502), .Y(n_900) );
INVx2_ASAP7_75t_L g1443 ( .A(n_502), .Y(n_1443) );
INVx1_ASAP7_75t_L g580 ( .A(n_504), .Y(n_580) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g728 ( .A(n_505), .Y(n_728) );
INVx1_ASAP7_75t_L g1309 ( .A(n_505), .Y(n_1309) );
BUFx3_ASAP7_75t_L g1417 ( .A(n_505), .Y(n_1417) );
INVx1_ASAP7_75t_L g634 ( .A(n_506), .Y(n_634) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_506), .Y(n_1172) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_509), .B1(n_511), .B2(n_512), .Y(n_507) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g590 ( .A(n_510), .Y(n_590) );
INVx2_ASAP7_75t_SL g726 ( .A(n_510), .Y(n_726) );
INVx2_ASAP7_75t_SL g1135 ( .A(n_510), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_512), .A2(n_692), .B1(n_697), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_512), .A2(n_728), .B1(n_1261), .B2(n_1262), .Y(n_1274) );
INVx2_ASAP7_75t_L g1310 ( .A(n_512), .Y(n_1310) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
BUFx3_ASAP7_75t_L g579 ( .A(n_513), .Y(n_579) );
BUFx2_ASAP7_75t_L g1458 ( .A(n_513), .Y(n_1458) );
AOI31xp33_ASAP7_75t_L g718 ( .A1(n_514), .A2(n_719), .A3(n_725), .B(n_727), .Y(n_718) );
CKINVDCx14_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
OAI31xp33_ASAP7_75t_L g1468 ( .A1(n_515), .A2(n_1469), .A3(n_1470), .B(n_1474), .Y(n_1468) );
AND2x4_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
AND2x2_ASAP7_75t_L g593 ( .A(n_516), .B(n_518), .Y(n_593) );
AND2x2_ASAP7_75t_L g796 ( .A(n_516), .B(n_518), .Y(n_796) );
AND2x2_ASAP7_75t_SL g895 ( .A(n_516), .B(n_518), .Y(n_895) );
AND2x2_ASAP7_75t_L g986 ( .A(n_516), .B(n_518), .Y(n_986) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI31xp67_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_531), .A3(n_548), .B(n_556), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g573 ( .A(n_524), .Y(n_573) );
AND2x4_ASAP7_75t_L g553 ( .A(n_525), .B(n_554), .Y(n_553) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g574 ( .A(n_528), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g1260 ( .A1(n_528), .A2(n_693), .B1(n_1261), .B2(n_1262), .Y(n_1260) );
INVxp67_ASAP7_75t_SL g1408 ( .A(n_528), .Y(n_1408) );
INVx1_ASAP7_75t_L g1774 ( .A(n_528), .Y(n_1774) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g700 ( .A(n_529), .Y(n_700) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_529), .Y(n_1083) );
AND2x4_ASAP7_75t_L g541 ( .A(n_530), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g568 ( .A(n_530), .B(n_542), .Y(n_568) );
AND2x2_ASAP7_75t_L g693 ( .A(n_530), .B(n_694), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g852 ( .A1(n_530), .A2(n_853), .B(n_854), .C(n_855), .Y(n_852) );
INVx1_ASAP7_75t_L g860 ( .A(n_530), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g1361 ( .A1(n_532), .A2(n_1317), .B1(n_1348), .B2(n_1351), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_532), .A2(n_1345), .B1(n_1358), .B2(n_1363), .Y(n_1362) );
OAI22xp5_ASAP7_75t_L g1390 ( .A1(n_532), .A2(n_607), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
OAI22xp5_ASAP7_75t_L g1428 ( .A1(n_532), .A2(n_1317), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_532), .A2(n_607), .B1(n_1488), .B2(n_1489), .Y(n_1487) );
INVx5_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
BUFx3_ASAP7_75t_L g566 ( .A(n_534), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_534), .A2(n_1074), .B1(n_1102), .B2(n_1103), .Y(n_1101) );
OAI22xp5_ASAP7_75t_L g1229 ( .A1(n_534), .A2(n_761), .B1(n_1215), .B2(n_1224), .Y(n_1229) );
BUFx2_ASAP7_75t_SL g1320 ( .A(n_534), .Y(n_1320) );
NAND3xp33_ASAP7_75t_L g1767 ( .A(n_535), .B(n_1768), .C(n_1771), .Y(n_1767) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_536), .A2(n_685), .B(n_688), .C(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g1149 ( .A(n_536), .Y(n_1149) );
INVx1_ASAP7_75t_L g1332 ( .A(n_536), .Y(n_1332) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AND2x2_ASAP7_75t_L g772 ( .A(n_537), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g857 ( .A(n_537), .B(n_542), .Y(n_857) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_538), .Y(n_687) );
BUFx3_ASAP7_75t_L g854 ( .A(n_538), .Y(n_854) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g774 ( .A(n_539), .Y(n_774) );
INVx1_ASAP7_75t_L g690 ( .A(n_541), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_541), .A2(n_833), .B1(n_834), .B2(n_835), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_541), .A2(n_835), .B1(n_1198), .B2(n_1199), .Y(n_1197) );
AOI222xp33_ASAP7_75t_L g1263 ( .A1(n_541), .A2(n_835), .B1(n_854), .B2(n_1264), .C1(n_1265), .C2(n_1266), .Y(n_1263) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_541), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g1404 ( .A1(n_541), .A2(n_778), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1150 ( .A1(n_543), .A2(n_568), .B1(n_1140), .B2(n_1151), .Y(n_1150) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g570 ( .A(n_544), .Y(n_570) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g779 ( .A(n_545), .Y(n_779) );
BUFx3_ASAP7_75t_L g835 ( .A(n_545), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_545), .A2(n_857), .B1(n_970), .B2(n_971), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_545), .A2(n_568), .B1(n_1298), .B2(n_1299), .Y(n_1297) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVxp67_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g965 ( .A(n_550), .Y(n_965) );
BUFx3_ASAP7_75t_L g820 ( .A(n_551), .Y(n_820) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_551), .Y(n_939) );
BUFx3_ASAP7_75t_L g1325 ( .A(n_551), .Y(n_1325) );
INVx2_ASAP7_75t_SL g1495 ( .A(n_551), .Y(n_1495) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
INVx4_ASAP7_75t_L g838 ( .A(n_553), .Y(n_838) );
INVx3_ASAP7_75t_SL g851 ( .A(n_553), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_553), .A2(n_964), .B1(n_965), .B2(n_966), .Y(n_963) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_554), .Y(n_877) );
BUFx3_ASAP7_75t_L g1238 ( .A(n_554), .Y(n_1238) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI31xp33_ASAP7_75t_L g768 ( .A1(n_557), .A2(n_769), .A3(n_780), .B(n_781), .Y(n_768) );
OAI31xp33_ASAP7_75t_SL g1045 ( .A1(n_557), .A2(n_1046), .A3(n_1047), .B(n_1050), .Y(n_1045) );
OAI31xp33_ASAP7_75t_L g1077 ( .A1(n_557), .A2(n_1078), .A3(n_1082), .B(n_1084), .Y(n_1077) );
OAI31xp33_ASAP7_75t_L g1115 ( .A1(n_557), .A2(n_1116), .A3(n_1120), .B(n_1121), .Y(n_1115) );
OAI31xp33_ASAP7_75t_SL g1294 ( .A1(n_557), .A2(n_1295), .A3(n_1296), .B(n_1300), .Y(n_1294) );
OAI31xp33_ASAP7_75t_L g1402 ( .A1(n_557), .A2(n_1403), .A3(n_1407), .B(n_1409), .Y(n_1402) );
OAI31xp33_ASAP7_75t_L g1765 ( .A1(n_557), .A2(n_1766), .A3(n_1767), .B(n_1773), .Y(n_1765) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx2_ASAP7_75t_SL g576 ( .A(n_558), .Y(n_576) );
INVx1_ASAP7_75t_L g701 ( .A(n_558), .Y(n_701) );
OAI31xp33_ASAP7_75t_L g828 ( .A1(n_558), .A2(n_829), .A3(n_831), .B(n_836), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g949 ( .A1(n_558), .A2(n_950), .B(n_957), .Y(n_949) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_558), .Y(n_1156) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g648 ( .A(n_562), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g563 ( .A(n_564), .B(n_577), .C(n_594), .Y(n_563) );
OAI31xp33_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_572), .A3(n_575), .B(n_576), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_566), .A2(n_662), .B1(n_670), .B2(n_705), .C(n_706), .Y(n_704) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_566), .A2(n_660), .B1(n_679), .B2(n_713), .C(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g1148 ( .A(n_566), .Y(n_1148) );
BUFx2_ASAP7_75t_L g1331 ( .A(n_566), .Y(n_1331) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B1(n_570), .B2(n_571), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g775 ( .A1(n_568), .A2(n_776), .B1(n_777), .B2(n_778), .Y(n_775) );
AOI222xp33_ASAP7_75t_L g951 ( .A1(n_568), .A2(n_835), .B1(n_854), .B2(n_945), .C1(n_946), .C2(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_568), .A2(n_778), .B1(n_1042), .B2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g1478 ( .A1(n_568), .A2(n_570), .B1(n_1472), .B2(n_1479), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g1768 ( .A1(n_568), .A2(n_835), .B1(n_1769), .B2(n_1770), .Y(n_1768) );
OAI31xp33_ASAP7_75t_SL g1194 ( .A1(n_576), .A2(n_1195), .A3(n_1200), .B(n_1201), .Y(n_1194) );
OAI21xp5_ASAP7_75t_L g1258 ( .A1(n_576), .A2(n_1259), .B(n_1267), .Y(n_1258) );
OAI31xp33_ASAP7_75t_L g1476 ( .A1(n_576), .A2(n_1477), .A3(n_1480), .B(n_1481), .Y(n_1476) );
OAI31xp33_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .A3(n_588), .B(n_593), .Y(n_577) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
NAND3xp33_ASAP7_75t_L g1205 ( .A(n_584), .B(n_1206), .C(n_1208), .Y(n_1205) );
INVx1_ASAP7_75t_L g723 ( .A(n_586), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_586), .A2(n_791), .B1(n_1198), .B2(n_1207), .Y(n_1206) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_592), .A2(n_682), .B1(n_683), .B2(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g1204 ( .A(n_592), .Y(n_1204) );
INVx1_ASAP7_75t_L g1475 ( .A(n_592), .Y(n_1475) );
OAI31xp33_ASAP7_75t_L g1410 ( .A1(n_593), .A2(n_1411), .A3(n_1412), .B(n_1416), .Y(n_1410) );
NOR2xp33_ASAP7_75t_SL g594 ( .A(n_595), .B(n_622), .Y(n_594) );
OAI33xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_604), .A3(n_605), .B1(n_611), .B2(n_615), .B3(n_619), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_601), .B2(n_602), .Y(n_596) );
OAI22xp33_ASAP7_75t_L g624 ( .A1(n_597), .A2(n_612), .B1(n_625), .B2(n_628), .Y(n_624) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_598), .A2(n_602), .B1(n_620), .B2(n_621), .Y(n_619) );
OAI22xp33_ASAP7_75t_L g1484 ( .A1(n_598), .A2(n_868), .B1(n_1485), .B2(n_1486), .Y(n_1484) );
INVx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g1366 ( .A(n_599), .Y(n_1366) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx4_ASAP7_75t_L g758 ( .A(n_600), .Y(n_758) );
INVx3_ASAP7_75t_L g1182 ( .A(n_600), .Y(n_1182) );
OAI22xp33_ASAP7_75t_L g642 ( .A1(n_601), .A2(n_613), .B1(n_643), .B2(n_645), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_602), .A2(n_1160), .B1(n_1175), .B2(n_1180), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1186 ( .A1(n_602), .A2(n_1167), .B1(n_1173), .B2(n_1180), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_602), .A2(n_1285), .B1(n_1290), .B2(n_1325), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1425 ( .A1(n_602), .A2(n_1325), .B1(n_1426), .B2(n_1427), .Y(n_1425) );
INVx6_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx5_ASAP7_75t_L g868 ( .A(n_603), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B1(n_609), .B2(n_610), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_606), .A2(n_620), .B1(n_630), .B2(n_632), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_607), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_607), .A2(n_922), .B1(n_932), .B2(n_937), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g1490 ( .A1(n_607), .A2(n_614), .B1(n_1491), .B2(n_1492), .Y(n_1490) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g761 ( .A(n_608), .Y(n_761) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_610), .A2(n_621), .B1(n_632), .B2(n_636), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g1386 ( .A1(n_614), .A2(n_1387), .B1(n_1388), .B2(n_1389), .Y(n_1386) );
INVx1_ASAP7_75t_L g1450 ( .A(n_614), .Y(n_1450) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_615), .A2(n_703), .B1(n_704), .B2(n_712), .Y(n_702) );
OAI33xp33_ASAP7_75t_L g1177 ( .A1(n_615), .A2(n_1178), .A3(n_1179), .B1(n_1183), .B2(n_1185), .B3(n_1186), .Y(n_1177) );
OA33x2_ASAP7_75t_L g1311 ( .A1(n_615), .A2(n_1312), .A3(n_1313), .B1(n_1316), .B2(n_1321), .B3(n_1324), .Y(n_1311) );
OAI33xp33_ASAP7_75t_L g1483 ( .A1(n_615), .A2(n_1178), .A3(n_1484), .B1(n_1487), .B2(n_1490), .B3(n_1493), .Y(n_1483) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g1368 ( .A(n_616), .Y(n_1368) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI33xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .A3(n_629), .B1(n_635), .B2(n_637), .B3(n_642), .Y(n_622) );
OAI33xp33_ASAP7_75t_L g1397 ( .A1(n_623), .A2(n_637), .A3(n_1398), .B1(n_1399), .B2(n_1400), .B3(n_1401), .Y(n_1397) );
OAI22xp33_ASAP7_75t_L g1398 ( .A1(n_625), .A2(n_1304), .B1(n_1384), .B2(n_1391), .Y(n_1398) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_625), .A2(n_628), .B1(n_1385), .B2(n_1392), .Y(n_1401) );
OAI22xp33_ASAP7_75t_L g1499 ( .A1(n_625), .A2(n_1485), .B1(n_1491), .B2(n_1500), .Y(n_1499) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g644 ( .A(n_627), .Y(n_644) );
INVxp67_ASAP7_75t_SL g1344 ( .A(n_627), .Y(n_1344) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g1441 ( .A(n_631), .Y(n_1441) );
INVx3_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g746 ( .A(n_634), .Y(n_746) );
OAI22xp33_ASAP7_75t_SL g1400 ( .A1(n_636), .A2(n_912), .B1(n_1389), .B2(n_1396), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1281 ( .A1(n_637), .A2(n_653), .B1(n_1282), .B2(n_1288), .Y(n_1281) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g909 ( .A(n_638), .Y(n_909) );
INVx2_ASAP7_75t_L g1355 ( .A(n_638), .Y(n_1355) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx3_ASAP7_75t_L g674 ( .A(n_639), .Y(n_674) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g889 ( .A(n_646), .Y(n_889) );
INVx1_ASAP7_75t_L g1304 ( .A(n_646), .Y(n_1304) );
INVx1_ASAP7_75t_L g1346 ( .A(n_646), .Y(n_1346) );
INVx1_ASAP7_75t_L g1413 ( .A(n_646), .Y(n_1413) );
INVx1_ASAP7_75t_L g729 ( .A(n_649), .Y(n_729) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NOR4xp25_ASAP7_75t_L g651 ( .A(n_652), .B(n_680), .C(n_702), .D(n_718), .Y(n_651) );
OAI33xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .A3(n_661), .B1(n_668), .B2(n_672), .B3(n_675), .Y(n_652) );
BUFx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OAI33xp33_ASAP7_75t_L g738 ( .A1(n_654), .A2(n_739), .A3(n_743), .B1(n_748), .B2(n_752), .B3(n_755), .Y(n_738) );
OAI33xp33_ASAP7_75t_L g800 ( .A1(n_654), .A2(n_755), .A3(n_801), .B1(n_804), .B2(n_809), .B3(n_814), .Y(n_800) );
OAI33xp33_ASAP7_75t_L g1019 ( .A1(n_654), .A2(n_755), .A3(n_1020), .B1(n_1023), .B2(n_1026), .B3(n_1029), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g1057 ( .A1(n_654), .A2(n_755), .A3(n_1058), .B1(n_1061), .B2(n_1064), .B3(n_1068), .Y(n_1057) );
OAI33xp33_ASAP7_75t_L g1110 ( .A1(n_654), .A2(n_755), .A3(n_1111), .B1(n_1112), .B2(n_1113), .B3(n_1114), .Y(n_1110) );
OAI33xp33_ASAP7_75t_L g1212 ( .A1(n_654), .A2(n_755), .A3(n_1213), .B1(n_1216), .B2(n_1219), .B3(n_1222), .Y(n_1212) );
OAI33xp33_ASAP7_75t_L g1340 ( .A1(n_654), .A2(n_1341), .A3(n_1347), .B1(n_1350), .B2(n_1355), .B3(n_1356), .Y(n_1340) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_659), .A2(n_676), .B1(n_677), .B2(n_679), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g1068 ( .A1(n_659), .A2(n_678), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
OAI22xp33_ASAP7_75t_L g1114 ( .A1(n_659), .A2(n_678), .B1(n_1100), .B2(n_1106), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_665), .B2(n_666), .Y(n_661) );
INVx2_ASAP7_75t_L g1003 ( .A(n_663), .Y(n_1003) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g749 ( .A(n_664), .Y(n_749) );
INVx2_ASAP7_75t_SL g811 ( .A(n_664), .Y(n_811) );
INVx5_ASAP7_75t_L g1166 ( .A(n_664), .Y(n_1166) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_664), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g926 ( .A1(n_666), .A2(n_927), .B1(n_928), .B2(n_929), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_666), .A2(n_811), .B1(n_1103), .B2(n_1109), .Y(n_1113) );
INVx3_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx3_ASAP7_75t_L g808 ( .A(n_667), .Y(n_808) );
INVx3_ASAP7_75t_L g813 ( .A(n_667), .Y(n_813) );
CKINVDCx8_ASAP7_75t_R g912 ( .A(n_667), .Y(n_912) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_674), .Y(n_1256) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_678), .A2(n_741), .B1(n_753), .B2(n_754), .Y(n_752) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_678), .A2(n_741), .B1(n_815), .B2(n_816), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g1026 ( .A1(n_678), .A2(n_741), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp33_ASAP7_75t_L g1222 ( .A1(n_678), .A2(n_741), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
OAI22xp33_ASAP7_75t_L g1764 ( .A1(n_678), .A2(n_741), .B1(n_1750), .B2(n_1757), .Y(n_1764) );
AOI31xp33_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_684), .A3(n_691), .B(n_701), .Y(n_680) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_697), .B2(n_698), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_693), .A2(n_954), .B1(n_955), .B2(n_956), .Y(n_953) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_694), .Y(n_717) );
INVx3_ASAP7_75t_L g1241 ( .A(n_694), .Y(n_1241) );
BUFx6f_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g708 ( .A(n_695), .Y(n_708) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_700), .B(n_863), .Y(n_862) );
AO21x1_ASAP7_75t_L g962 ( .A1(n_701), .A2(n_963), .B(n_967), .Y(n_962) );
OAI33xp33_ASAP7_75t_L g756 ( .A1(n_703), .A2(n_757), .A3(n_760), .B1(n_763), .B2(n_764), .B3(n_767), .Y(n_756) );
OAI33xp33_ASAP7_75t_L g933 ( .A1(n_703), .A2(n_767), .A3(n_934), .B1(n_935), .B2(n_936), .B3(n_938), .Y(n_933) );
OAI33xp33_ASAP7_75t_L g1032 ( .A1(n_703), .A2(n_767), .A3(n_1033), .B1(n_1035), .B2(n_1036), .B3(n_1037), .Y(n_1032) );
OAI33xp33_ASAP7_75t_L g1225 ( .A1(n_703), .A2(n_767), .A3(n_1226), .B1(n_1228), .B2(n_1229), .B3(n_1230), .Y(n_1225) );
INVx1_ASAP7_75t_L g1364 ( .A(n_705), .Y(n_1364) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g881 ( .A(n_708), .Y(n_881) );
INVx2_ASAP7_75t_SL g990 ( .A(n_708), .Y(n_990) );
INVx1_ASAP7_75t_L g1000 ( .A(n_708), .Y(n_1000) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx3_ASAP7_75t_L g882 ( .A(n_711), .Y(n_882) );
INVx2_ASAP7_75t_L g992 ( .A(n_711), .Y(n_992) );
INVx3_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_715), .A2(n_803), .B1(n_816), .B2(n_826), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_715), .A2(n_770), .B1(n_924), .B2(n_928), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1755 ( .A1(n_715), .A2(n_824), .B1(n_1756), .B2(n_1757), .Y(n_1755) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_721), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1270 ( .A(n_726), .Y(n_1270) );
INVx2_ASAP7_75t_L g948 ( .A(n_728), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_1129), .B2(n_1187), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
XOR2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_958), .Y(n_732) );
XNOR2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_846), .Y(n_733) );
XNOR2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_797), .Y(n_734) );
NAND3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_768), .C(n_782), .Y(n_736) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_738), .B(n_756), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_740), .A2(n_753), .B1(n_758), .B2(n_759), .Y(n_757) );
OAI22xp33_ASAP7_75t_L g920 ( .A1(n_741), .A2(n_889), .B1(n_921), .B2(n_922), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_742), .A2(n_754), .B1(n_761), .B2(n_762), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_744), .A2(n_750), .B1(n_761), .B2(n_762), .Y(n_760) );
OAI22xp5_ASAP7_75t_L g1029 ( .A1(n_746), .A2(n_811), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_746), .A2(n_1065), .B1(n_1066), .B2(n_1067), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_746), .A2(n_927), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
OAI22xp33_ASAP7_75t_SL g1760 ( .A1(n_746), .A2(n_1166), .B1(n_1746), .B2(n_1753), .Y(n_1760) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_747), .A2(n_751), .B1(n_759), .B2(n_765), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g1020 ( .A1(n_749), .A2(n_813), .B1(n_1021), .B2(n_1022), .Y(n_1020) );
INVx2_ASAP7_75t_L g1170 ( .A(n_749), .Y(n_1170) );
OAI22xp33_ASAP7_75t_L g1033 ( .A1(n_758), .A2(n_1024), .B1(n_1027), .B2(n_1034), .Y(n_1033) );
OAI22xp5_ASAP7_75t_L g1037 ( .A1(n_758), .A2(n_759), .B1(n_1022), .B2(n_1031), .Y(n_1037) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_758), .A2(n_821), .B1(n_1059), .B2(n_1069), .Y(n_1072) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_758), .A2(n_759), .B1(n_1063), .B2(n_1067), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_758), .A2(n_821), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
OAI22xp33_ASAP7_75t_L g1226 ( .A1(n_758), .A2(n_1214), .B1(n_1223), .B2(n_1227), .Y(n_1226) );
OAI22xp33_ASAP7_75t_L g1748 ( .A1(n_758), .A2(n_1034), .B1(n_1749), .B2(n_1750), .Y(n_1748) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_759), .A2(n_807), .B1(n_812), .B2(n_820), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g934 ( .A1(n_759), .A2(n_820), .B1(n_921), .B2(n_931), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_759), .A2(n_765), .B1(n_1218), .B2(n_1221), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g823 ( .A1(n_761), .A2(n_805), .B1(n_810), .B2(n_824), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_761), .A2(n_762), .B1(n_1025), .B2(n_1028), .Y(n_1036) );
OAI22xp5_ASAP7_75t_L g1228 ( .A1(n_761), .A2(n_762), .B1(n_1217), .B2(n_1220), .Y(n_1228) );
OAI22xp5_ASAP7_75t_L g1745 ( .A1(n_761), .A2(n_937), .B1(n_1746), .B2(n_1747), .Y(n_1745) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_762), .A2(n_1062), .B1(n_1065), .B2(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI33xp33_ASAP7_75t_L g817 ( .A1(n_767), .A2(n_818), .A3(n_819), .B1(n_823), .B2(n_825), .B3(n_827), .Y(n_817) );
NAND3xp33_ASAP7_75t_SL g950 ( .A(n_771), .B(n_951), .C(n_953), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g1259 ( .A(n_771), .B(n_1260), .C(n_1263), .Y(n_1259) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g972 ( .A(n_772), .Y(n_972) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
BUFx2_ASAP7_75t_L g975 ( .A(n_774), .Y(n_975) );
AOI32xp33_ASAP7_75t_L g785 ( .A1(n_777), .A2(n_786), .A3(n_789), .B1(n_791), .B2(n_792), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g1079 ( .A1(n_778), .A2(n_857), .B1(n_1080), .B2(n_1081), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_778), .A2(n_1334), .B1(n_1335), .B2(n_1336), .Y(n_1333) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
OAI31xp33_ASAP7_75t_SL g782 ( .A1(n_783), .A2(n_784), .A3(n_794), .B(n_796), .Y(n_782) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVxp67_ASAP7_75t_L g843 ( .A(n_791), .Y(n_843) );
INVxp67_ASAP7_75t_L g891 ( .A(n_791), .Y(n_891) );
INVx1_ASAP7_75t_L g982 ( .A(n_791), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g1271 ( .A(n_793), .B(n_1272), .C(n_1274), .Y(n_1271) );
NAND3xp33_ASAP7_75t_L g1777 ( .A(n_793), .B(n_1778), .C(n_1779), .Y(n_1777) );
OAI31xp33_ASAP7_75t_SL g839 ( .A1(n_796), .A2(n_840), .A3(n_841), .B(n_842), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g940 ( .A1(n_796), .A2(n_941), .B(n_947), .Y(n_940) );
OAI31xp33_ASAP7_75t_L g1038 ( .A1(n_796), .A2(n_1039), .A3(n_1040), .B(n_1044), .Y(n_1038) );
OAI31xp33_ASAP7_75t_SL g1085 ( .A1(n_796), .A2(n_1086), .A3(n_1087), .B(n_1093), .Y(n_1085) );
OAI31xp33_ASAP7_75t_SL g1122 ( .A1(n_796), .A2(n_1123), .A3(n_1124), .B(n_1127), .Y(n_1122) );
OAI31xp33_ASAP7_75t_L g1202 ( .A1(n_796), .A2(n_1203), .A3(n_1205), .B(n_1210), .Y(n_1202) );
OAI21xp5_ASAP7_75t_L g1268 ( .A1(n_796), .A2(n_1269), .B(n_1271), .Y(n_1268) );
NAND3xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_828), .C(n_839), .Y(n_798) );
NOR2xp33_ASAP7_75t_SL g799 ( .A(n_800), .B(n_817), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_802), .A2(n_815), .B1(n_820), .B2(n_821), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_806), .A2(n_808), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1112 ( .A1(n_806), .A2(n_808), .B1(n_1102), .B2(n_1108), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_806), .A2(n_1172), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_809) );
BUFx6f_ASAP7_75t_L g1312 ( .A(n_818), .Y(n_1312) );
OAI33xp33_ASAP7_75t_L g1359 ( .A1(n_818), .A2(n_1360), .A3(n_1361), .B1(n_1362), .B2(n_1365), .B3(n_1368), .Y(n_1359) );
OAI22xp5_ASAP7_75t_L g1752 ( .A1(n_820), .A2(n_821), .B1(n_1753), .B2(n_1754), .Y(n_1752) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_821), .A2(n_925), .B1(n_929), .B2(n_939), .Y(n_938) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g956 ( .A(n_830), .Y(n_956) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_835), .A2(n_857), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1451 ( .A1(n_835), .A2(n_1334), .B1(n_1452), .B2(n_1453), .Y(n_1451) );
XOR2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_916), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_883), .B(n_885), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_854), .B(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_869), .B(n_872), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g910 ( .A1(n_867), .A2(n_873), .B1(n_911), .B2(n_912), .C(n_913), .Y(n_910) );
OAI22xp5_ASAP7_75t_L g1493 ( .A1(n_868), .A2(n_1494), .B1(n_1496), .B2(n_1497), .Y(n_1493) );
OAI211xp5_ASAP7_75t_SL g872 ( .A1(n_873), .A2(n_874), .B(n_875), .C(n_880), .Y(n_872) );
BUFx6f_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g995 ( .A(n_877), .Y(n_995) );
INVx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
BUFx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_895), .B(n_896), .Y(n_885) );
NAND2xp5_ASAP7_75t_SL g886 ( .A(n_887), .B(n_893), .Y(n_886) );
BUFx2_ASAP7_75t_L g1144 ( .A(n_895), .Y(n_1144) );
OAI31xp33_ASAP7_75t_L g1301 ( .A1(n_895), .A2(n_1302), .A3(n_1303), .B(n_1307), .Y(n_1301) );
OAI31xp33_ASAP7_75t_L g1369 ( .A1(n_895), .A2(n_1370), .A3(n_1371), .B(n_1374), .Y(n_1369) );
OAI211xp5_ASAP7_75t_L g897 ( .A1(n_898), .A2(n_899), .B(n_901), .C(n_906), .Y(n_897) );
OAI221xp5_ASAP7_75t_L g1288 ( .A1(n_899), .A2(n_1172), .B1(n_1289), .B2(n_1290), .C(n_1291), .Y(n_1288) );
OAI22xp33_ASAP7_75t_L g1501 ( .A1(n_899), .A2(n_912), .B1(n_1488), .B2(n_1496), .Y(n_1501) );
INVx2_ASAP7_75t_SL g899 ( .A(n_900), .Y(n_899) );
BUFx3_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx8_ASAP7_75t_L g915 ( .A(n_903), .Y(n_915) );
BUFx3_ASAP7_75t_L g1252 ( .A(n_903), .Y(n_1252) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx12f_ASAP7_75t_L g1004 ( .A(n_908), .Y(n_1004) );
BUFx3_ASAP7_75t_L g1248 ( .A(n_908), .Y(n_1248) );
OAI22xp5_ASAP7_75t_L g1163 ( .A1(n_912), .A2(n_1164), .B1(n_1165), .B2(n_1167), .Y(n_1163) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx8_ASAP7_75t_L g1006 ( .A(n_915), .Y(n_1006) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_940), .C(n_949), .Y(n_917) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_919), .B(n_933), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1761 ( .A1(n_927), .A2(n_1747), .B1(n_1754), .B2(n_1762), .Y(n_1761) );
OAI22xp5_ASAP7_75t_L g1104 ( .A1(n_937), .A2(n_1074), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
HB1xp67_ASAP7_75t_L g1196 ( .A(n_937), .Y(n_1196) );
AOI22xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_1051), .B1(n_1052), .B2(n_1128), .Y(n_958) );
INVx1_ASAP7_75t_L g1128 ( .A(n_959), .Y(n_1128) );
XNOR2x1_ASAP7_75t_SL g959 ( .A(n_960), .B(n_1016), .Y(n_959) );
NAND4xp75_ASAP7_75t_L g961 ( .A(n_962), .B(n_978), .C(n_987), .D(n_1001), .Y(n_961) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_968), .B(n_977), .Y(n_967) );
NAND3xp33_ASAP7_75t_L g968 ( .A(n_969), .B(n_972), .C(n_973), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_976), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx2_ASAP7_75t_L g996 ( .A(n_975), .Y(n_996) );
INVx1_ASAP7_75t_L g998 ( .A(n_975), .Y(n_998) );
AO21x1_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_980), .B(n_985), .Y(n_978) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
OAI31xp33_ASAP7_75t_L g1775 ( .A1(n_986), .A2(n_1776), .A3(n_1777), .B(n_1780), .Y(n_1775) );
NAND3xp33_ASAP7_75t_L g1234 ( .A(n_988), .B(n_1235), .C(n_1239), .Y(n_1234) );
INVx1_ASAP7_75t_L g1751 ( .A(n_988), .Y(n_1751) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
AOI32xp33_ASAP7_75t_L g1001 ( .A1(n_1002), .A2(n_1005), .A3(n_1009), .B1(n_1010), .B2(n_1012), .Y(n_1001) );
BUFx2_ASAP7_75t_L g1292 ( .A(n_1006), .Y(n_1292) );
INVx2_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1008), .Y(n_1253) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1011), .Y(n_1066) );
INVx2_ASAP7_75t_L g1283 ( .A(n_1011), .Y(n_1283) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NAND3xp33_ASAP7_75t_L g1245 ( .A(n_1014), .B(n_1246), .C(n_1249), .Y(n_1245) );
AND3x1_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1038), .C(n_1045), .Y(n_1017) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1032), .Y(n_1018) );
BUFx3_ASAP7_75t_L g1367 ( .A(n_1034), .Y(n_1367) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
XNOR2x1_ASAP7_75t_L g1052 ( .A(n_1053), .B(n_1094), .Y(n_1052) );
XNOR2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1055), .Y(n_1053) );
AND3x1_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1077), .C(n_1085), .Y(n_1055) );
NOR2xp33_ASAP7_75t_SL g1056 ( .A(n_1057), .B(n_1071), .Y(n_1056) );
INVx2_ASAP7_75t_SL g1154 ( .A(n_1083), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1338 ( .A(n_1083), .Y(n_1338) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1090), .Y(n_1446) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1090), .Y(n_1461) );
AND3x1_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1115), .C(n_1122), .Y(n_1095) );
NOR2xp33_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1110), .Y(n_1096) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1187 ( .A(n_1130), .Y(n_1187) );
NAND3xp33_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1145), .C(n_1157), .Y(n_1131) );
OAI31xp33_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1136), .A3(n_1143), .B(n_1144), .Y(n_1132) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1140), .B1(n_1141), .B2(n_1142), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1462 ( .A1(n_1138), .A2(n_1141), .B1(n_1452), .B2(n_1463), .Y(n_1462) );
BUFx3_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
BUFx3_ASAP7_75t_L g1273 ( .A(n_1139), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_1141), .A2(n_1273), .B1(n_1298), .B2(n_1306), .Y(n_1305) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_1141), .A2(n_1273), .B1(n_1335), .B2(n_1373), .Y(n_1372) );
OAI31xp33_ASAP7_75t_L g1456 ( .A1(n_1144), .A2(n_1457), .A3(n_1459), .B(n_1464), .Y(n_1456) );
OAI31xp33_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1152), .A3(n_1155), .B(n_1156), .Y(n_1145) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
OAI31xp33_ASAP7_75t_L g1328 ( .A1(n_1156), .A2(n_1329), .A3(n_1330), .B(n_1337), .Y(n_1328) );
OAI31xp33_ASAP7_75t_L g1447 ( .A1(n_1156), .A2(n_1448), .A3(n_1454), .B(n_1455), .Y(n_1447) );
NOR2xp33_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1177), .Y(n_1157) );
BUFx3_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx8_ASAP7_75t_L g1353 ( .A(n_1166), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1171), .B1(n_1172), .B2(n_1173), .Y(n_1168) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
OAI221xp5_ASAP7_75t_L g1282 ( .A1(n_1172), .A2(n_1283), .B1(n_1284), .B2(n_1285), .C(n_1286), .Y(n_1282) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_1172), .A2(n_1351), .B1(n_1352), .B2(n_1354), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1399 ( .A1(n_1172), .A2(n_1283), .B1(n_1387), .B2(n_1394), .Y(n_1399) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_1172), .A2(n_1429), .B1(n_1435), .B2(n_1441), .Y(n_1440) );
OAI22xp5_ASAP7_75t_L g1442 ( .A1(n_1172), .A2(n_1430), .B1(n_1436), .B2(n_1443), .Y(n_1442) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_1172), .A2(n_1283), .B1(n_1489), .B2(n_1497), .Y(n_1502) );
OAI22xp33_ASAP7_75t_L g1360 ( .A1(n_1180), .A2(n_1227), .B1(n_1342), .B2(n_1357), .Y(n_1360) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx2_ASAP7_75t_SL g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1188), .Y(n_1506) );
XNOR2xp5_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1375), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_1190), .A2(n_1191), .B1(n_1275), .B2(n_1276), .Y(n_1189) );
INVx2_ASAP7_75t_SL g1190 ( .A(n_1191), .Y(n_1190) );
XNOR2x1_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1231), .Y(n_1191) );
NAND3xp33_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1202), .C(n_1211), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1208 ( .A(n_1199), .B(n_1209), .Y(n_1208) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1225), .Y(n_1211) );
NAND3xp33_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1258), .C(n_1268), .Y(n_1232) );
AND4x1_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1242), .C(n_1245), .D(n_1254), .Y(n_1233) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
BUFx2_ASAP7_75t_L g1287 ( .A(n_1252), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1254 ( .A(n_1255), .B(n_1256), .C(n_1257), .Y(n_1254) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
BUFx2_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
XNOR2x1_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1326), .Y(n_1277) );
NAND4xp75_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1294), .C(n_1301), .D(n_1311), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_1284), .A2(n_1289), .B1(n_1317), .B2(n_1320), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1779 ( .A(n_1293), .B(n_1770), .Y(n_1779) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
OAI33xp33_ASAP7_75t_L g1424 ( .A1(n_1312), .A2(n_1368), .A3(n_1425), .B1(n_1428), .B2(n_1431), .B3(n_1434), .Y(n_1424) );
INVx2_ASAP7_75t_L g1317 ( .A(n_1318), .Y(n_1317) );
INVx2_ASAP7_75t_L g1388 ( .A(n_1318), .Y(n_1388) );
INVx4_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1431 ( .A1(n_1320), .A2(n_1363), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
OAI22xp5_ASAP7_75t_L g1393 ( .A1(n_1325), .A2(n_1394), .B1(n_1395), .B2(n_1396), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1434 ( .A1(n_1325), .A2(n_1367), .B1(n_1435), .B2(n_1436), .Y(n_1434) );
AND3x1_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1339), .C(n_1369), .Y(n_1327) );
NOR2xp33_ASAP7_75t_SL g1339 ( .A(n_1340), .B(n_1359), .Y(n_1339) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1343), .B1(n_1345), .B2(n_1346), .Y(n_1341) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g1365 ( .A1(n_1349), .A2(n_1354), .B1(n_1366), .B2(n_1367), .Y(n_1365) );
INVx2_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
XNOR2xp5_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1418), .Y(n_1375) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
NAND3xp33_ASAP7_75t_L g1380 ( .A(n_1381), .B(n_1402), .C(n_1410), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1397), .Y(n_1381) );
INVx2_ASAP7_75t_SL g1418 ( .A(n_1419), .Y(n_1418) );
OA22x2_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1421), .B1(n_1465), .B2(n_1466), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1421), .Y(n_1420) );
NAND3xp33_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1447), .C(n_1456), .Y(n_1422) );
NOR2xp33_ASAP7_75t_SL g1423 ( .A(n_1424), .B(n_1437), .Y(n_1423) );
INVxp67_ASAP7_75t_SL g1445 ( .A(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVxp67_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1461), .Y(n_1500) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1467), .Y(n_1504) );
NAND3xp33_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1476), .C(n_1482), .Y(n_1467) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1498), .Y(n_1482) );
INVx2_ASAP7_75t_L g1494 ( .A(n_1495), .Y(n_1494) );
OAI221xp5_ASAP7_75t_SL g1507 ( .A1(n_1508), .A2(n_1737), .B1(n_1740), .B2(n_1783), .C(n_1786), .Y(n_1507) );
AOI21xp5_ASAP7_75t_L g1508 ( .A1(n_1509), .A2(n_1651), .B(n_1704), .Y(n_1508) );
NAND4xp25_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1621), .C(n_1637), .D(n_1643), .Y(n_1509) );
NOR5xp2_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1575), .C(n_1588), .D(n_1595), .E(n_1618), .Y(n_1510) );
OAI21xp5_ASAP7_75t_SL g1511 ( .A1(n_1512), .A2(n_1532), .B(n_1551), .Y(n_1511) );
NOR2xp33_ASAP7_75t_L g1552 ( .A(n_1512), .B(n_1533), .Y(n_1552) );
OAI31xp33_ASAP7_75t_L g1729 ( .A1(n_1512), .A2(n_1730), .A3(n_1731), .B(n_1732), .Y(n_1729) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
AND2x2_ASAP7_75t_L g1650 ( .A(n_1513), .B(n_1608), .Y(n_1650) );
AOI221xp5_ASAP7_75t_L g1667 ( .A1(n_1513), .A2(n_1591), .B1(n_1668), .B2(n_1669), .C(n_1671), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1514), .B(n_1528), .Y(n_1513) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1514), .Y(n_1578) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1514), .Y(n_1590) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1514), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1640 ( .A(n_1514), .B(n_1566), .Y(n_1640) );
NAND2xp5_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1522), .Y(n_1514) );
AND2x6_ASAP7_75t_L g1516 ( .A(n_1517), .B(n_1518), .Y(n_1516) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1517), .B(n_1521), .Y(n_1520) );
AND2x4_ASAP7_75t_L g1523 ( .A(n_1517), .B(n_1524), .Y(n_1523) );
AND2x6_ASAP7_75t_L g1526 ( .A(n_1517), .B(n_1527), .Y(n_1526) );
AND2x2_ASAP7_75t_L g1530 ( .A(n_1517), .B(n_1521), .Y(n_1530) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1517), .B(n_1521), .Y(n_1612) );
NAND2xp5_ASAP7_75t_L g1739 ( .A(n_1517), .B(n_1524), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1519), .B(n_1525), .Y(n_1524) );
HB1xp67_ASAP7_75t_L g1797 ( .A(n_1524), .Y(n_1797) );
CKINVDCx5p33_ASAP7_75t_R g1566 ( .A(n_1528), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1587 ( .A(n_1528), .B(n_1563), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1615 ( .A(n_1528), .B(n_1578), .Y(n_1615) );
HB1xp67_ASAP7_75t_SL g1633 ( .A(n_1528), .Y(n_1633) );
NAND2xp5_ASAP7_75t_L g1697 ( .A(n_1528), .B(n_1608), .Y(n_1697) );
NAND2xp5_ASAP7_75t_L g1709 ( .A(n_1528), .B(n_1535), .Y(n_1709) );
AND2x4_ASAP7_75t_L g1528 ( .A(n_1529), .B(n_1531), .Y(n_1528) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1532), .Y(n_1720) );
NAND2xp5_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1538), .Y(n_1532) );
AND2x2_ASAP7_75t_L g1644 ( .A(n_1533), .B(n_1570), .Y(n_1644) );
NAND2xp5_ASAP7_75t_L g1727 ( .A(n_1533), .B(n_1616), .Y(n_1727) );
CKINVDCx14_ASAP7_75t_R g1533 ( .A(n_1534), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1534), .B(n_1586), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1593 ( .A(n_1534), .B(n_1563), .Y(n_1593) );
NAND2xp5_ASAP7_75t_L g1601 ( .A(n_1534), .B(n_1555), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1647 ( .A(n_1534), .B(n_1583), .Y(n_1647) );
AND2x2_ASAP7_75t_L g1661 ( .A(n_1534), .B(n_1662), .Y(n_1661) );
NOR2xp33_ASAP7_75t_L g1673 ( .A(n_1534), .B(n_1587), .Y(n_1673) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1534), .B(n_1629), .Y(n_1693) );
NOR2xp33_ASAP7_75t_L g1703 ( .A(n_1534), .B(n_1596), .Y(n_1703) );
INVx3_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
CKINVDCx5p33_ASAP7_75t_R g1567 ( .A(n_1535), .Y(n_1567) );
NOR2xp33_ASAP7_75t_L g1604 ( .A(n_1535), .B(n_1572), .Y(n_1604) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1535), .B(n_1540), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1642 ( .A(n_1535), .B(n_1556), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1677 ( .A(n_1535), .B(n_1649), .Y(n_1677) );
NAND2xp5_ASAP7_75t_L g1699 ( .A(n_1535), .B(n_1658), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1535), .B(n_1583), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1731 ( .A(n_1535), .B(n_1629), .Y(n_1731) );
AND2x4_ASAP7_75t_SL g1535 ( .A(n_1536), .B(n_1537), .Y(n_1535) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
OR2x2_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1543), .Y(n_1539) );
INVx2_ASAP7_75t_L g1555 ( .A(n_1540), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1540), .B(n_1548), .Y(n_1558) );
AND2x2_ASAP7_75t_L g1574 ( .A(n_1540), .B(n_1557), .Y(n_1574) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1540), .B(n_1556), .Y(n_1632) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1540), .B(n_1656), .Y(n_1655) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1540), .B(n_1545), .Y(n_1670) );
OAI322xp33_ASAP7_75t_L g1671 ( .A1(n_1540), .A2(n_1554), .A3(n_1649), .B1(n_1672), .B2(n_1674), .C1(n_1678), .C2(n_1680), .Y(n_1671) );
OR2x2_ASAP7_75t_L g1707 ( .A(n_1540), .B(n_1642), .Y(n_1707) );
OR2x2_ASAP7_75t_L g1718 ( .A(n_1540), .B(n_1545), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1542), .Y(n_1540) );
OR2x2_ASAP7_75t_L g1617 ( .A(n_1543), .B(n_1555), .Y(n_1617) );
INVx1_ASAP7_75t_L g1658 ( .A(n_1543), .Y(n_1658) );
OR2x2_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1548), .Y(n_1543) );
AND2x2_ASAP7_75t_L g1556 ( .A(n_1544), .B(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1572 ( .A(n_1545), .B(n_1573), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1545), .B(n_1548), .Y(n_1583) );
AND2x2_ASAP7_75t_L g1635 ( .A(n_1545), .B(n_1555), .Y(n_1635) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1547), .Y(n_1545) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1548), .Y(n_1557) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1548), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1690 ( .A(n_1548), .B(n_1555), .Y(n_1690) );
NAND2x1_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1550), .Y(n_1548) );
AOI22xp33_ASAP7_75t_L g1551 ( .A1(n_1552), .A2(n_1553), .B1(n_1559), .B2(n_1568), .Y(n_1551) );
NAND2xp5_ASAP7_75t_L g1553 ( .A(n_1554), .B(n_1558), .Y(n_1553) );
NAND2xp5_ASAP7_75t_L g1554 ( .A(n_1555), .B(n_1556), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1570 ( .A(n_1555), .B(n_1571), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1582 ( .A(n_1555), .B(n_1583), .Y(n_1582) );
OR2x2_ASAP7_75t_L g1627 ( .A(n_1555), .B(n_1628), .Y(n_1627) );
OR2x2_ASAP7_75t_L g1663 ( .A(n_1555), .B(n_1572), .Y(n_1663) );
NOR2xp33_ASAP7_75t_L g1675 ( .A(n_1555), .B(n_1676), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1556), .B(n_1600), .Y(n_1599) );
NAND2xp5_ASAP7_75t_L g1606 ( .A(n_1556), .B(n_1607), .Y(n_1606) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_1556), .B(n_1567), .Y(n_1656) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1558), .Y(n_1620) );
OAI21xp5_ASAP7_75t_L g1708 ( .A1(n_1558), .A2(n_1709), .B(n_1710), .Y(n_1708) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
NAND2xp5_ASAP7_75t_L g1560 ( .A(n_1561), .B(n_1567), .Y(n_1560) );
INVx1_ASAP7_75t_L g1736 ( .A(n_1561), .Y(n_1736) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1562), .Y(n_1561) );
OR2x2_ASAP7_75t_L g1576 ( .A(n_1562), .B(n_1577), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1563), .B(n_1566), .Y(n_1562) );
INVx2_ASAP7_75t_SL g1597 ( .A(n_1563), .Y(n_1597) );
INVx1_ASAP7_75t_L g1608 ( .A(n_1563), .Y(n_1608) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1565), .Y(n_1563) );
OR2x2_ASAP7_75t_L g1596 ( .A(n_1566), .B(n_1597), .Y(n_1596) );
AND2x2_ASAP7_75t_L g1603 ( .A(n_1566), .B(n_1590), .Y(n_1603) );
NOR2xp33_ASAP7_75t_L g1622 ( .A(n_1566), .B(n_1623), .Y(n_1622) );
OAI22xp5_ASAP7_75t_L g1653 ( .A1(n_1566), .A2(n_1633), .B1(n_1654), .B2(n_1657), .Y(n_1653) );
NAND3xp33_ASAP7_75t_L g1692 ( .A(n_1566), .B(n_1583), .C(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1567), .Y(n_1581) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_1567), .B(n_1689), .Y(n_1688) );
INVxp33_ASAP7_75t_SL g1568 ( .A(n_1569), .Y(n_1568) );
NOR2xp33_ASAP7_75t_SL g1569 ( .A(n_1570), .B(n_1574), .Y(n_1569) );
INVx2_ASAP7_75t_L g1594 ( .A(n_1570), .Y(n_1594) );
AOI222xp33_ASAP7_75t_L g1643 ( .A1(n_1571), .A2(n_1644), .B1(n_1645), .B2(n_1646), .C1(n_1648), .C2(n_1650), .Y(n_1643) );
NOR2xp33_ASAP7_75t_L g1679 ( .A(n_1571), .B(n_1658), .Y(n_1679) );
A2O1A1Ixp33_ASAP7_75t_L g1732 ( .A1(n_1571), .A2(n_1581), .B(n_1650), .C(n_1662), .Y(n_1732) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1572), .Y(n_1571) );
A2O1A1Ixp33_ASAP7_75t_L g1733 ( .A1(n_1574), .A2(n_1645), .B(n_1673), .C(n_1734), .Y(n_1733) );
OAI21xp5_ASAP7_75t_SL g1575 ( .A1(n_1576), .A2(n_1579), .B(n_1584), .Y(n_1575) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1576), .Y(n_1728) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1578), .Y(n_1649) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1578), .B(n_1625), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1668 ( .A(n_1578), .B(n_1586), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1578), .B(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
AND2x2_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1582), .Y(n_1580) );
AOI221xp5_ASAP7_75t_L g1719 ( .A1(n_1582), .A2(n_1685), .B1(n_1720), .B2(n_1721), .C(n_1722), .Y(n_1719) );
NAND2xp5_ASAP7_75t_L g1584 ( .A(n_1583), .B(n_1585), .Y(n_1584) );
INVx1_ASAP7_75t_L g1628 ( .A(n_1583), .Y(n_1628) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1583), .B(n_1607), .Y(n_1712) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1585), .B(n_1620), .Y(n_1619) );
NAND2xp5_ASAP7_75t_L g1634 ( .A(n_1585), .B(n_1635), .Y(n_1634) );
NAND2xp5_ASAP7_75t_L g1686 ( .A(n_1586), .B(n_1645), .Y(n_1686) );
INVx2_ASAP7_75t_L g1586 ( .A(n_1587), .Y(n_1586) );
AOI21xp33_ASAP7_75t_L g1652 ( .A1(n_1587), .A2(n_1653), .B(n_1659), .Y(n_1652) );
INVxp67_ASAP7_75t_SL g1588 ( .A(n_1589), .Y(n_1588) );
NAND2xp5_ASAP7_75t_L g1589 ( .A(n_1590), .B(n_1591), .Y(n_1589) );
NOR2xp33_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1594), .Y(n_1591) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
OAI21xp33_ASAP7_75t_L g1614 ( .A1(n_1593), .A2(n_1615), .B(n_1616), .Y(n_1614) );
OAI211xp5_ASAP7_75t_SL g1595 ( .A1(n_1596), .A2(n_1598), .B(n_1602), .C(n_1614), .Y(n_1595) );
INVx1_ASAP7_75t_L g1721 ( .A(n_1596), .Y(n_1721) );
INVx2_ASAP7_75t_L g1629 ( .A(n_1597), .Y(n_1629) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1597), .B(n_1712), .Y(n_1711) );
O2A1O1Ixp33_ASAP7_75t_SL g1722 ( .A1(n_1597), .A2(n_1664), .B(n_1723), .C(n_1724), .Y(n_1722) );
CKINVDCx14_ASAP7_75t_R g1598 ( .A(n_1599), .Y(n_1598) );
NAND2xp5_ASAP7_75t_L g1657 ( .A(n_1600), .B(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
OR2x2_ASAP7_75t_L g1664 ( .A(n_1601), .B(n_1628), .Y(n_1664) );
AOI211xp5_ASAP7_75t_L g1713 ( .A1(n_1601), .A2(n_1714), .B(n_1715), .C(n_1717), .Y(n_1713) );
AOI221xp5_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1604), .B1(n_1605), .B2(n_1608), .C(n_1609), .Y(n_1602) );
NOR2xp33_ASAP7_75t_L g1626 ( .A(n_1603), .B(n_1627), .Y(n_1626) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1603), .Y(n_1680) );
O2A1O1Ixp33_ASAP7_75t_L g1725 ( .A1(n_1604), .A2(n_1726), .B(n_1728), .C(n_1729), .Y(n_1725) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
NAND2xp5_ASAP7_75t_L g1624 ( .A(n_1606), .B(n_1625), .Y(n_1624) );
INVx2_ASAP7_75t_L g1625 ( .A(n_1608), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_1609), .B(n_1692), .Y(n_1691) );
INVx3_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
AND2x2_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1613), .Y(n_1610) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1615), .Y(n_1724) );
INVx2_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
INVxp67_ASAP7_75t_SL g1618 ( .A(n_1619), .Y(n_1618) );
O2A1O1Ixp33_ASAP7_75t_L g1621 ( .A1(n_1622), .A2(n_1626), .B(n_1629), .C(n_1630), .Y(n_1621) );
OAI31xp33_ASAP7_75t_L g1637 ( .A1(n_1622), .A2(n_1626), .A3(n_1638), .B(n_1641), .Y(n_1637) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
AND2x2_ASAP7_75t_L g1648 ( .A(n_1625), .B(n_1649), .Y(n_1648) );
OR2x2_ASAP7_75t_L g1684 ( .A(n_1625), .B(n_1649), .Y(n_1684) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1627), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1639 ( .A(n_1629), .B(n_1640), .Y(n_1639) );
O2A1O1Ixp33_ASAP7_75t_L g1630 ( .A1(n_1631), .A2(n_1633), .B(n_1634), .C(n_1636), .Y(n_1630) );
AOI21xp33_ASAP7_75t_L g1734 ( .A1(n_1631), .A2(n_1735), .B(n_1736), .Y(n_1734) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
NAND2xp5_ASAP7_75t_L g1702 ( .A(n_1635), .B(n_1703), .Y(n_1702) );
CKINVDCx14_ASAP7_75t_R g1730 ( .A(n_1635), .Y(n_1730) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1636), .Y(n_1645) );
AOI221xp5_ASAP7_75t_L g1705 ( .A1(n_1636), .A2(n_1668), .B1(n_1706), .B2(n_1708), .C(n_1713), .Y(n_1705) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1641), .Y(n_1723) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1644), .Y(n_1735) );
INVx1_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
AOI222xp33_ASAP7_75t_L g1694 ( .A1(n_1648), .A2(n_1683), .B1(n_1695), .B2(n_1696), .C1(n_1698), .C2(n_1700), .Y(n_1694) );
NAND5xp2_ASAP7_75t_L g1651 ( .A(n_1652), .B(n_1667), .C(n_1681), .D(n_1694), .E(n_1702), .Y(n_1651) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVxp67_ASAP7_75t_SL g1714 ( .A(n_1656), .Y(n_1714) );
AOI21xp33_ASAP7_75t_L g1659 ( .A1(n_1660), .A2(n_1664), .B(n_1665), .Y(n_1659) );
INVx1_ASAP7_75t_L g1660 ( .A(n_1661), .Y(n_1660) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1664), .Y(n_1695) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVxp67_ASAP7_75t_SL g1672 ( .A(n_1673), .Y(n_1672) );
INVxp67_ASAP7_75t_L g1674 ( .A(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
HB1xp67_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
AOI221xp5_ASAP7_75t_L g1681 ( .A1(n_1682), .A2(n_1683), .B1(n_1685), .B2(n_1687), .C(n_1691), .Y(n_1681) );
INVx1_ASAP7_75t_L g1683 ( .A(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx1_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
INVx1_ASAP7_75t_L g1716 ( .A(n_1697), .Y(n_1716) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1699), .Y(n_1698) );
INVxp67_ASAP7_75t_SL g1700 ( .A(n_1701), .Y(n_1700) );
NAND4xp25_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1719), .C(n_1725), .D(n_1733), .Y(n_1704) );
INVxp67_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
INVx1_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1717 ( .A(n_1718), .Y(n_1717) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
CKINVDCx20_ASAP7_75t_R g1737 ( .A(n_1738), .Y(n_1737) );
CKINVDCx5p33_ASAP7_75t_R g1738 ( .A(n_1739), .Y(n_1738) );
INVx3_ASAP7_75t_SL g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1742), .Y(n_1782) );
NAND3xp33_ASAP7_75t_L g1742 ( .A(n_1743), .B(n_1765), .C(n_1775), .Y(n_1742) );
NOR2xp33_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1758), .Y(n_1743) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
HB1xp67_ASAP7_75t_L g1792 ( .A(n_1782), .Y(n_1792) );
CKINVDCx5p33_ASAP7_75t_R g1783 ( .A(n_1784), .Y(n_1783) );
HB1xp67_ASAP7_75t_SL g1787 ( .A(n_1788), .Y(n_1787) );
BUFx3_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
INVxp33_ASAP7_75t_SL g1790 ( .A(n_1791), .Y(n_1790) );
HB1xp67_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
HB1xp67_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
OAI21xp5_ASAP7_75t_L g1795 ( .A1(n_1796), .A2(n_1797), .B(n_1798), .Y(n_1795) );
INVx1_ASAP7_75t_L g1798 ( .A(n_1799), .Y(n_1798) );
endmodule