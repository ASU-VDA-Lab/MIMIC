module fake_jpeg_5103_n_213 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_213);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_213;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_34),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_25),
.B(n_27),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_49),
.C(n_56),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_31),
.B1(n_29),
.B2(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_58),
.B1(n_60),
.B2(n_24),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_20),
.B1(n_30),
.B2(n_26),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_45),
.A2(n_52),
.B1(n_35),
.B2(n_42),
.Y(n_82)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_31),
.Y(n_49)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_17),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_55)
);

OAI22x1_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_27),
.B1(n_39),
.B2(n_22),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_30),
.B1(n_26),
.B2(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_28),
.B1(n_21),
.B2(n_23),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_28),
.B1(n_21),
.B2(n_23),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_64),
.Y(n_67)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_68),
.Y(n_89)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_71),
.Y(n_87)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_74),
.B(n_1),
.Y(n_106)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_76),
.B(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_82),
.B1(n_56),
.B2(n_15),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_15),
.B1(n_17),
.B2(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_38),
.C(n_32),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_49),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_49),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_98),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_27),
.B(n_46),
.C(n_18),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_69),
.A2(n_84),
.B(n_74),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_102),
.B1(n_46),
.B2(n_57),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_81),
.B(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_15),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_46),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_93),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_114),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_71),
.B1(n_80),
.B2(n_108),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_78),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_38),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_96),
.B1(n_99),
.B2(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_68),
.Y(n_122)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_100),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_103),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_97),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_148),
.C(n_38),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_131),
.A2(n_139),
.B(n_142),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_135),
.A2(n_144),
.B1(n_113),
.B2(n_110),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_86),
.B(n_92),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_143),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_94),
.B(n_102),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_101),
.Y(n_143)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_105),
.B(n_87),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_67),
.B1(n_108),
.B2(n_107),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_52),
.B1(n_59),
.B2(n_118),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_105),
.B(n_107),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_67),
.B(n_38),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_91),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_147),
.B(n_117),
.Y(n_150)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_47),
.C(n_48),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_157),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_154),
.B1(n_160),
.B2(n_145),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_165),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_141),
.A2(n_113),
.B1(n_129),
.B2(n_128),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_38),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_135),
.C(n_142),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_52),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_109),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_172),
.C(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_149),
.C(n_148),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_137),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_175),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_179),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_145),
.B(n_144),
.C(n_143),
.D(n_131),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_176),
.A2(n_144),
.B(n_153),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_165),
.B(n_158),
.C(n_160),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_133),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_177),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_187),
.B1(n_172),
.B2(n_167),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_190),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_156),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_170),
.C(n_173),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_171),
.A2(n_70),
.B(n_18),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_196),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_175),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_198),
.C(n_188),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_186),
.A2(n_88),
.B1(n_14),
.B2(n_13),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_189),
.B(n_119),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_27),
.C(n_14),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_203),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_181),
.C(n_185),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_193),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_207),
.B(n_12),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_180),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_192),
.B1(n_191),
.B2(n_199),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_205),
.A3(n_204),
.B1(n_10),
.B2(n_11),
.C1(n_9),
.C2(n_8),
.Y(n_211)
);

AOI321xp33_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_76),
.C(n_209),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_210),
.Y(n_213)
);


endmodule