module fake_jpeg_24543_n_304 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_156;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_288;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_265;
wire n_115;
wire n_123;
wire n_273;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx11_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_12),
.B(n_5),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_2),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_53),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_26),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_34),
.B1(n_35),
.B2(n_32),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_28),
.B1(n_34),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_55),
.A2(n_84),
.B1(n_24),
.B2(n_19),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_35),
.B1(n_21),
.B2(n_25),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_77),
.B1(n_11),
.B2(n_12),
.Y(n_113)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_23),
.B1(n_25),
.B2(n_21),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_1),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_69),
.B(n_73),
.C(n_85),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_23),
.B1(n_31),
.B2(n_22),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_78),
.B1(n_24),
.B2(n_19),
.Y(n_98)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_80),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_36),
.B(n_29),
.C(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_36),
.B(n_19),
.C(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_36),
.B1(n_33),
.B2(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_43),
.B(n_38),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_49),
.B(n_2),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_3),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_33),
.B1(n_29),
.B2(n_24),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_40),
.B(n_4),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_6),
.Y(n_90)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_105),
.B1(n_110),
.B2(n_115),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_98),
.A2(n_102),
.B1(n_85),
.B2(n_112),
.Y(n_127)
);

NOR4xp25_ASAP7_75t_SL g101 ( 
.A(n_69),
.B(n_17),
.C(n_7),
.D(n_9),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_13),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_18),
.B1(n_36),
.B2(n_10),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_6),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_80),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_73),
.A2(n_36),
.B1(n_10),
.B2(n_11),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_9),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx2_ASAP7_75t_SL g138 ( 
.A(n_107),
.Y(n_138)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

BUFx2_ASAP7_75t_SL g144 ( 
.A(n_108),
.Y(n_144)
);

AND2x6_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_9),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_117),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_86),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_59),
.A2(n_58),
.B1(n_74),
.B2(n_77),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_121),
.B1(n_51),
.B2(n_82),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_74),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_122),
.Y(n_166)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_127),
.A2(n_141),
.B1(n_154),
.B2(n_108),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_67),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_116),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_140),
.Y(n_163)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_50),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_66),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_70),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_87),
.Y(n_146)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_121),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_95),
.A2(n_117),
.B1(n_118),
.B2(n_60),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_151),
.B(n_114),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_14),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_60),
.B1(n_71),
.B2(n_61),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_111),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_94),
.B(n_80),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_153),
.B(n_15),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_99),
.A2(n_77),
.B1(n_84),
.B2(n_55),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_105),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_158),
.B(n_167),
.Y(n_204)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_152),
.A2(n_110),
.B(n_75),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_16),
.B(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_175),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_94),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_170),
.B(n_172),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_130),
.B(n_100),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_100),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_180),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_97),
.B1(n_119),
.B2(n_113),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_174),
.A2(n_186),
.B1(n_139),
.B2(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_93),
.B(n_102),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_178),
.B(n_182),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_181),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_93),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_141),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_103),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_125),
.B(n_123),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_133),
.A2(n_65),
.B(n_103),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_184),
.Y(n_196)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_132),
.B1(n_150),
.B2(n_135),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_77),
.B1(n_76),
.B2(n_109),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_157),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_132),
.B1(n_150),
.B2(n_142),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_189),
.A2(n_191),
.B1(n_213),
.B2(n_178),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_207),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_200),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_206),
.C(n_208),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_166),
.B(n_139),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_202),
.B(n_166),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_125),
.B(n_123),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_205),
.A2(n_210),
.B(n_169),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_134),
.C(n_143),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_158),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_136),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_211),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_16),
.B(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_182),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_174),
.A2(n_126),
.B1(n_109),
.B2(n_16),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_225),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_164),
.B1(n_165),
.B2(n_184),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_221),
.A2(n_234),
.B1(n_235),
.B2(n_210),
.Y(n_244)
);

BUFx12_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_230),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_204),
.C(n_188),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_192),
.Y(n_236)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx2_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_196),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_197),
.B1(n_213),
.B2(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_232),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_237),
.C(n_250),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_212),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_231),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_246),
.Y(n_260)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_249),
.B(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

A2O1A1O1Ixp25_ASAP7_75t_L g250 ( 
.A1(n_235),
.A2(n_207),
.B(n_170),
.C(n_172),
.D(n_163),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_173),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_252),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_180),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_254),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_247),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_255),
.A2(n_258),
.B(n_259),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_215),
.B1(n_228),
.B2(n_214),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_256),
.A2(n_257),
.B1(n_220),
.B2(n_240),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_219),
.B(n_226),
.Y(n_259)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_217),
.CI(n_220),
.CON(n_261),
.SN(n_261)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_261),
.Y(n_272)
);

BUFx12_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_219),
.B(n_222),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_252),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_273),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_236),
.C(n_237),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_278),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_258),
.B1(n_239),
.B2(n_260),
.Y(n_271)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_271),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_248),
.B(n_223),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_275),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_282),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_232),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_229),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_270),
.A2(n_259),
.B(n_265),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_203),
.B(n_261),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_230),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_286),
.A2(n_263),
.B1(n_273),
.B2(n_225),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_281),
.B(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_293),
.B(n_288),
.Y(n_297)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_223),
.B(n_272),
.Y(n_296)
);

OAI32xp33_ASAP7_75t_SL g298 ( 
.A1(n_296),
.A2(n_203),
.A3(n_163),
.B1(n_175),
.B2(n_161),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_297),
.A2(n_298),
.B1(n_295),
.B2(n_161),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_285),
.Y(n_299)
);

OAI221xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_285),
.B1(n_268),
.B2(n_294),
.C(n_269),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_301),
.C(n_298),
.Y(n_302)
);

OAI221xp5_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_223),
.B1(n_156),
.B2(n_181),
.C(n_160),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_304)
);


endmodule