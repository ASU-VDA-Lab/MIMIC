module fake_jpeg_26410_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_26),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_43),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_54),
.Y(n_68)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_53),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_28),
.B1(n_22),
.B2(n_16),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_38),
.Y(n_66)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_28),
.B1(n_22),
.B2(n_25),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_22),
.B1(n_19),
.B2(n_30),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_62),
.A2(n_70),
.B1(n_45),
.B2(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_69),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_42),
.B1(n_36),
.B2(n_39),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_42),
.C(n_36),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_90),
.C(n_46),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_44),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_35),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_29),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_43),
.B1(n_22),
.B2(n_16),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_52),
.B1(n_19),
.B2(n_32),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_20),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_17),
.B1(n_25),
.B2(n_30),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_31),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_92),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_89),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_17),
.B1(n_25),
.B2(n_30),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_19),
.B1(n_23),
.B2(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_50),
.B(n_17),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_47),
.B(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_46),
.B(n_23),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_93),
.A2(n_101),
.B(n_109),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_98),
.B1(n_100),
.B2(n_103),
.Y(n_122)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_75),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_69),
.A2(n_56),
.B1(n_53),
.B2(n_58),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_26),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_53),
.B1(n_58),
.B2(n_52),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_88),
.B1(n_78),
.B2(n_87),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_80),
.Y(n_109)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_91),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_117),
.A2(n_85),
.B1(n_92),
.B2(n_90),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_46),
.C(n_60),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_118),
.B(n_60),
.C(n_75),
.Y(n_134)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_87),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_89),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_0),
.B(n_1),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_32),
.B(n_18),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_121),
.A2(n_64),
.B(n_63),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_108),
.B(n_120),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_142),
.B1(n_97),
.B2(n_110),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_98),
.A2(n_72),
.B1(n_74),
.B2(n_83),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_125),
.A2(n_141),
.B1(n_151),
.B2(n_110),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_95),
.A2(n_67),
.B1(n_78),
.B2(n_66),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_128),
.A2(n_133),
.B1(n_147),
.B2(n_106),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_65),
.Y(n_130)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_65),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_131),
.B(n_111),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_132),
.B(n_134),
.C(n_146),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_136),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_118),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_137),
.A2(n_144),
.B(n_101),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_139),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_104),
.A2(n_33),
.B1(n_32),
.B2(n_18),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_33),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_149),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_32),
.B1(n_18),
.B2(n_21),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_108),
.B(n_99),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_60),
.C(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_27),
.B1(n_24),
.B2(n_32),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_101),
.A2(n_103),
.B1(n_109),
.B2(n_100),
.Y(n_151)
);

AO22x1_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_109),
.B1(n_93),
.B2(n_107),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_141),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_155),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_147),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_112),
.B1(n_96),
.B2(n_116),
.Y(n_160)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_160),
.A2(n_14),
.B1(n_15),
.B2(n_155),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_162),
.B1(n_175),
.B2(n_181),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_150),
.A2(n_97),
.B(n_102),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_165),
.A2(n_168),
.B(n_171),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_117),
.B1(n_106),
.B2(n_96),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_169),
.B1(n_170),
.B2(n_9),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_178),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_150),
.A2(n_114),
.B(n_32),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_112),
.B1(n_115),
.B2(n_27),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_21),
.B1(n_18),
.B2(n_60),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_128),
.A2(n_21),
.B(n_18),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_21),
.B(n_1),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_174),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_122),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_136),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_126),
.B(n_132),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_151),
.A2(n_0),
.B(n_2),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_129),
.B1(n_125),
.B2(n_144),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_185),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_130),
.A2(n_2),
.B(n_3),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_124),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_3),
.B(n_8),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_131),
.A2(n_8),
.B(n_9),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_188),
.A2(n_207),
.B(n_171),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_138),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_192),
.B(n_193),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_195),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_167),
.B(n_138),
.C(n_140),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_198),
.C(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_199),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_140),
.C(n_148),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_182),
.B1(n_175),
.B2(n_181),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_202),
.A2(n_212),
.B1(n_179),
.B2(n_185),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_11),
.C(n_13),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_160),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_14),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_183),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_14),
.B1(n_15),
.B2(n_161),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_153),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_15),
.Y(n_215)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_215),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_225),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_187),
.B1(n_212),
.B2(n_211),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_177),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_232),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_178),
.B(n_168),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_235),
.B(n_186),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_203),
.B(n_163),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_152),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_156),
.B(n_174),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_166),
.C(n_154),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_187),
.C(n_154),
.Y(n_250)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_235),
.B(n_188),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_241),
.A2(n_251),
.B(n_228),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_242),
.B(n_219),
.Y(n_261)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_203),
.B(n_190),
.C(n_206),
.D(n_200),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_249),
.Y(n_263)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_255),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_259),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_206),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_225),
.B(n_180),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_176),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_158),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_236),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_158),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_223),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_217),
.A2(n_186),
.B1(n_208),
.B2(n_210),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_218),
.B1(n_238),
.B2(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_248),
.B(n_218),
.C(n_237),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_275),
.C(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_227),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_262),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_272),
.Y(n_281)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_276),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_271),
.B1(n_253),
.B2(n_257),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_153),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_222),
.B1(n_239),
.B2(n_220),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_240),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_233),
.C(n_204),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_252),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_256),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_283),
.Y(n_291)
);

NAND2x1_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_252),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_241),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_269),
.C(n_274),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_264),
.C(n_273),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_254),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_295),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_273),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_301),
.C(n_290),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_264),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_246),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_285),
.A2(n_272),
.B1(n_245),
.B2(n_266),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_298),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_262),
.C(n_263),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_262),
.B(n_246),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_302),
.A2(n_292),
.B(n_293),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_304),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_311),
.C(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_288),
.C(n_281),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_310),
.B(n_291),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_301),
.A2(n_281),
.B1(n_276),
.B2(n_243),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_316),
.Y(n_318)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_319),
.C(n_312),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_315),
.A2(n_306),
.B(n_303),
.Y(n_319)
);

O2A1O1Ixp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_318),
.B(n_305),
.C(n_299),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_300),
.C(n_263),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_202),
.B(n_240),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_170),
.Y(n_324)
);


endmodule