module fake_jpeg_12203_n_613 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_613);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_483;
wire n_236;
wire n_291;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_15),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_68),
.Y(n_126)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_63),
.B(n_64),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_14),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_65),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_25),
.B(n_14),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_71),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_75),
.Y(n_167)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_76),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_82),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_18),
.Y(n_84)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_88),
.Y(n_170)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_90),
.Y(n_134)
);

HAxp5_ASAP7_75t_SL g91 ( 
.A(n_40),
.B(n_0),
.CON(n_91),
.SN(n_91)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_91),
.A2(n_0),
.B(n_3),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_14),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_104),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_18),
.Y(n_94)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_96),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_24),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_18),
.Y(n_102)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_103),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_37),
.B(n_12),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_107),
.Y(n_149)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_37),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_121),
.Y(n_178)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_20),
.B(n_11),
.C(n_2),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_113),
.B(n_29),
.C(n_50),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_32),
.Y(n_115)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_116),
.Y(n_197)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_117),
.Y(n_200)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_26),
.Y(n_119)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_39),
.Y(n_122)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_41),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_33),
.Y(n_131)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_84),
.A2(n_55),
.B1(n_57),
.B2(n_48),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_129),
.A2(n_146),
.B1(n_177),
.B2(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_131),
.B(n_160),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_88),
.A2(n_26),
.B1(n_48),
.B2(n_19),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_133),
.A2(n_165),
.B(n_172),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_61),
.A2(n_45),
.B1(n_34),
.B2(n_51),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_153),
.B(n_183),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_94),
.A2(n_45),
.B1(n_34),
.B2(n_51),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_157),
.A2(n_206),
.B1(n_93),
.B2(n_75),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_29),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_88),
.A2(n_48),
.B1(n_32),
.B2(n_51),
.Y(n_165)
);

INVx6_ASAP7_75t_SL g166 ( 
.A(n_71),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_91),
.A2(n_49),
.B(n_48),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_90),
.A2(n_34),
.B1(n_45),
.B2(n_35),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_180),
.B(n_191),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_90),
.A2(n_27),
.B1(n_35),
.B2(n_38),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_82),
.B(n_46),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_99),
.A2(n_38),
.B1(n_27),
.B2(n_46),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_188),
.B1(n_195),
.B2(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_87),
.B(n_50),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_187),
.B(n_89),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_102),
.A2(n_49),
.B1(n_33),
.B2(n_52),
.Y(n_188)
);

AND2x4_ASAP7_75t_L g191 ( 
.A(n_118),
.B(n_54),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_96),
.B(n_108),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_192),
.B(n_3),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_110),
.A2(n_52),
.B1(n_54),
.B2(n_23),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_199),
.B(n_3),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_115),
.A2(n_52),
.B1(n_28),
.B2(n_54),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_77),
.A2(n_79),
.B1(n_112),
.B2(n_103),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_80),
.B1(n_83),
.B2(n_85),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_207),
.A2(n_249),
.B1(n_251),
.B2(n_272),
.Y(n_295)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_208),
.Y(n_299)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_209),
.Y(n_279)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_212),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_130),
.A2(n_105),
.B1(n_107),
.B2(n_119),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_139),
.Y(n_215)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_144),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_216),
.B(n_219),
.Y(n_298)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_218),
.Y(n_283)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_130),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_220),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_170),
.A2(n_81),
.B1(n_117),
.B2(n_114),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_126),
.B(n_0),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_223),
.B(n_276),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_129),
.A2(n_100),
.B1(n_98),
.B2(n_95),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_224),
.A2(n_225),
.B1(n_270),
.B2(n_133),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_228),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_191),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_229),
.B(n_230),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_170),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_231),
.B(n_236),
.Y(n_317)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_169),
.Y(n_232)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_232),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_234),
.Y(n_286)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_147),
.Y(n_235)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_235),
.Y(n_288)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_136),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_238),
.Y(n_328)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_239),
.Y(n_329)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_240),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_152),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_245),
.Y(n_290)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_145),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_244),
.A2(n_250),
.B1(n_254),
.B2(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_246),
.B(n_247),
.Y(n_313)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_176),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_178),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_248),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_177),
.A2(n_66),
.B1(n_60),
.B2(n_70),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_171),
.A2(n_52),
.B1(n_23),
.B2(n_22),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_252),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_175),
.A2(n_52),
.B1(n_23),
.B2(n_22),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_253),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_194),
.A2(n_22),
.B1(n_28),
.B2(n_5),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_255),
.Y(n_305)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_127),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_256),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_195),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_257),
.Y(n_310)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_258),
.Y(n_321)
);

OR2x2_ASAP7_75t_SL g316 ( 
.A(n_259),
.B(n_264),
.Y(n_316)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_127),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_260),
.Y(n_331)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_261),
.Y(n_332)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

CKINVDCx12_ASAP7_75t_R g303 ( 
.A(n_262),
.Y(n_303)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_199),
.A2(n_28),
.B(n_4),
.C(n_5),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_132),
.B(n_3),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_265),
.B(n_268),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_266),
.A2(n_267),
.B1(n_273),
.B2(n_275),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_179),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_135),
.B(n_197),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_277),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_128),
.A2(n_28),
.B1(n_5),
.B2(n_6),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_148),
.B(n_4),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_271),
.B(n_274),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_165),
.A2(n_28),
.B1(n_8),
.B2(n_9),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_184),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_163),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_163),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_182),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_140),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_278),
.A2(n_173),
.B(n_138),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_284),
.A2(n_324),
.B1(n_327),
.B2(n_7),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_213),
.B(n_181),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_293),
.A2(n_314),
.B(n_208),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_154),
.C(n_155),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_315),
.C(n_143),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_226),
.A2(n_233),
.B1(n_249),
.B2(n_242),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_304),
.A2(n_278),
.B1(n_270),
.B2(n_264),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_231),
.A2(n_142),
.B1(n_151),
.B2(n_137),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_306),
.A2(n_307),
.B1(n_141),
.B2(n_276),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_253),
.A2(n_151),
.B1(n_190),
.B2(n_137),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_242),
.B(n_182),
.C(n_149),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_222),
.B(n_168),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_318),
.B(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_227),
.B(n_202),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_211),
.A2(n_128),
.B1(n_205),
.B2(n_190),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_205),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_326),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_259),
.B(n_179),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_211),
.A2(n_204),
.B1(n_138),
.B2(n_162),
.Y(n_327)
);

AO22x1_ASAP7_75t_SL g335 ( 
.A1(n_225),
.A2(n_167),
.B1(n_162),
.B2(n_161),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_220),
.Y(n_349)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_330),
.Y(n_336)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_337),
.A2(n_342),
.B1(n_359),
.B2(n_374),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_338),
.B(n_339),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_313),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_304),
.A2(n_223),
.B1(n_167),
.B2(n_161),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_287),
.B(n_252),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_343),
.B(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_330),
.Y(n_344)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_310),
.A2(n_213),
.B1(n_145),
.B2(n_267),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_346),
.A2(n_349),
.B1(n_351),
.B2(n_360),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_347),
.B(n_356),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_348),
.A2(n_353),
.B(n_371),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_311),
.B(n_255),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_362),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_312),
.A2(n_258),
.B(n_239),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_312),
.A2(n_263),
.B1(n_261),
.B2(n_210),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_298),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_361),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_294),
.B(n_235),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_300),
.B(n_215),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_357),
.B(n_363),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_280),
.A2(n_141),
.B1(n_236),
.B2(n_218),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_295),
.A2(n_238),
.B1(n_232),
.B2(n_244),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_282),
.A2(n_141),
.B1(n_218),
.B2(n_236),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_298),
.Y(n_361)
);

NOR2x1p5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_262),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_320),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_313),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_369),
.Y(n_394)
);

AOI32xp33_ASAP7_75t_L g365 ( 
.A1(n_300),
.A2(n_217),
.A3(n_209),
.B1(n_240),
.B2(n_247),
.Y(n_365)
);

AOI32xp33_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_325),
.A3(n_320),
.B1(n_323),
.B2(n_332),
.Y(n_392)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_315),
.B(n_241),
.C(n_266),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_367),
.B(n_281),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_287),
.B(n_228),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_311),
.B(n_7),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_313),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_376),
.Y(n_403)
);

OAI21xp33_ASAP7_75t_SL g371 ( 
.A1(n_314),
.A2(n_326),
.B(n_293),
.Y(n_371)
);

O2A1O1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_293),
.A2(n_250),
.B(n_273),
.C(n_10),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_372),
.A2(n_379),
.B(n_285),
.Y(n_414)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_297),
.Y(n_373)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_295),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_378),
.B1(n_322),
.B2(n_302),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_323),
.B(n_8),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_377),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_284),
.A2(n_8),
.B1(n_10),
.B2(n_324),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_319),
.B(n_10),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_375),
.A2(n_310),
.B1(n_335),
.B2(n_318),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_398),
.B1(n_405),
.B2(n_413),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_337),
.A2(n_327),
.B1(n_290),
.B2(n_335),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_390),
.A2(n_415),
.B1(n_339),
.B2(n_370),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_392),
.A2(n_341),
.B(n_365),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_378),
.A2(n_335),
.B1(n_285),
.B2(n_308),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_343),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_407),
.Y(n_442)
);

MAJx2_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_290),
.C(n_316),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_367),
.C(n_362),
.Y(n_427)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_406),
.B(n_416),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_350),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_346),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_408),
.Y(n_435)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_290),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_286),
.C(n_302),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_376),
.B(n_352),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_412),
.B(n_414),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_349),
.A2(n_285),
.B1(n_328),
.B2(n_296),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_371),
.A2(n_328),
.B1(n_296),
.B2(n_332),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_352),
.B(n_333),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_357),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_427),
.C(n_430),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_418),
.A2(n_382),
.B1(n_385),
.B2(n_392),
.Y(n_451)
);

XOR2x2_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_341),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g454 ( 
.A1(n_420),
.A2(n_437),
.B(n_444),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_398),
.A2(n_359),
.B1(n_374),
.B2(n_342),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_422),
.A2(n_436),
.B1(n_445),
.B2(n_408),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_411),
.A2(n_368),
.B1(n_358),
.B2(n_360),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_423),
.Y(n_462)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_424),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_390),
.A2(n_381),
.B1(n_415),
.B2(n_382),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_426),
.A2(n_432),
.B1(n_443),
.B2(n_385),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_429),
.B(n_394),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_410),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_395),
.Y(n_431)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_381),
.A2(n_364),
.B1(n_355),
.B2(n_361),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_416),
.C(n_401),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_433),
.B(n_439),
.C(n_449),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_396),
.B(n_369),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_440),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_372),
.B1(n_348),
.B2(n_353),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_401),
.A2(n_354),
.B(n_362),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_391),
.B(n_362),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_413),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_399),
.B(n_379),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_441),
.B(n_402),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_407),
.A2(n_351),
.B1(n_372),
.B2(n_336),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_411),
.A2(n_345),
.B(n_344),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_380),
.A2(n_377),
.B1(n_373),
.B2(n_334),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_404),
.Y(n_446)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_393),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_389),
.Y(n_458)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_329),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_433),
.C(n_428),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_451),
.A2(n_452),
.B1(n_457),
.B2(n_466),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_453),
.A2(n_425),
.B(n_420),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_456),
.A2(n_463),
.B1(n_435),
.B2(n_429),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_414),
.B1(n_394),
.B2(n_403),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_458),
.B(n_469),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_444),
.A2(n_436),
.B(n_442),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_459),
.A2(n_454),
.B(n_451),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_441),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_461),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_419),
.A2(n_403),
.B1(n_389),
.B2(n_384),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_430),
.B(n_388),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_464),
.B(n_474),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_388),
.B1(n_386),
.B2(n_384),
.Y(n_466)
);

NOR2x1_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_386),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_471),
.B(n_476),
.C(n_477),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_472),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_434),
.B(n_331),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_331),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_427),
.B(n_428),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_420),
.B(n_281),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_417),
.B(n_402),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_443),
.A2(n_383),
.B1(n_340),
.B2(n_373),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_478),
.A2(n_334),
.B1(n_297),
.B2(n_301),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_425),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_435),
.Y(n_489)
);

XNOR2x1_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_449),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_481),
.B(n_437),
.Y(n_486)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_421),
.Y(n_482)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_482),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_452),
.A2(n_419),
.B1(n_422),
.B2(n_440),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_483),
.A2(n_496),
.B1(n_455),
.B2(n_475),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_484),
.B(n_504),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_485),
.A2(n_299),
.B1(n_292),
.B2(n_305),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_486),
.B(n_468),
.Y(n_514)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_489),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_491),
.A2(n_494),
.B(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_492),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_467),
.B(n_448),
.C(n_446),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_493),
.B(n_501),
.C(n_490),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_454),
.A2(n_445),
.B(n_438),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_460),
.Y(n_495)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_495),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_457),
.A2(n_431),
.B1(n_424),
.B2(n_421),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_482),
.Y(n_498)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_498),
.Y(n_534)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_460),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_499),
.A2(n_505),
.B1(n_507),
.B2(n_510),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_459),
.A2(n_383),
.B(n_340),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_500),
.A2(n_506),
.B(n_511),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_467),
.B(n_279),
.C(n_291),
.Y(n_501)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_479),
.B(n_309),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_462),
.A2(n_299),
.B(n_291),
.Y(n_508)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_465),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_455),
.B(n_309),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_512),
.B(n_515),
.C(n_517),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_481),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_513),
.B(n_484),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_514),
.B(n_516),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_501),
.B(n_471),
.C(n_474),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_486),
.B(n_468),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_490),
.B(n_477),
.C(n_464),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_476),
.C(n_466),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_522),
.C(n_526),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_463),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_519),
.B(n_531),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_491),
.B(n_456),
.C(n_478),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_500),
.B(n_496),
.Y(n_523)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_524),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_462),
.C(n_475),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_480),
.B1(n_470),
.B2(n_469),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_528),
.A2(n_509),
.B1(n_502),
.B2(n_492),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_497),
.A2(n_480),
.B1(n_470),
.B2(n_301),
.Y(n_529)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_529),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g531 ( 
.A(n_497),
.B(n_303),
.Y(n_531)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_535),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_533),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_542),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_523),
.B(n_489),
.Y(n_540)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_540),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_520),
.A2(n_502),
.B(n_485),
.Y(n_541)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_541),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_520),
.A2(n_509),
.B(n_488),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_545),
.A2(n_535),
.B1(n_526),
.B2(n_527),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g570 ( 
.A(n_546),
.B(n_554),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_512),
.B(n_488),
.C(n_508),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_552),
.Y(n_563)
);

AOI22x1_ASAP7_75t_L g551 ( 
.A1(n_523),
.A2(n_507),
.B1(n_487),
.B2(n_510),
.Y(n_551)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_551),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_528),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_524),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_553),
.A2(n_541),
.B1(n_539),
.B2(n_542),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_521),
.A2(n_504),
.B1(n_506),
.B2(n_511),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_537),
.B(n_515),
.C(n_513),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_555),
.B(n_556),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_544),
.A2(n_525),
.B1(n_530),
.B2(n_522),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_557),
.A2(n_562),
.B1(n_538),
.B2(n_548),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_516),
.C(n_517),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_558),
.B(n_560),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_514),
.C(n_519),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_543),
.B(n_518),
.C(n_531),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_561),
.B(n_564),
.C(n_566),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_538),
.A2(n_534),
.B1(n_532),
.B2(n_487),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_505),
.C(n_495),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_549),
.B(n_499),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_551),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_498),
.C(n_283),
.Y(n_566)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_571),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_570),
.B(n_546),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_574),
.B(n_321),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_575),
.A2(n_566),
.B1(n_561),
.B2(n_283),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_568),
.A2(n_540),
.B(n_539),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_576),
.A2(n_577),
.B(n_567),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_559),
.A2(n_569),
.B(n_557),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_555),
.B(n_547),
.C(n_548),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_578),
.B(n_582),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_563),
.A2(n_540),
.B1(n_551),
.B2(n_549),
.Y(n_580)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_580),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_564),
.B(n_305),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_562),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_583),
.A2(n_575),
.B1(n_579),
.B2(n_584),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_584),
.B(n_565),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_573),
.B(n_558),
.C(n_560),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_588),
.Y(n_596)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_586),
.Y(n_595)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_587),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_573),
.B(n_279),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_578),
.C(n_589),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_292),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_592),
.B(n_593),
.Y(n_598)
);

AO21x1_ASAP7_75t_L g599 ( 
.A1(n_594),
.A2(n_580),
.B(n_581),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_599),
.B(n_600),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_585),
.B(n_577),
.C(n_576),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_601),
.B(n_591),
.Y(n_603)
);

OAI321xp33_ASAP7_75t_L g607 ( 
.A1(n_603),
.A2(n_595),
.A3(n_598),
.B1(n_587),
.B2(n_333),
.C(n_329),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_596),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_604),
.A2(n_605),
.B(n_588),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_597),
.B(n_590),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_606),
.A2(n_607),
.B(n_598),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_608),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_609),
.B(n_602),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_299),
.B(n_321),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_303),
.C(n_292),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_612),
.A2(n_286),
.B1(n_289),
.B2(n_609),
.Y(n_613)
);


endmodule