module fake_jpeg_2759_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_0),
.B(n_1),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_41),
.A2(n_5),
.B(n_7),
.Y(n_111)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_10),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_47),
.B(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_50),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_62),
.Y(n_88)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_23),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g113 ( 
.A(n_59),
.Y(n_113)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_28),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_8),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_70),
.Y(n_118)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_18),
.B(n_2),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_3),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_5),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_77),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_17),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g116 ( 
.A(n_78),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_24),
.B1(n_27),
.B2(n_39),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_81),
.A2(n_89),
.B1(n_105),
.B2(n_64),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_114),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_24),
.B1(n_27),
.B2(n_38),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_61),
.B(n_20),
.C(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_100),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_20),
.C(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_46),
.B1(n_78),
.B2(n_57),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_75),
.A2(n_38),
.B1(n_7),
.B2(n_5),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_106),
.A2(n_45),
.B1(n_42),
.B2(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_9),
.Y(n_126)
);

CKINVDCx12_ASAP7_75t_R g112 ( 
.A(n_71),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_68),
.B(n_9),
.Y(n_114)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_127),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_141),
.B1(n_85),
.B2(n_94),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_63),
.B1(n_69),
.B2(n_60),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_125),
.B1(n_142),
.B2(n_134),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_89),
.B(n_90),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_118),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_128),
.Y(n_154)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_40),
.B(n_56),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_135),
.Y(n_149)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_79),
.B(n_78),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_147),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_113),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_134),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_117),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_137),
.Y(n_153)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_105),
.B(n_87),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_84),
.B1(n_97),
.B2(n_92),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_80),
.B1(n_95),
.B2(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_144),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_82),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_110),
.B1(n_102),
.B2(n_93),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_131),
.C(n_133),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_108),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_164),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_84),
.B1(n_104),
.B2(n_103),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_133),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_104),
.B1(n_122),
.B2(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_162),
.B1(n_165),
.B2(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_147),
.B1(n_124),
.B2(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_167),
.Y(n_182)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_169),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_151),
.B1(n_155),
.B2(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_176),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_166),
.B(n_140),
.Y(n_173)
);

XOR2x2_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_164),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_130),
.B1(n_123),
.B2(n_137),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_179),
.B1(n_181),
.B2(n_158),
.Y(n_191)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_178),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_143),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_159),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_149),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_146),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_191),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_151),
.B1(n_155),
.B2(n_161),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_130),
.B(n_149),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_180),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_157),
.B1(n_130),
.B2(n_156),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_172),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_184),
.B(n_173),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_197),
.B(n_201),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_154),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_202),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_200),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_180),
.C(n_168),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_183),
.Y(n_209)
);

AO32x1_ASAP7_75t_L g204 ( 
.A1(n_186),
.A2(n_169),
.A3(n_178),
.B1(n_175),
.B2(n_176),
.Y(n_204)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_190),
.CI(n_187),
.CON(n_208),
.SN(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_205),
.B(n_209),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_197),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_211),
.B(n_182),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_217),
.C(n_192),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_199),
.B1(n_182),
.B2(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_207),
.C(n_177),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_202),
.B(n_204),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_208),
.B(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_216),
.B(n_212),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_188),
.B(n_136),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_218),
.A2(n_203),
.A3(n_207),
.B1(n_188),
.B2(n_179),
.C1(n_156),
.C2(n_170),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_224),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_132),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_225),
.B(n_222),
.C(n_120),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_138),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_129),
.Y(n_231)
);


endmodule