module fake_jpeg_19129_n_205 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_27),
.Y(n_35)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_26),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_19),
.B1(n_13),
.B2(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_33),
.Y(n_57)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_49),
.Y(n_64)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_38),
.B1(n_28),
.B2(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_52),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_55),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_11),
.B(n_21),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_36),
.B1(n_37),
.B2(n_30),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_51),
.B1(n_24),
.B2(n_53),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_35),
.B(n_34),
.C(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_29),
.B(n_32),
.C(n_27),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_71),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_49),
.Y(n_72)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_51),
.B1(n_45),
.B2(n_54),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_29),
.B(n_1),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_83),
.A2(n_57),
.B(n_71),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_93),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_66),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_88),
.B(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_77),
.B(n_69),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_58),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_94),
.B(n_17),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_65),
.B(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_101),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_61),
.B1(n_58),
.B2(n_67),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_98),
.A2(n_56),
.B1(n_76),
.B2(n_75),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_68),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_62),
.B(n_70),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_74),
.B1(n_80),
.B2(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_91),
.B1(n_95),
.B2(n_15),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_109),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_100),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_114),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_115),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_95),
.B(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_76),
.B1(n_60),
.B2(n_67),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_113),
.B1(n_119),
.B2(n_99),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_67),
.B1(n_60),
.B2(n_19),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_88),
.B(n_29),
.Y(n_115)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_16),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_29),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.C(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_38),
.C(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_20),
.B1(n_18),
.B2(n_15),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_121),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_90),
.B(n_18),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_124),
.B(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_103),
.A2(n_22),
.B1(n_14),
.B2(n_17),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_22),
.B1(n_27),
.B2(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_27),
.C(n_12),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_123),
.C(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_139),
.A2(n_140),
.B(n_141),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_145),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_0),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_111),
.B(n_122),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_131),
.B(n_129),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_107),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_17),
.C(n_16),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_135),
.C(n_131),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_16),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_14),
.B1(n_6),
.B2(n_7),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_5),
.B(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_164),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_162),
.B(n_154),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_132),
.C(n_126),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_165),
.C(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_138),
.C(n_16),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_142),
.C(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_171),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_161),
.B(n_149),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_146),
.B1(n_149),
.B2(n_2),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_0),
.Y(n_183)
);

NOR2x1_ASAP7_75t_SL g173 ( 
.A(n_165),
.B(n_146),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_168),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_177),
.B(n_6),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_174),
.B(n_160),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_14),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_157),
.C(n_160),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_14),
.C(n_3),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_185),
.B1(n_4),
.B2(n_8),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_4),
.B(n_9),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_184),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_172),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_190),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_3),
.B(n_4),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_1),
.C(n_2),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_192),
.B(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_196),
.C(n_197),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_8),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_189),
.A2(n_0),
.B(n_1),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_1),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_198),
.C(n_195),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.C(n_200),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g205 ( 
.A(n_204),
.Y(n_205)
);


endmodule