module fake_jpeg_6046_n_25 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_16;
wire n_24;
wire n_17;
wire n_15;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_5),
.A2(n_13),
.B1(n_11),
.B2(n_1),
.Y(n_17)
);

OAI22xp33_ASAP7_75t_L g18 ( 
.A1(n_3),
.A2(n_9),
.B1(n_4),
.B2(n_2),
.Y(n_18)
);

AND2x4_ASAP7_75t_SL g19 ( 
.A(n_7),
.B(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

XOR2x2_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_16),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_18),
.A2(n_6),
.B1(n_17),
.B2(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_23),
.B(n_22),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_15),
.Y(n_25)
);


endmodule