module fake_jpeg_10258_n_228 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_46),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_50),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_28),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_20),
.Y(n_63)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_64)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_61),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_29),
.B1(n_27),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_55),
.A2(n_30),
.B1(n_19),
.B2(n_33),
.Y(n_103)
);

CKINVDCx9p33_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_23),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_69),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_29),
.B(n_28),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

AND2x4_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_29),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_36),
.B(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx4f_ASAP7_75t_SL g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_23),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_76),
.Y(n_79)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_94),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_43),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_93),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_86),
.B1(n_109),
.B2(n_83),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_86),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_45),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_88),
.B(n_89),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_31),
.B1(n_22),
.B2(n_33),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_102),
.B1(n_106),
.B2(n_53),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_22),
.B(n_31),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_34),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_101),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_34),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_28),
.B(n_18),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_57),
.B1(n_80),
.B2(n_62),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_65),
.B(n_19),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_19),
.B1(n_18),
.B2(n_28),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_0),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_1),
.Y(n_133)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_108),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_121),
.B1(n_129),
.B2(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_58),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_120),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_18),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_18),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_124),
.Y(n_143)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_102),
.B1(n_86),
.B2(n_85),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_87),
.B1(n_99),
.B2(n_108),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_86),
.A2(n_62),
.B1(n_74),
.B2(n_37),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_130),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_82),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_132),
.A2(n_94),
.B1(n_88),
.B2(n_104),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_93),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_127),
.B1(n_126),
.B2(n_113),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_139),
.B(n_152),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_91),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_81),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_1),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_111),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_151),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_112),
.A2(n_74),
.B(n_109),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_153),
.B(n_116),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_99),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g153 ( 
.A(n_112),
.B(n_81),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_126),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_126),
.B1(n_113),
.B2(n_133),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_163),
.B1(n_164),
.B2(n_170),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_159),
.A2(n_90),
.B1(n_142),
.B2(n_68),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_162),
.A2(n_168),
.B(n_172),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_127),
.B1(n_114),
.B2(n_122),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_135),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_169),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_87),
.B(n_90),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_110),
.B1(n_130),
.B2(n_76),
.Y(n_170)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_12),
.B1(n_16),
.B2(n_13),
.C(n_10),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_100),
.B(n_67),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_66),
.Y(n_173)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_145),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_149),
.C(n_153),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_179),
.C(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_143),
.B1(n_153),
.B2(n_152),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_186),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_157),
.B(n_140),
.C(n_150),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_136),
.C(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_164),
.B(n_146),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_185),
.B(n_189),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_134),
.A3(n_155),
.B1(n_148),
.B2(n_143),
.C1(n_138),
.C2(n_137),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_144),
.C(n_142),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_168),
.C(n_173),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_165),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_188),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_194),
.Y(n_201)
);

AOI211xp5_ASAP7_75t_SL g197 ( 
.A1(n_176),
.A2(n_163),
.B(n_162),
.C(n_170),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_178),
.B1(n_158),
.B2(n_175),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_183),
.C(n_179),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_203),
.A2(n_206),
.B1(n_194),
.B2(n_199),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_195),
.A2(n_176),
.B(n_180),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_207),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_165),
.Y(n_209)
);

XOR2x2_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_196),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_191),
.B1(n_199),
.B2(n_171),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_204),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_2),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_201),
.A3(n_212),
.B1(n_213),
.B2(n_209),
.C1(n_160),
.C2(n_12),
.Y(n_218)
);

AOI321xp33_ASAP7_75t_L g215 ( 
.A1(n_208),
.A2(n_190),
.A3(n_160),
.B1(n_169),
.B2(n_100),
.C(n_174),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_215),
.A2(n_190),
.B(n_205),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_218),
.A2(n_219),
.B(n_220),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_16),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_217),
.A2(n_214),
.B(n_10),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_4),
.C(n_5),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_224),
.A2(n_225),
.B(n_6),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_6),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_226),
.A2(n_7),
.A3(n_8),
.B1(n_100),
.B2(n_222),
.C1(n_203),
.C2(n_220),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_7),
.Y(n_228)
);


endmodule