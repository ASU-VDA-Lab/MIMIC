module real_jpeg_20398_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_0),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_0),
.A2(n_29),
.B1(n_71),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_0),
.A2(n_29),
.B1(n_45),
.B2(n_46),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_37),
.B1(n_71),
.B2(n_77),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_71),
.B1(n_77),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_2),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_95),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_95),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_95),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_71),
.B1(n_77),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_3),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_149),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_149),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_149),
.Y(n_202)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_70),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_6),
.A2(n_86),
.B(n_156),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_8),
.A2(n_71),
.B1(n_77),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_8),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_127),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_127),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_9),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_9),
.A2(n_14),
.B(n_33),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_147),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_9),
.A2(n_58),
.B1(n_202),
.B2(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_9),
.B(n_45),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_45),
.B(n_229),
.Y(n_233)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_11),
.A2(n_45),
.B1(n_46),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_117)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_28),
.B(n_31),
.C(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_130),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_20),
.B(n_104),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_82),
.B2(n_103),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_54),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_41),
.B(n_53),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_24),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_35),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_25),
.A2(n_39),
.B(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_26),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_43),
.B2(n_44),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_27),
.A2(n_34),
.B(n_147),
.C(n_194),
.Y(n_193)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_27),
.B(n_43),
.Y(n_230)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g228 ( 
.A1(n_28),
.A2(n_44),
.A3(n_46),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_30),
.B(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_31),
.A2(n_39),
.B1(n_63),
.B2(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_31),
.A2(n_35),
.B(n_91),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_31),
.A2(n_39),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_31),
.B(n_147),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_31),
.A2(n_39),
.B1(n_198),
.B2(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_31),
.A2(n_39),
.B1(n_220),
.B2(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_32),
.B(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_38),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_39),
.A2(n_63),
.B(n_64),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_39),
.A2(n_64),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_41)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_42),
.A2(n_48),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_42),
.A2(n_48),
.B1(n_143),
.B2(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_42),
.A2(n_48),
.B1(n_174),
.B2(n_233),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_45),
.Y(n_47)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_45),
.B(n_70),
.Y(n_153)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_46),
.A2(n_73),
.B1(n_146),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_49),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_48),
.B(n_122),
.Y(n_165)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_48),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_62),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_67),
.B1(n_80),
.B2(n_81),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_62),
.B1(n_81),
.B2(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B(n_60),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_58),
.A2(n_117),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_58),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_58),
.A2(n_188),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_58),
.A2(n_88),
.B(n_190),
.Y(n_221)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_59),
.B(n_147),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_61),
.A2(n_119),
.B(n_186),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_75),
.B(n_78),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_68),
.A2(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_94),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_68),
.A2(n_126),
.B1(n_128),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_69),
.A2(n_74),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

HAxp5_ASAP7_75t_SL g146 ( 
.A(n_71),
.B(n_147),
.CON(n_146),
.SN(n_146)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_74),
.B(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_74),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_92),
.C(n_97),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_90),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_84),
.B(n_90),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_89),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_93),
.B1(n_97),
.B2(n_98),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_121),
.B(n_123),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_100),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_279),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_108),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_110),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.C(n_124),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_111),
.A2(n_112),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_120),
.A2(n_124),
.B1(n_125),
.B2(n_271),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_120),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_147),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_275),
.B(n_280),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_178),
.B(n_260),
.C(n_274),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_167),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_133),
.B(n_167),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_150),
.B2(n_166),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_137),
.C(n_166),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_145),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_148),
.Y(n_161)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_158),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_151),
.B(n_159),
.C(n_163),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_168),
.B(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_172),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_175),
.C(n_176),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_173),
.B(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_175),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_259),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_253),
.B(n_258),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_241),
.B(n_252),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_223),
.B(n_240),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_211),
.B(n_222),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_199),
.B(n_210),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_191),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_191),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_205),
.B(n_209),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_221),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_219),
.C(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_225),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_231),
.B1(n_238),
.B2(n_239),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_232),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_237),
.C(n_238),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_242),
.B(n_243),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_248),
.B2(n_249),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_250),
.C(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_261),
.B(n_262),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_268),
.C(n_273),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_272),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);


endmodule