module fake_jpeg_5385_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_38),
.B(n_40),
.Y(n_85)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_49),
.A2(n_18),
.B1(n_16),
.B2(n_19),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_54),
.Y(n_64)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_13),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_61),
.Y(n_98)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_14),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_16),
.B1(n_19),
.B2(n_45),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_63),
.A2(n_71),
.B1(n_89),
.B2(n_93),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_66),
.A2(n_97),
.B1(n_33),
.B2(n_26),
.Y(n_135)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_77),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_70),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_53),
.A2(n_19),
.B1(n_16),
.B2(n_36),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_35),
.B(n_24),
.C(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_76),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_49),
.A2(n_36),
.B1(n_35),
.B2(n_24),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_78),
.A2(n_79),
.B1(n_95),
.B2(n_21),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_46),
.A2(n_29),
.B1(n_25),
.B2(n_31),
.Y(n_79)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_83),
.Y(n_122)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_86),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_29),
.C(n_25),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_33),
.Y(n_126)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_54),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_90),
.B(n_107),
.Y(n_136)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_52),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_94),
.A2(n_104),
.B1(n_33),
.B2(n_26),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_97)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_45),
.A2(n_32),
.B1(n_30),
.B2(n_22),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_38),
.B(n_33),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_38),
.B(n_14),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_121),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_32),
.B1(n_22),
.B2(n_21),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_130),
.B1(n_140),
.B2(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_0),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_117),
.B(n_89),
.Y(n_160)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_131),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_83),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_66),
.A2(n_21),
.B1(n_33),
.B2(n_26),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_73),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_133),
.Y(n_149)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_134),
.A2(n_109),
.B1(n_67),
.B2(n_26),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_81),
.B1(n_74),
.B2(n_80),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_137),
.Y(n_148)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_138),
.A2(n_139),
.B1(n_100),
.B2(n_101),
.Y(n_147)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_145),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_85),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_146),
.A2(n_173),
.B(n_159),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_96),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_176),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_152),
.A2(n_170),
.B1(n_175),
.B2(n_139),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_98),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_134),
.A2(n_104),
.B1(n_71),
.B2(n_94),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_169),
.B1(n_172),
.B2(n_178),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_106),
.B1(n_92),
.B2(n_100),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_158),
.B1(n_113),
.B2(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_162),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_130),
.B1(n_124),
.B2(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_124),
.B(n_62),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_160),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_142),
.A2(n_26),
.B(n_33),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_161),
.A2(n_137),
.B(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_165),
.Y(n_207)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_86),
.C(n_108),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_179),
.C(n_160),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_65),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_118),
.A2(n_77),
.B1(n_91),
.B2(n_74),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_119),
.B(n_81),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_173),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_80),
.B1(n_109),
.B2(n_67),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_143),
.B(n_0),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_86),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_174),
.B(n_137),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_108),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_123),
.B(n_14),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_6),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_115),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_153),
.C(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_182),
.Y(n_225)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_115),
.B1(n_131),
.B2(n_120),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_187),
.A2(n_212),
.B1(n_216),
.B2(n_7),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_188),
.A2(n_194),
.B1(n_202),
.B2(n_204),
.Y(n_227)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_200),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_83),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_206),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_209),
.C(n_210),
.Y(n_224)
);

AOI32xp33_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_128),
.A3(n_138),
.B1(n_133),
.B2(n_141),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_163),
.C(n_148),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_177),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_199),
.Y(n_238)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_201),
.B(n_211),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_156),
.A2(n_113),
.B1(n_129),
.B2(n_3),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_1),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_203),
.A2(n_205),
.B(n_151),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_158),
.A2(n_149),
.B1(n_157),
.B2(n_161),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_213),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_1),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_1),
.C(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_151),
.B(n_144),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_168),
.B(n_6),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_214),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_215),
.B(n_7),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_172),
.A2(n_178),
.B1(n_171),
.B2(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

AO21x2_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_164),
.B(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_221),
.A2(n_210),
.B1(n_211),
.B2(n_199),
.Y(n_268)
);

OAI21x1_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_205),
.B(n_184),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_196),
.B(n_200),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_213),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_148),
.Y(n_229)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_145),
.C(n_8),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_234),
.C(n_209),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_236),
.B1(n_240),
.B2(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_7),
.Y(n_233)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_233),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_7),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_181),
.Y(n_235)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_235),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_183),
.A2(n_190),
.B1(n_187),
.B2(n_216),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_241),
.Y(n_267)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_10),
.B1(n_11),
.B2(n_183),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_259),
.Y(n_269)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_251),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_256),
.C(n_257),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_190),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_234),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_260),
.C(n_224),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_221),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_203),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_220),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_262),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_236),
.A2(n_189),
.B1(n_203),
.B2(n_185),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_263),
.A2(n_268),
.B1(n_240),
.B2(n_227),
.Y(n_274)
);

XOR2x1_ASAP7_75t_L g264 ( 
.A(n_221),
.B(n_223),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_264),
.B(n_229),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_196),
.B(n_189),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_242),
.B1(n_226),
.B2(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_267),
.B(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_276),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_272),
.B(n_263),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_260),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_274),
.A2(n_266),
.B1(n_249),
.B2(n_227),
.Y(n_294)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_217),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_277),
.Y(n_293)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_280),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_254),
.B1(n_255),
.B2(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_282),
.C(n_258),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_224),
.C(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_220),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_284),
.A2(n_233),
.B(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_286),
.B(n_235),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_271),
.B(n_239),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_248),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_282),
.C(n_281),
.Y(n_306)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_246),
.B(n_286),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_297),
.B(n_300),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_298),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_294),
.A2(n_296),
.B1(n_272),
.B2(n_243),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_279),
.B1(n_285),
.B2(n_269),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_273),
.Y(n_298)
);

INVx11_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_287),
.B1(n_274),
.B2(n_290),
.Y(n_302)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_302),
.A2(n_292),
.B(n_228),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_270),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_284),
.B(n_250),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_308),
.B(n_312),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_307),
.C(n_247),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_278),
.C(n_280),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_257),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_238),
.Y(n_321)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_317),
.B(n_320),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_295),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_312),
.B(n_309),
.Y(n_324)
);

HAxp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_246),
.CON(n_317),
.SN(n_317)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_301),
.A2(n_283),
.B1(n_296),
.B2(n_294),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_318),
.A2(n_302),
.B1(n_308),
.B2(n_303),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_305),
.Y(n_323)
);

AO21x1_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_316),
.B(n_314),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_324),
.B(n_325),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_320),
.A2(n_307),
.B(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_326),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_328),
.A2(n_329),
.B(n_331),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_306),
.C(n_311),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_315),
.B(n_319),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_332),
.B(n_318),
.Y(n_335)
);

OAI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_317),
.B(n_321),
.Y(n_336)
);

AO21x2_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_305),
.B(n_265),
.Y(n_337)
);


endmodule