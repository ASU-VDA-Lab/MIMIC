module real_jpeg_3739_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_0),
.A2(n_44),
.B1(n_45),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_0),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_57),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_0),
.A2(n_57),
.B1(n_63),
.B2(n_65),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_1),
.A2(n_27),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_1),
.B(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_43),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_1),
.A2(n_35),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_1),
.B(n_60),
.C(n_63),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_44),
.B1(n_45),
.B2(n_125),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_1),
.B(n_78),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_69),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_54),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_2),
.A2(n_54),
.B1(n_63),
.B2(n_65),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_63),
.B1(n_65),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_5),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_80),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_63),
.B1(n_65),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_11),
.A2(n_63),
.B1(n_65),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_12),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_12),
.A2(n_39),
.B1(n_63),
.B2(n_65),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_13),
.A2(n_33),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_13),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_13),
.A2(n_51),
.B1(n_63),
.B2(n_65),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_14),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_114),
.B1(n_188),
.B2(n_189),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_19),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_113),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_93),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_84),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_22),
.B(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_23),
.B(n_41),
.C(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_24),
.A2(n_32),
.B1(n_38),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g73 ( 
.A1(n_28),
.A2(n_31),
.A3(n_35),
.B1(n_37),
.B2(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_33),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_32),
.Y(n_89)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_33),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_33),
.B(n_125),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI32xp33_ASAP7_75t_L g123 ( 
.A1(n_35),
.A2(n_45),
.A3(n_47),
.B1(n_124),
.B2(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_40)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_42),
.A2(n_50),
.B1(n_52),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_42),
.A2(n_52),
.B1(n_53),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_42),
.A2(n_52),
.B1(n_86),
.B2(n_147),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AO22x1_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_45),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_44),
.B(n_48),
.Y(n_126)
);

INVx5_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_45),
.B(n_156),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_47),
.Y(n_48)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_66),
.B2(n_69),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_56),
.A2(n_58),
.B1(n_69),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_58),
.A2(n_69),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_58),
.A2(n_69),
.B1(n_138),
.B2(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_62),
.A2(n_67),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_62),
.A2(n_110),
.B1(n_121),
.B2(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_63),
.B(n_166),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_84),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_75),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_76),
.A2(n_78),
.B1(n_129),
.B2(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_76),
.A2(n_78),
.B1(n_125),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_76),
.A2(n_78),
.B1(n_168),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_82),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_77),
.A2(n_106),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_77),
.A2(n_106),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.C(n_90),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_133),
.B(n_187),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_131),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_131),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_119),
.B(n_122),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_127),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_182),
.B(n_186),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_151),
.B(n_181),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_143),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_143),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_141),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_140),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_146),
.C(n_149),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_162),
.B(n_180),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_155),
.B1(n_157),
.B2(n_158),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_174),
.B(n_179),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_169),
.B(n_173),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_178),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_185),
.Y(n_186)
);


endmodule