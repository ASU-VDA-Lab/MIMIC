module fake_jpeg_31390_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_15),
.B(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_7),
.B(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_8),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_12),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_11),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_15),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_30),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_16),
.B1(n_17),
.B2(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_19),
.Y(n_32)
);

AO22x1_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_13),
.B1(n_9),
.B2(n_11),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_34),
.C(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_39),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_12),
.C(n_14),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_31),
.B1(n_33),
.B2(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_10),
.B(n_14),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_21),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.C(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_48),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_40),
.C(n_43),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_49),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_3),
.A3(n_4),
.B1(n_6),
.B2(n_21),
.C1(n_45),
.C2(n_49),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_3),
.Y(n_52)
);


endmodule