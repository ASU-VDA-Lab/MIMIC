module fake_ariane_1075_n_844 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_844);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_844;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_779;
wire n_731;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_804;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_767;
wire n_736;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g164 ( 
.A(n_24),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_40),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_42),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_21),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_104),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_106),
.Y(n_170)
);

BUFx2_ASAP7_75t_SL g171 ( 
.A(n_111),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_55),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_78),
.Y(n_173)
);

BUFx10_ASAP7_75t_L g174 ( 
.A(n_2),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_139),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_98),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_126),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_18),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_152),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_116),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_0),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_70),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_137),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_154),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_110),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_3),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_145),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_89),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_1),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_81),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_24),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_30),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_16),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_14),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_163),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_45),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_108),
.Y(n_207)
);

CKINVDCx12_ASAP7_75t_R g208 ( 
.A(n_122),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_29),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_83),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_76),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_48),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_60),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_57),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_71),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_65),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_20),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_92),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_67),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_52),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_86),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_84),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_143),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_133),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_8),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_172),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

NOR2xp67_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_228),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_175),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_187),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_200),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_174),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_166),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_206),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_182),
.Y(n_249)
);

INVxp33_ASAP7_75t_SL g250 ( 
.A(n_168),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_228),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_199),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_0),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_214),
.B(n_1),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_201),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_202),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_209),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_171),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_220),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_169),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_208),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_221),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_165),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_222),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_165),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_167),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_170),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_167),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_176),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_177),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_178),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_181),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_173),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_273),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_231),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_180),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_236),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_251),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_238),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_266),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_259),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_239),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_267),
.B(n_185),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_253),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_239),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_274),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_252),
.B(n_212),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_260),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_277),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_186),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_270),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_279),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

NAND2x1_ASAP7_75t_L g315 ( 
.A(n_237),
.B(n_212),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_275),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_275),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_234),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_256),
.Y(n_320)
);

AND2x4_ASAP7_75t_L g321 ( 
.A(n_230),
.B(n_212),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_264),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_240),
.B(n_2),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_246),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_248),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_254),
.B(n_188),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_255),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_262),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_250),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_268),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_285),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_329),
.B(n_250),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_R g336 ( 
.A(n_305),
.B(n_268),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_321),
.B(n_261),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_306),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_284),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_306),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_329),
.B(n_261),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_329),
.B(n_263),
.Y(n_342)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_294),
.B(n_212),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_329),
.B(n_263),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_212),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_329),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_284),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_241),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_189),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_294),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_294),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_295),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_309),
.B(n_241),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_295),
.B(n_191),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_283),
.B(n_192),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_295),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_194),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_295),
.B(n_198),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_290),
.Y(n_363)
);

OR2x6_ASAP7_75t_L g364 ( 
.A(n_304),
.B(n_3),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_308),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_301),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_203),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_317),
.B(n_204),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_308),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

AND2x4_ASAP7_75t_L g373 ( 
.A(n_321),
.B(n_4),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g374 ( 
.A1(n_320),
.A2(n_227),
.B1(n_226),
.B2(n_225),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g375 ( 
.A(n_282),
.B(n_4),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_288),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_313),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_328),
.B(n_205),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_296),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_313),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_315),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_292),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_293),
.A2(n_224),
.B1(n_223),
.B2(n_219),
.Y(n_383)
);

NAND2xp33_ASAP7_75t_L g384 ( 
.A(n_325),
.B(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_303),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_322),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_287),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_211),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_L g391 ( 
.A(n_331),
.B(n_213),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_286),
.B(n_330),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_L g393 ( 
.A(n_299),
.B(n_215),
.Y(n_393)
);

AO22x2_ASAP7_75t_L g394 ( 
.A1(n_319),
.A2(n_281),
.B1(n_324),
.B2(n_316),
.Y(n_394)
);

XNOR2x2_ASAP7_75t_SL g395 ( 
.A(n_324),
.B(n_5),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_287),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_289),
.A2(n_218),
.B1(n_216),
.B2(n_7),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_304),
.B(n_5),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_289),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_297),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_L g402 ( 
.A1(n_326),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_297),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_356),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_349),
.B(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_356),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_359),
.B(n_316),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_318),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_6),
.Y(n_410)
);

NAND2x1p5_ASAP7_75t_L g411 ( 
.A(n_352),
.B(n_332),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_389),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_337),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_350),
.A2(n_291),
.B(n_300),
.Y(n_415)
);

OAI221xp5_ASAP7_75t_L g416 ( 
.A1(n_402),
.A2(n_307),
.B1(n_318),
.B2(n_332),
.C(n_12),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_339),
.B(n_348),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_9),
.Y(n_418)
);

NAND3xp33_ASAP7_75t_SL g419 ( 
.A(n_348),
.B(n_312),
.C(n_302),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_351),
.Y(n_420)
);

AND2x6_ASAP7_75t_SL g421 ( 
.A(n_364),
.B(n_10),
.Y(n_421)
);

INVx8_ASAP7_75t_L g422 ( 
.A(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_338),
.B(n_10),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_373),
.B(n_11),
.Y(n_426)
);

OAI22xp33_ASAP7_75t_L g427 ( 
.A1(n_398),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_344),
.B(n_13),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_353),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_373),
.B(n_14),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_397),
.B(n_162),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_338),
.B(n_15),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_15),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_386),
.B(n_16),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_353),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_334),
.B(n_17),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_402),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_386),
.B(n_19),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_384),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_440)
);

AND2x6_ASAP7_75t_SL g441 ( 
.A(n_364),
.B(n_22),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_375),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_442)
);

BUFx8_ASAP7_75t_L g443 ( 
.A(n_367),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_344),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_336),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_23),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_333),
.Y(n_449)
);

NOR3xp33_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_25),
.C(n_26),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_352),
.B(n_355),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_344),
.Y(n_452)
);

AND2x6_ASAP7_75t_SL g453 ( 
.A(n_364),
.B(n_27),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_355),
.B(n_27),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_388),
.B(n_28),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

NAND2x1p5_ASAP7_75t_L g457 ( 
.A(n_347),
.B(n_28),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_361),
.B(n_376),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_385),
.B(n_29),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_387),
.B(n_30),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_371),
.B(n_31),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_354),
.B(n_31),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_32),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_354),
.B(n_32),
.Y(n_465)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_394),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_360),
.B(n_36),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_L g468 ( 
.A1(n_346),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_401),
.B(n_41),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_360),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_366),
.B(n_43),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_390),
.B(n_44),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_346),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_SL g475 ( 
.A(n_377),
.B(n_46),
.C(n_47),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_369),
.B(n_370),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_L g477 ( 
.A(n_380),
.B(n_49),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_422),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_407),
.B(n_400),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_414),
.B(n_341),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_459),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_405),
.B(n_403),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_417),
.B(n_342),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_443),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_444),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_412),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_420),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

OR2x4_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_395),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_443),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_456),
.Y(n_493)
);

NAND2x1p5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_366),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_425),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_408),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

OR2x6_ASAP7_75t_L g500 ( 
.A(n_422),
.B(n_366),
.Y(n_500)
);

BUFx4f_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_409),
.B(n_345),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_446),
.B(n_399),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_458),
.B(n_399),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_444),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_422),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_429),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_447),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_381),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_369),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_445),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_447),
.B(n_381),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_476),
.B(n_370),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_381),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_418),
.B(n_391),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_448),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_452),
.B(n_343),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_423),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_424),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_404),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_406),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_452),
.B(n_343),
.Y(n_527)
);

BUFx6f_ASAP7_75t_SL g528 ( 
.A(n_419),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_418),
.B(n_410),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_410),
.B(n_394),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_455),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_460),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_474),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_471),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_433),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g536 ( 
.A1(n_489),
.A2(n_474),
.B(n_473),
.Y(n_536)
);

AO31x2_ASAP7_75t_L g537 ( 
.A1(n_529),
.A2(n_464),
.A3(n_461),
.B(n_439),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_478),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_511),
.A2(n_516),
.B(n_518),
.Y(n_539)
);

OAI21xp33_ASAP7_75t_L g540 ( 
.A1(n_504),
.A2(n_464),
.B(n_438),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_480),
.B(n_436),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_531),
.A2(n_454),
.B(n_469),
.Y(n_542)
);

BUFx12f_ASAP7_75t_L g543 ( 
.A(n_486),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_532),
.B(n_471),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_479),
.B(n_428),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_489),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_483),
.B(n_436),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g548 ( 
.A1(n_535),
.A2(n_434),
.B(n_463),
.Y(n_548)
);

OAI21x1_ASAP7_75t_L g549 ( 
.A1(n_533),
.A2(n_467),
.B(n_472),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_496),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_483),
.B(n_394),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_500),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_502),
.B(n_461),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_496),
.A2(n_465),
.B(n_467),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_499),
.A2(n_472),
.B(n_457),
.Y(n_555)
);

OAI21x1_ASAP7_75t_L g556 ( 
.A1(n_499),
.A2(n_457),
.B(n_428),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_513),
.A2(n_451),
.B(n_432),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_515),
.B(n_426),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_515),
.B(n_430),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_482),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_515),
.A2(n_438),
.B1(n_442),
.B2(n_440),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

NAND3xp33_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_442),
.C(n_450),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_533),
.A2(n_466),
.B(n_468),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_525),
.A2(n_477),
.B(n_350),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_L g567 ( 
.A(n_485),
.B(n_416),
.C(n_415),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_513),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_484),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_491),
.A2(n_498),
.B1(n_395),
.B2(n_486),
.Y(n_570)
);

CKINVDCx11_ASAP7_75t_R g571 ( 
.A(n_498),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_530),
.B(n_374),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_512),
.Y(n_573)
);

NOR2x1_ASAP7_75t_L g574 ( 
.A(n_510),
.B(n_431),
.Y(n_574)
);

OAI21x1_ASAP7_75t_L g575 ( 
.A1(n_514),
.A2(n_466),
.B(n_358),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_525),
.A2(n_358),
.B(n_362),
.Y(n_576)
);

AO31x2_ASAP7_75t_L g577 ( 
.A1(n_514),
.A2(n_519),
.A3(n_522),
.B(n_497),
.Y(n_577)
);

AOI21x1_ASAP7_75t_L g578 ( 
.A1(n_488),
.A2(n_495),
.B(n_490),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_519),
.A2(n_362),
.B(n_475),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_530),
.A2(n_393),
.B(n_378),
.C(n_383),
.Y(n_580)
);

A2O1A1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_501),
.A2(n_524),
.B(n_522),
.C(n_521),
.Y(n_581)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_541),
.A2(n_501),
.B(n_383),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_577),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_557),
.A2(n_523),
.B(n_526),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_536),
.A2(n_523),
.B(n_494),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_539),
.B(n_517),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_554),
.A2(n_494),
.B(n_501),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_549),
.A2(n_534),
.B(n_507),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

O2A1O1Ixp33_ASAP7_75t_SL g590 ( 
.A1(n_553),
.A2(n_427),
.B(n_479),
.C(n_509),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_570),
.A2(n_491),
.B1(n_453),
.B2(n_421),
.Y(n_591)
);

O2A1O1Ixp5_ASAP7_75t_L g592 ( 
.A1(n_542),
.A2(n_487),
.B(n_505),
.C(n_510),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_546),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_549),
.A2(n_534),
.B(n_507),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_552),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_561),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_543),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

A2O1A1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_540),
.A2(n_521),
.B(n_517),
.C(n_510),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_564),
.B(n_508),
.C(n_506),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_567),
.A2(n_517),
.B(n_481),
.C(n_520),
.Y(n_601)
);

AOI21x1_ASAP7_75t_L g602 ( 
.A1(n_548),
.A2(n_527),
.B(n_520),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g603 ( 
.A1(n_562),
.A2(n_481),
.B(n_487),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_547),
.B(n_572),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_561),
.B(n_500),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_573),
.B(n_506),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_577),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_552),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_580),
.A2(n_508),
.B1(n_558),
.B2(n_559),
.Y(n_610)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_550),
.B(n_487),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_563),
.B(n_520),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_551),
.A2(n_481),
.B1(n_528),
.B2(n_493),
.Y(n_613)
);

AND2x2_ASAP7_75t_SL g614 ( 
.A(n_563),
.B(n_527),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_563),
.B(n_493),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_556),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_543),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_555),
.A2(n_575),
.B(n_579),
.Y(n_618)
);

AO21x2_ASAP7_75t_L g619 ( 
.A1(n_576),
.A2(n_527),
.B(n_343),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_571),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_563),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_571),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_550),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_565),
.A2(n_528),
.B1(n_441),
.B2(n_492),
.Y(n_625)
);

AOI221xp5_ASAP7_75t_L g626 ( 
.A1(n_591),
.A2(n_580),
.B1(n_528),
.B2(n_560),
.C(n_538),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_605),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_604),
.B(n_569),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_597),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_SL g630 ( 
.A(n_582),
.B(n_581),
.C(n_545),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_591),
.A2(n_565),
.B1(n_574),
.B2(n_544),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_593),
.Y(n_632)
);

AOI21xp33_ASAP7_75t_L g633 ( 
.A1(n_610),
.A2(n_565),
.B(n_544),
.Y(n_633)
);

OAI211xp5_ASAP7_75t_L g634 ( 
.A1(n_590),
.A2(n_492),
.B(n_566),
.C(n_581),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_618),
.A2(n_578),
.B(n_545),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_SL g636 ( 
.A1(n_603),
.A2(n_537),
.B1(n_568),
.B2(n_493),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_615),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_593),
.Y(n_638)
);

CKINVDCx6p67_ASAP7_75t_R g639 ( 
.A(n_622),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_625),
.A2(n_505),
.B1(n_493),
.B2(n_507),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_595),
.B(n_537),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_R g642 ( 
.A(n_605),
.B(n_568),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_604),
.A2(n_507),
.B1(n_537),
.B2(n_505),
.Y(n_643)
);

AOI22x1_ASAP7_75t_L g644 ( 
.A1(n_620),
.A2(n_537),
.B1(n_343),
.B2(n_577),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_605),
.B(n_615),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_600),
.A2(n_343),
.B1(n_51),
.B2(n_53),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_598),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_586),
.A2(n_50),
.B1(n_54),
.B2(n_56),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_598),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_615),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_623),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_L g652 ( 
.A1(n_606),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_586),
.B(n_62),
.Y(n_653)
);

INVx3_ASAP7_75t_SL g654 ( 
.A(n_597),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_618),
.A2(n_63),
.B(n_64),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_623),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_595),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_583),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_583),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_605),
.B(n_161),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_622),
.Y(n_661)
);

CKINVDCx8_ASAP7_75t_R g662 ( 
.A(n_617),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_607),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_SL g664 ( 
.A1(n_601),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_664)
);

CKINVDCx14_ASAP7_75t_R g665 ( 
.A(n_620),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_608),
.B(n_158),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_596),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_615),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_623),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_607),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_612),
.B(n_157),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_617),
.Y(n_672)
);

INVx3_ASAP7_75t_SL g673 ( 
.A(n_614),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_621),
.B(n_75),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_SL g675 ( 
.A1(n_599),
.A2(n_77),
.B(n_79),
.C(n_82),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_613),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_584),
.Y(n_677)
);

OAI211xp5_ASAP7_75t_L g678 ( 
.A1(n_626),
.A2(n_616),
.B(n_621),
.C(n_584),
.Y(n_678)
);

OAI221xp5_ASAP7_75t_SL g679 ( 
.A1(n_648),
.A2(n_612),
.B1(n_621),
.B2(n_589),
.C(n_609),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_640),
.A2(n_630),
.B1(n_628),
.B2(n_631),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_648),
.A2(n_614),
.B1(n_612),
.B2(n_596),
.Y(n_681)
);

AOI221xp5_ASAP7_75t_L g682 ( 
.A1(n_643),
.A2(n_624),
.B1(n_592),
.B2(n_623),
.C(n_616),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_634),
.A2(n_614),
.B1(n_596),
.B2(n_589),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_635),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_658),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_646),
.A2(n_612),
.B1(n_596),
.B2(n_611),
.Y(n_686)
);

AO21x2_ASAP7_75t_L g687 ( 
.A1(n_633),
.A2(n_624),
.B(n_588),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_645),
.Y(n_688)
);

OAI21xp33_ASAP7_75t_L g689 ( 
.A1(n_657),
.A2(n_616),
.B(n_602),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_666),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_661),
.B(n_612),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_641),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_659),
.Y(n_693)
);

AOI221xp5_ASAP7_75t_L g694 ( 
.A1(n_643),
.A2(n_623),
.B1(n_619),
.B2(n_609),
.C(n_584),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_630),
.A2(n_619),
.B1(n_611),
.B2(n_584),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_645),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_631),
.A2(n_619),
.B1(n_596),
.B2(n_609),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_638),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_673),
.A2(n_596),
.B1(n_585),
.B2(n_594),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_677),
.B(n_594),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_649),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_644),
.A2(n_671),
.B1(n_660),
.B2(n_653),
.Y(n_702)
);

BUFx2_ASAP7_75t_L g703 ( 
.A(n_677),
.Y(n_703)
);

AOI22xp33_ASAP7_75t_L g704 ( 
.A1(n_673),
.A2(n_585),
.B1(n_588),
.B2(n_587),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_SL g705 ( 
.A1(n_671),
.A2(n_587),
.B1(n_602),
.B2(n_93),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_627),
.Y(n_706)
);

OAI211xp5_ASAP7_75t_SL g707 ( 
.A1(n_662),
.A2(n_665),
.B(n_646),
.C(n_636),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_663),
.B(n_90),
.Y(n_708)
);

AOI222xp33_ASAP7_75t_L g709 ( 
.A1(n_676),
.A2(n_156),
.B1(n_94),
.B2(n_95),
.C1(n_96),
.C2(n_97),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_654),
.B(n_91),
.Y(n_710)
);

OAI211xp5_ASAP7_75t_L g711 ( 
.A1(n_636),
.A2(n_99),
.B(n_101),
.C(n_102),
.Y(n_711)
);

OAI21x1_ASAP7_75t_L g712 ( 
.A1(n_655),
.A2(n_656),
.B(n_669),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_660),
.A2(n_103),
.B1(n_105),
.B2(n_109),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_671),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_714)
);

BUFx12f_ASAP7_75t_L g715 ( 
.A(n_629),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_670),
.Y(n_716)
);

HB1xp67_ASAP7_75t_L g717 ( 
.A(n_637),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_692),
.B(n_685),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_716),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_685),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_692),
.B(n_651),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_703),
.B(n_650),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_693),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_700),
.B(n_650),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_700),
.B(n_668),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_L g727 ( 
.A1(n_707),
.A2(n_709),
.B(n_667),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_703),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_690),
.A2(n_660),
.B1(n_667),
.B2(n_676),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_693),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_698),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_717),
.B(n_701),
.Y(n_732)
);

BUFx2_ASAP7_75t_L g733 ( 
.A(n_684),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_684),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_689),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_684),
.B(n_637),
.Y(n_736)
);

AND2x4_ASAP7_75t_L g737 ( 
.A(n_706),
.B(n_668),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_687),
.B(n_647),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_712),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_712),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_687),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_687),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_688),
.B(n_627),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_708),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_694),
.B(n_632),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_706),
.Y(n_746)
);

AO21x2_ASAP7_75t_L g747 ( 
.A1(n_678),
.A2(n_664),
.B(n_675),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_728),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_719),
.Y(n_749)
);

AND2x6_ASAP7_75t_SL g750 ( 
.A(n_743),
.B(n_710),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_727),
.A2(n_686),
.B1(n_681),
.B2(n_708),
.Y(n_751)
);

NOR5xp2_ASAP7_75t_SL g752 ( 
.A(n_727),
.B(n_682),
.C(n_642),
.D(n_652),
.E(n_639),
.Y(n_752)
);

NOR2x1_ASAP7_75t_L g753 ( 
.A(n_718),
.B(n_629),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_719),
.Y(n_754)
);

OAI211xp5_ASAP7_75t_L g755 ( 
.A1(n_729),
.A2(n_680),
.B(n_714),
.C(n_702),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_725),
.B(n_696),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_719),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_718),
.B(n_696),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_747),
.A2(n_664),
.B(n_679),
.Y(n_759)
);

OAI211xp5_ASAP7_75t_L g760 ( 
.A1(n_735),
.A2(n_705),
.B(n_713),
.C(n_711),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_749),
.Y(n_761)
);

INVx6_ASAP7_75t_L g762 ( 
.A(n_750),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_748),
.Y(n_763)
);

OR2x2_ASAP7_75t_L g764 ( 
.A(n_758),
.B(n_728),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_753),
.B(n_654),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_756),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_748),
.Y(n_767)
);

OR2x2_ASAP7_75t_L g768 ( 
.A(n_754),
.B(n_732),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_757),
.B(n_732),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_768),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_766),
.B(n_726),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_SL g772 ( 
.A1(n_762),
.A2(n_759),
.B1(n_735),
.B2(n_744),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_762),
.B(n_715),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_769),
.B(n_764),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_765),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_771),
.B(n_763),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_775),
.B(n_763),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_770),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_774),
.B(n_767),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_773),
.B(n_726),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_780),
.B(n_773),
.Y(n_781)
);

OAI22xp33_ASAP7_75t_L g782 ( 
.A1(n_778),
.A2(n_751),
.B1(n_759),
.B2(n_772),
.Y(n_782)
);

INVxp67_ASAP7_75t_SL g783 ( 
.A(n_777),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_776),
.Y(n_784)
);

OAI211xp5_ASAP7_75t_SL g785 ( 
.A1(n_783),
.A2(n_755),
.B(n_760),
.C(n_777),
.Y(n_785)
);

AOI321xp33_ASAP7_75t_L g786 ( 
.A1(n_782),
.A2(n_755),
.A3(n_760),
.B1(n_776),
.B2(n_752),
.C(n_779),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_785),
.B(n_783),
.Y(n_787)
);

NAND4xp25_ASAP7_75t_L g788 ( 
.A(n_786),
.B(n_781),
.C(n_784),
.D(n_733),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_785),
.B(n_731),
.Y(n_789)
);

INVx2_ASAP7_75t_SL g790 ( 
.A(n_787),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_788),
.B(n_672),
.C(n_731),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_789),
.B(n_720),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_787),
.B(n_720),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_789),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_789),
.Y(n_795)
);

AOI221x1_ASAP7_75t_L g796 ( 
.A1(n_791),
.A2(n_674),
.B1(n_742),
.B2(n_741),
.C(n_724),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_790),
.A2(n_747),
.B(n_744),
.C(n_741),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_794),
.B(n_795),
.C(n_793),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_SL g799 ( 
.A1(n_792),
.A2(n_715),
.B(n_733),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_SL g800 ( 
.A(n_790),
.B(n_706),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_791),
.A2(n_739),
.B(n_683),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_798),
.B(n_726),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_797),
.A2(n_747),
.B(n_739),
.Y(n_803)
);

AOI222xp33_ASAP7_75t_L g804 ( 
.A1(n_800),
.A2(n_742),
.B1(n_745),
.B2(n_738),
.C1(n_761),
.C2(n_697),
.Y(n_804)
);

NOR2x1_ASAP7_75t_L g805 ( 
.A(n_799),
.B(n_747),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_796),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_801),
.A2(n_746),
.B(n_739),
.Y(n_807)
);

NAND3xp33_ASAP7_75t_SL g808 ( 
.A(n_798),
.B(n_691),
.C(n_723),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_806),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_802),
.Y(n_810)
);

NAND5xp2_ASAP7_75t_L g811 ( 
.A(n_807),
.B(n_736),
.C(n_725),
.D(n_724),
.E(n_730),
.Y(n_811)
);

NAND4xp75_ASAP7_75t_L g812 ( 
.A(n_805),
.B(n_721),
.C(n_736),
.D(n_730),
.Y(n_812)
);

NAND4xp75_ASAP7_75t_L g813 ( 
.A(n_803),
.B(n_721),
.C(n_736),
.D(n_746),
.Y(n_813)
);

NOR3xp33_ASAP7_75t_L g814 ( 
.A(n_808),
.B(n_740),
.C(n_746),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_804),
.B(n_734),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_L g816 ( 
.A(n_806),
.B(n_740),
.C(n_745),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_802),
.A2(n_734),
.B1(n_723),
.B2(n_740),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_810),
.B(n_734),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_809),
.A2(n_737),
.B(n_738),
.Y(n_819)
);

NOR3xp33_ASAP7_75t_L g820 ( 
.A(n_816),
.B(n_738),
.C(n_745),
.Y(n_820)
);

OAI211xp5_ASAP7_75t_SL g821 ( 
.A1(n_814),
.A2(n_695),
.B(n_699),
.C(n_704),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_811),
.A2(n_737),
.B(n_743),
.Y(n_822)
);

AOI221xp5_ASAP7_75t_L g823 ( 
.A1(n_817),
.A2(n_722),
.B1(n_737),
.B2(n_706),
.C(n_688),
.Y(n_823)
);

NAND5xp2_ASAP7_75t_L g824 ( 
.A(n_815),
.B(n_115),
.C(n_117),
.D(n_118),
.E(n_119),
.Y(n_824)
);

AOI211x1_ASAP7_75t_L g825 ( 
.A1(n_813),
.A2(n_812),
.B(n_737),
.C(n_124),
.Y(n_825)
);

NOR4xp25_ASAP7_75t_L g826 ( 
.A(n_810),
.B(n_722),
.C(n_123),
.D(n_125),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_SL g827 ( 
.A(n_809),
.B(n_722),
.C(n_127),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_827),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_SL g829 ( 
.A(n_826),
.B(n_120),
.C(n_128),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_818),
.Y(n_830)
);

XNOR2xp5_ASAP7_75t_L g831 ( 
.A(n_825),
.B(n_129),
.Y(n_831)
);

BUFx2_ASAP7_75t_L g832 ( 
.A(n_823),
.Y(n_832)
);

OR3x2_ASAP7_75t_L g833 ( 
.A(n_824),
.B(n_130),
.C(n_131),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_820),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_831),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_828),
.A2(n_819),
.B1(n_822),
.B2(n_821),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_830),
.B(n_832),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_837),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_838),
.B(n_835),
.Y(n_839)
);

AOI222xp33_ASAP7_75t_L g840 ( 
.A1(n_839),
.A2(n_836),
.B1(n_829),
.B2(n_834),
.C1(n_833),
.C2(n_706),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_840),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_132),
.B(n_134),
.Y(n_842)
);

AOI221xp5_ASAP7_75t_L g843 ( 
.A1(n_842),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.C(n_147),
.Y(n_843)
);

AOI211xp5_ASAP7_75t_L g844 ( 
.A1(n_843),
.A2(n_148),
.B(n_149),
.C(n_150),
.Y(n_844)
);


endmodule