module fake_jpeg_27834_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_31),
.Y(n_52)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_52),
.Y(n_68)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_31),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_45),
.A2(n_56),
.B(n_41),
.C(n_16),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_18),
.B1(n_19),
.B2(n_28),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_31),
.C(n_19),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_18),
.C(n_30),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_25),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_40),
.B1(n_33),
.B2(n_35),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_62),
.B(n_64),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_27),
.B(n_20),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_79),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_36),
.B1(n_18),
.B2(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_66),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_74),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_70),
.B(n_71),
.Y(n_103)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_44),
.Y(n_72)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_73),
.A2(n_75),
.B1(n_77),
.B2(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_43),
.A2(n_29),
.B1(n_25),
.B2(n_27),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_20),
.B1(n_16),
.B2(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_53),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_17),
.C(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_17),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_54),
.B1(n_45),
.B2(n_57),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_104),
.B1(n_73),
.B2(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_98),
.B1(n_72),
.B2(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_46),
.B1(n_51),
.B2(n_24),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_101),
.A2(n_105),
.B(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_24),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_32),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_65),
.Y(n_106)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_1),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_1),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_2),
.B(n_4),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_122),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_68),
.C(n_85),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_119),
.C(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_106),
.B1(n_103),
.B2(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_63),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_69),
.C(n_60),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_88),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_128),
.B(n_109),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_65),
.B1(n_74),
.B2(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_86),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_64),
.B1(n_60),
.B2(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR4xp25_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_61),
.C(n_4),
.D(n_5),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

NAND2x1_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_101),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_107),
.B(n_105),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_126),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_118),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g136 ( 
.A1(n_130),
.A2(n_99),
.A3(n_101),
.B1(n_108),
.B2(n_107),
.C1(n_91),
.C2(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_140),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_139),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_99),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_95),
.C(n_98),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_146),
.C(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_148),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_104),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_105),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

AO221x1_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_96),
.B1(n_61),
.B2(n_117),
.C(n_125),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_115),
.B1(n_114),
.B2(n_110),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_161),
.B1(n_144),
.B2(n_149),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_118),
.C(n_127),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_160),
.C(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_158),
.B(n_162),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_113),
.C(n_114),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_144),
.B1(n_132),
.B2(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_113),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_116),
.C(n_123),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_156),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_159),
.C(n_151),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_173),
.C(n_174),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_147),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_172),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_164),
.B(n_140),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_157),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_141),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_150),
.C(n_135),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_163),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_177),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_154),
.B1(n_150),
.B2(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_179),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_175),
.A2(n_171),
.B1(n_161),
.B2(n_129),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_180),
.A2(n_186),
.B(n_2),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_183),
.Y(n_187)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_176),
.Y(n_183)
);

AOI211xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_128),
.B(n_122),
.C(n_121),
.Y(n_186)
);

OAI31xp33_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_166),
.A3(n_170),
.B(n_173),
.Y(n_188)
);

OAI321xp33_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_189),
.A3(n_186),
.B1(n_185),
.B2(n_8),
.C(n_9),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_182),
.A2(n_166),
.B(n_15),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_5),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.C(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_15),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_198),
.Y(n_199)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_197),
.B(n_8),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_193),
.C(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_187),
.C(n_10),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_188),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.C(n_12),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_196),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_202),
.A2(n_199),
.B(n_12),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);


endmodule