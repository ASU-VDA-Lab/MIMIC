module real_jpeg_1035_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_1),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_71),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_1),
.A2(n_33),
.B1(n_36),
.B2(n_71),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_2),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_2),
.A2(n_52),
.B1(n_67),
.B2(n_68),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_2),
.A2(n_33),
.B1(n_36),
.B2(n_52),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_6),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_33),
.C(n_48),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_8),
.A2(n_35),
.B1(n_50),
.B2(n_53),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_8),
.B(n_46),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_8),
.A2(n_35),
.B1(n_67),
.B2(n_68),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_8),
.B(n_26),
.C(n_28),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_68),
.C(n_88),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_8),
.B(n_24),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_8),
.B(n_65),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_139),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_33),
.B1(n_36),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_10),
.A2(n_41),
.B1(n_50),
.B2(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_41),
.B1(n_67),
.B2(n_68),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_253),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_230),
.B(n_251),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_207),
.B(n_227),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_124),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_108),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_18),
.B(n_108),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_75),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_19),
.B(n_76),
.C(n_100),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_44),
.B2(n_58),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_21),
.B(n_58),
.C(n_59),
.Y(n_210)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_32),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_40),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_24),
.A2(n_32),
.B(n_157),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_24),
.A2(n_96),
.B(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_25),
.B(n_97),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_25)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_26),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_27),
.A2(n_28),
.B1(n_87),
.B2(n_88),
.Y(n_92)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2x1_ASAP7_75t_SL g165 ( 
.A(n_28),
.B(n_166),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_32),
.B(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_33),
.B(n_134),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_38),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_42),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_42),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_54),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_46),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_46),
.B(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_46),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_56)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_49),
.B(n_55),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_62),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_54),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_72),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_64),
.B(n_73),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_64),
.A2(n_74),
.B(n_123),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_64),
.B(n_174),
.Y(n_188)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_65),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_66),
.A2(n_74),
.B(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_68),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_68),
.B(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_72),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_72),
.B(n_170),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_74),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_100),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_83),
.C(n_95),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_79),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_81),
.A2(n_82),
.B(n_266),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_82),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_84),
.B1(n_95),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21x1_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_90),
.B(n_93),
.Y(n_84)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_85),
.A2(n_154),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_90),
.A2(n_106),
.B(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_91),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_91),
.B(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_94),
.B(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_101),
.B(n_104),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_102),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_103),
.B(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_105),
.B(n_153),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_106),
.B(n_140),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_115),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_110),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_115),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.C(n_119),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_117),
.B(n_245),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_122),
.B(n_188),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_145),
.B(n_206),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_142),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_126),
.B(n_142),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.C(n_136),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_127),
.A2(n_128),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_136),
.B1(n_137),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_135),
.A2(n_159),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_135),
.B(n_248),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_135),
.A2(n_159),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_138),
.B(n_154),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_139),
.B(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_160),
.B(n_205),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_147),
.B(n_151),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_148),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_158),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_200),
.B(n_204),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_182),
.B(n_199),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_175),
.B1(n_176),
.B2(n_181),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_178),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_179),
.C(n_181),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_189),
.B(n_198),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_186),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_197),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_202),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_226),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_212),
.C(n_222),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_221),
.B2(n_222),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_218),
.C(n_219),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_250),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_250),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_235),
.C(n_247),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_246),
.B2(n_247),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_239),
.C(n_244),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_248),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_273),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_257),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_267),
.B2(n_268),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B(n_272),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);


endmodule