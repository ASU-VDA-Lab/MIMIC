module fake_jpeg_9265_n_116 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx13_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx11_ASAP7_75t_SL g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_30),
.Y(n_32)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_24),
.A2(n_30),
.B(n_29),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_25),
.B(n_30),
.Y(n_43)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_24),
.A2(n_13),
.B1(n_11),
.B2(n_16),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_13),
.B1(n_25),
.B2(n_19),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_20),
.B(n_12),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_45),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_33),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_47),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_52),
.B1(n_55),
.B2(n_33),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_12),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_25),
.B1(n_28),
.B2(n_26),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_58),
.Y(n_78)
);

A2O1A1O1Ixp25_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_41),
.B(n_18),
.C(n_27),
.D(n_26),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_51),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_34),
.B1(n_38),
.B2(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_10),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_52),
.A2(n_34),
.B1(n_39),
.B2(n_36),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_67),
.C(n_68),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_21),
.B(n_16),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_37),
.C(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_51),
.B1(n_54),
.B2(n_17),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_57),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_0),
.Y(n_79)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_79),
.B(n_0),
.CI(n_2),
.CON(n_83),
.SN(n_83)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_57),
.B1(n_67),
.B2(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_86),
.B1(n_60),
.B2(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_87),
.Y(n_90)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_71),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_91),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_70),
.C(n_78),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_97),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_69),
.B1(n_70),
.B2(n_62),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_60),
.B1(n_65),
.B2(n_14),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_95),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_102),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_85),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_86),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_91),
.C(n_83),
.Y(n_107)
);

AOI31xp67_ASAP7_75t_SL g104 ( 
.A1(n_101),
.A2(n_90),
.A3(n_88),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_98),
.A2(n_93),
.B1(n_94),
.B2(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_2),
.Y(n_109)
);

NOR2xp67_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_99),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_108),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_105),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_111),
.A2(n_112),
.B(n_110),
.Y(n_113)
);

MAJx2_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_3),
.C(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_5),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_5),
.CI(n_113),
.CON(n_116),
.SN(n_116)
);


endmodule