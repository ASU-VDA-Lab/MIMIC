module fake_jpeg_356_n_394 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_394);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_394;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_46),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx4f_ASAP7_75t_SL g135 ( 
.A(n_50),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_51),
.B(n_52),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_56),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_55),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_13),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_40),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_79),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_64),
.Y(n_105)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_66),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_76),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_R g76 ( 
.A(n_18),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_20),
.Y(n_81)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_12),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_21),
.B1(n_20),
.B2(n_33),
.Y(n_94)
);

OA22x2_ASAP7_75t_L g158 ( 
.A1(n_94),
.A2(n_114),
.B1(n_132),
.B2(n_29),
.Y(n_158)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_57),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_45),
.A2(n_29),
.B1(n_26),
.B2(n_19),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_115),
.B(n_109),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_124),
.B1(n_133),
.B2(n_94),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_43),
.B1(n_39),
.B2(n_31),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_42),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_61),
.A2(n_16),
.B1(n_28),
.B2(n_23),
.Y(n_133)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_91),
.B(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_139),
.B(n_140),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_149),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_86),
.B(n_76),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_142),
.B(n_155),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_58),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_156),
.C(n_160),
.Y(n_199)
);

INVx11_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_163),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_161),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_49),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_99),
.B(n_66),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_98),
.A2(n_63),
.B1(n_23),
.B2(n_28),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_157),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_158),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_96),
.B(n_83),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_98),
.B(n_84),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_26),
.Y(n_163)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g182 ( 
.A(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_42),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_168),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_24),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_24),
.B(n_19),
.C(n_82),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_169),
.A2(n_37),
.B(n_41),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_124),
.B(n_47),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_171),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_73),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_172),
.A2(n_175),
.B1(n_93),
.B2(n_89),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_108),
.B(n_77),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_173),
.B(n_136),
.Y(n_191)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_90),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_118),
.A2(n_72),
.B1(n_69),
.B2(n_78),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_87),
.A2(n_70),
.B1(n_62),
.B2(n_55),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_179),
.A2(n_127),
.B1(n_88),
.B2(n_104),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_101),
.A2(n_53),
.B1(n_44),
.B2(n_67),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_37),
.B(n_41),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_183),
.A2(n_209),
.B1(n_214),
.B2(n_162),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_186),
.A2(n_197),
.B1(n_205),
.B2(n_208),
.Y(n_242)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_92),
.B1(n_101),
.B2(n_119),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_191),
.B(n_151),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_SL g195 ( 
.A1(n_158),
.A2(n_129),
.B(n_119),
.C(n_117),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_195),
.A2(n_160),
.B(n_156),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_127),
.B1(n_88),
.B2(n_122),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_200),
.A2(n_209),
.B(n_204),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_144),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_104),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_204),
.B(n_212),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_74),
.B1(n_65),
.B2(n_110),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_1),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_217),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_37),
.B1(n_41),
.B2(n_5),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_41),
.B1(n_3),
.B2(n_6),
.Y(n_209)
);

OR2x6_ASAP7_75t_SL g212 ( 
.A(n_142),
.B(n_41),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_14),
.B1(n_10),
.B2(n_7),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_161),
.B(n_2),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_213),
.B(n_207),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_220),
.A2(n_233),
.B(n_248),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_142),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_228),
.C(n_240),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_224),
.B1(n_232),
.B2(n_215),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_145),
.B1(n_165),
.B2(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_185),
.B(n_199),
.C(n_218),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_185),
.B(n_155),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_208),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_196),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_235),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_155),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_236),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_148),
.B1(n_147),
.B2(n_167),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_162),
.B(n_154),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_234),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_192),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_151),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_247),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_238),
.Y(n_262)
);

XOR2x2_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_160),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_159),
.C(n_137),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_156),
.C(n_166),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_243),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_210),
.C(n_196),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_245),
.C(n_143),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_138),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_212),
.A2(n_154),
.B(n_137),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_184),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_193),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_252),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_259),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_201),
.B1(n_215),
.B2(n_195),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_256),
.A2(n_267),
.B1(n_223),
.B2(n_249),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_190),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_212),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_261),
.B(n_263),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_194),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_231),
.C(n_240),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_236),
.A2(n_195),
.B1(n_214),
.B2(n_183),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_250),
.A2(n_189),
.B1(n_187),
.B2(n_182),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_246),
.A2(n_197),
.B1(n_205),
.B2(n_200),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_272),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_224),
.A2(n_189),
.B1(n_146),
.B2(n_178),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_242),
.A2(n_198),
.B1(n_182),
.B2(n_211),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_273),
.A2(n_236),
.B1(n_250),
.B2(n_222),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_246),
.A2(n_198),
.B1(n_138),
.B2(n_176),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_280),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_221),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_252),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_248),
.B(n_238),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_281),
.A2(n_304),
.B(n_276),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_265),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_289),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_232),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_268),
.B(n_257),
.Y(n_310)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_297),
.B1(n_257),
.B2(n_280),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_279),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_288),
.B(n_290),
.Y(n_305)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_244),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_293),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_294),
.A2(n_263),
.B1(n_278),
.B2(n_271),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_301),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_267),
.A2(n_223),
.B1(n_231),
.B2(n_241),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_229),
.C(n_245),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_298),
.B(n_299),
.C(n_261),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_256),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_226),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_303),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_262),
.A2(n_225),
.B(n_227),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_281),
.A2(n_268),
.B(n_257),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_306),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_308),
.B(n_323),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_310),
.Y(n_332)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_270),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_313),
.B(n_317),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_316),
.B(n_319),
.C(n_325),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_291),
.B(n_266),
.C(n_264),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_234),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_322),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_297),
.A2(n_277),
.B1(n_260),
.B2(n_225),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_324),
.C(n_304),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_277),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_291),
.B(n_260),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_174),
.B1(n_143),
.B2(n_159),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_292),
.B(n_2),
.C(n_3),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_299),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_340),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_334),
.B(n_325),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_319),
.B(n_298),
.C(n_293),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_336),
.B(n_337),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_301),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_295),
.C(n_282),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_339),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_312),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_294),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_323),
.B(n_296),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_341),
.B(n_317),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_300),
.C(n_296),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_343),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_342),
.B(n_283),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_344),
.B(n_345),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_338),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_347),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_348),
.A2(n_351),
.B1(n_354),
.B2(n_315),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_350),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_340),
.B(n_310),
.Y(n_350)
);

AO221x1_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_321),
.B1(n_327),
.B2(n_335),
.C(n_318),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_327),
.Y(n_352)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_352),
.Y(n_366)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_332),
.Y(n_353)
);

BUFx4f_ASAP7_75t_SL g365 ( 
.A(n_353),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_326),
.A2(n_286),
.B1(n_306),
.B2(n_309),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_357),
.A2(n_326),
.B(n_309),
.Y(n_358)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_355),
.A2(n_287),
.B1(n_324),
.B2(n_315),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_368),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_346),
.B(n_328),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_363),
.Y(n_371)
);

XOR2x2_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_328),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_364),
.B(n_354),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_356),
.B(n_331),
.C(n_341),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_367),
.B(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_373),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_370),
.B(n_374),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_331),
.C(n_348),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_365),
.B(n_303),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_284),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_377),
.C(n_363),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_289),
.Y(n_377)
);

XNOR2x1_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_359),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_378),
.B(n_359),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_372),
.A2(n_358),
.B(n_366),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_379),
.A2(n_374),
.B(n_370),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_381),
.B(n_383),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_361),
.C(n_346),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_380),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_384),
.A2(n_387),
.B(n_382),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_349),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_388),
.A2(n_389),
.B1(n_385),
.B2(n_382),
.Y(n_390)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_390),
.A2(n_302),
.B(n_7),
.C(n_8),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_391),
.A2(n_2),
.B(n_7),
.Y(n_392)
);

O2A1O1Ixp33_ASAP7_75t_SL g393 ( 
.A1(n_392),
.A2(n_9),
.B(n_2),
.C(n_8),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_8),
.Y(n_394)
);


endmodule