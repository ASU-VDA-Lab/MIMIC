module real_aes_8618_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_0), .A2(n_60), .B1(n_452), .B2(n_457), .Y(n_451) );
INVx1_ASAP7_75t_L g115 ( .A(n_1), .Y(n_115) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_2), .A2(n_29), .B1(n_105), .B2(n_153), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_3), .B(n_125), .Y(n_133) );
AND2x6_ASAP7_75t_L g120 ( .A(n_4), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g535 ( .A(n_4), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_4), .B(n_540), .Y(n_539) );
AO22x2_ASAP7_75t_L g441 ( .A1(n_5), .A2(n_25), .B1(n_433), .B2(n_438), .Y(n_441) );
INVx1_ASAP7_75t_L g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g99 ( .A(n_7), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_8), .B(n_101), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_9), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_10), .B(n_92), .Y(n_199) );
AO32x2_ASAP7_75t_L g169 ( .A1(n_11), .A2(n_91), .A3(n_125), .B1(n_144), .B2(n_170), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_12), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_13), .B(n_105), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_14), .B(n_92), .Y(n_122) );
AO22x2_ASAP7_75t_L g443 ( .A1(n_15), .A2(n_28), .B1(n_433), .B2(n_434), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_16), .A2(n_41), .B1(n_105), .B2(n_153), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g155 ( .A1(n_17), .A2(n_63), .B1(n_101), .B2(n_105), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_18), .B(n_105), .Y(n_185) );
INVx1_ASAP7_75t_L g546 ( .A(n_18), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_19), .A2(n_424), .B1(n_522), .B2(n_523), .Y(n_423) );
INVx1_ASAP7_75t_L g522 ( .A(n_19), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_20), .B(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g110 ( .A(n_21), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_22), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_23), .B(n_146), .Y(n_187) );
INVx2_ASAP7_75t_L g103 ( .A(n_24), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_26), .B(n_105), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_27), .B(n_146), .Y(n_168) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_28), .A2(n_47), .B1(n_58), .B2(n_528), .C(n_529), .Y(n_527) );
INVxp67_ASAP7_75t_L g530 ( .A(n_28), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_29), .A2(n_76), .B1(n_418), .B2(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_29), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_30), .A2(n_415), .B1(n_416), .B2(n_422), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_30), .Y(n_415) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_31), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_32), .A2(n_61), .B1(n_474), .B2(n_478), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_33), .B(n_105), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_34), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g152 ( .A1(n_35), .A2(n_72), .B1(n_153), .B2(n_154), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_36), .B(n_105), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_37), .B(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_38), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_39), .A2(n_424), .B1(n_523), .B2(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_39), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_40), .B(n_113), .Y(n_132) );
AOI22xp33_ASAP7_75t_SL g197 ( .A1(n_42), .A2(n_49), .B1(n_101), .B2(n_105), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_43), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g410 ( .A1(n_44), .A2(n_64), .B1(n_411), .B2(n_412), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g411 ( .A(n_44), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_45), .B(n_105), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_46), .B(n_105), .Y(n_161) );
AO22x2_ASAP7_75t_L g432 ( .A1(n_47), .A2(n_68), .B1(n_433), .B2(n_434), .Y(n_432) );
INVxp67_ASAP7_75t_L g531 ( .A(n_47), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_48), .A2(n_417), .B1(n_420), .B2(n_421), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_48), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_50), .Y(n_483) );
INVx1_ASAP7_75t_L g121 ( .A(n_51), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_52), .B(n_105), .Y(n_116) );
INVx1_ASAP7_75t_L g95 ( .A(n_53), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_54), .Y(n_528) );
AO32x2_ASAP7_75t_L g150 ( .A1(n_55), .A2(n_125), .A3(n_144), .B1(n_151), .B2(n_156), .Y(n_150) );
INVx1_ASAP7_75t_L g140 ( .A(n_56), .Y(n_140) );
INVx1_ASAP7_75t_L g182 ( .A(n_57), .Y(n_182) );
AO22x2_ASAP7_75t_L g437 ( .A1(n_58), .A2(n_74), .B1(n_433), .B2(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_59), .B(n_101), .Y(n_183) );
AOI22xp5_ASAP7_75t_SL g537 ( .A1(n_59), .A2(n_424), .B1(n_523), .B2(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_59), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_62), .Y(n_450) );
INVx1_ASAP7_75t_L g412 ( .A(n_64), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_65), .B(n_153), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_66), .B(n_101), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_67), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_69), .Y(n_510) );
INVx2_ASAP7_75t_L g93 ( .A(n_70), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_71), .B(n_101), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_73), .A2(n_77), .B1(n_101), .B2(n_102), .Y(n_196) );
INVx1_ASAP7_75t_L g433 ( .A(n_75), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_75), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_76), .B(n_101), .Y(n_138) );
INVx1_ASAP7_75t_L g419 ( .A(n_76), .Y(n_419) );
AOI221xp5_ASAP7_75t_SL g78 ( .A1(n_79), .A2(n_401), .B1(n_407), .B2(n_524), .C(n_536), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_80), .Y(n_79) );
AND2x2_ASAP7_75t_SL g80 ( .A(n_81), .B(n_367), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_271), .C(n_355), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_214), .C(n_236), .D(n_252), .Y(n_82) );
AOI221xp5_ASAP7_75t_L g83 ( .A1(n_84), .A2(n_147), .B1(n_173), .B2(n_192), .C(n_200), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_86), .B(n_123), .Y(n_85) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_86), .B(n_192), .Y(n_226) );
NAND4xp25_ASAP7_75t_L g266 ( .A(n_86), .B(n_254), .C(n_267), .D(n_269), .Y(n_266) );
INVxp67_ASAP7_75t_L g383 ( .A(n_86), .Y(n_383) );
INVx3_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
OR2x2_ASAP7_75t_L g265 ( .A(n_87), .B(n_203), .Y(n_265) );
AND2x2_ASAP7_75t_L g289 ( .A(n_87), .B(n_123), .Y(n_289) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g256 ( .A(n_88), .B(n_191), .Y(n_256) );
AND2x2_ASAP7_75t_L g296 ( .A(n_88), .B(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_L g313 ( .A(n_88), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_88), .B(n_124), .Y(n_337) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g190 ( .A(n_89), .B(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g208 ( .A(n_89), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g220 ( .A(n_89), .B(n_124), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_89), .B(n_134), .Y(n_242) );
OA21x2_ASAP7_75t_L g89 ( .A1(n_90), .A2(n_97), .B(n_122), .Y(n_89) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_90), .A2(n_135), .B(n_145), .Y(n_134) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_92), .Y(n_125) );
AND2x2_ASAP7_75t_L g92 ( .A(n_93), .B(n_94), .Y(n_92) );
AND2x2_ASAP7_75t_SL g146 ( .A(n_93), .B(n_94), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g94 ( .A(n_95), .B(n_96), .Y(n_94) );
OAI21xp5_ASAP7_75t_L g97 ( .A1(n_98), .A2(n_111), .B(n_120), .Y(n_97) );
O2A1O1Ixp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_100), .B(n_104), .C(n_107), .Y(n_98) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx2_ASAP7_75t_L g106 ( .A(n_103), .Y(n_106) );
INVx1_ASAP7_75t_L g114 ( .A(n_103), .Y(n_114) );
INVx3_ASAP7_75t_L g181 ( .A(n_105), .Y(n_181) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
BUFx3_ASAP7_75t_L g154 ( .A(n_106), .Y(n_154) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_108), .A2(n_185), .B(n_186), .Y(n_184) );
INVx4_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx3_ASAP7_75t_L g119 ( .A(n_110), .Y(n_119) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_110), .Y(n_143) );
INVx1_ASAP7_75t_L g164 ( .A(n_110), .Y(n_164) );
AND2x2_ASAP7_75t_L g406 ( .A(n_110), .B(n_114), .Y(n_406) );
O2A1O1Ixp33_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_115), .B(n_116), .C(n_117), .Y(n_111) );
O2A1O1Ixp5_ASAP7_75t_L g139 ( .A1(n_112), .A2(n_140), .B(n_141), .C(n_142), .Y(n_139) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_117), .A2(n_131), .B(n_132), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_117), .A2(n_143), .B1(n_171), .B2(n_172), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_117), .A2(n_143), .B1(n_196), .B2(n_197), .Y(n_195) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g127 ( .A1(n_118), .A2(n_128), .B(n_129), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_118), .A2(n_137), .B(n_138), .Y(n_136) );
O2A1O1Ixp5_ASAP7_75t_SL g180 ( .A1(n_118), .A2(n_181), .B(n_182), .C(n_183), .Y(n_180) );
INVx5_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g151 ( .A1(n_119), .A2(n_143), .B1(n_152), .B2(n_155), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g126 ( .A1(n_120), .A2(n_127), .B(n_130), .Y(n_126) );
BUFx3_ASAP7_75t_L g144 ( .A(n_120), .Y(n_144) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_120), .A2(n_160), .B(n_165), .Y(n_159) );
OAI21xp5_ASAP7_75t_L g179 ( .A1(n_120), .A2(n_180), .B(n_184), .Y(n_179) );
AND2x4_ASAP7_75t_L g405 ( .A(n_120), .B(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_121), .Y(n_533) );
AND2x2_ASAP7_75t_L g223 ( .A(n_123), .B(n_224), .Y(n_223) );
AOI221xp5_ASAP7_75t_L g272 ( .A1(n_123), .A2(n_273), .B1(n_276), .B2(n_278), .C(n_282), .Y(n_272) );
AND2x2_ASAP7_75t_L g331 ( .A(n_123), .B(n_296), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_123), .B(n_313), .Y(n_365) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_134), .Y(n_123) );
INVx3_ASAP7_75t_L g191 ( .A(n_124), .Y(n_191) );
AND2x2_ASAP7_75t_L g240 ( .A(n_124), .B(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g294 ( .A(n_124), .B(n_209), .Y(n_294) );
AND2x2_ASAP7_75t_L g352 ( .A(n_124), .B(n_353), .Y(n_352) );
OA21x2_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B(n_133), .Y(n_124) );
INVx4_ASAP7_75t_L g194 ( .A(n_125), .Y(n_194) );
AND2x2_ASAP7_75t_L g192 ( .A(n_134), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g209 ( .A(n_134), .Y(n_209) );
INVx1_ASAP7_75t_L g264 ( .A(n_134), .Y(n_264) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_134), .Y(n_270) );
AND2x2_ASAP7_75t_L g315 ( .A(n_134), .B(n_191), .Y(n_315) );
OR2x2_ASAP7_75t_L g354 ( .A(n_134), .B(n_193), .Y(n_354) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_139), .B(n_144), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_142), .A2(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND3xp33_ASAP7_75t_L g213 ( .A(n_144), .B(n_194), .C(n_195), .Y(n_213) );
INVx2_ASAP7_75t_L g156 ( .A(n_146), .Y(n_156) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_146), .A2(n_159), .B(n_168), .Y(n_158) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_146), .A2(n_179), .B(n_187), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_147), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_157), .Y(n_147) );
AND2x2_ASAP7_75t_L g350 ( .A(n_148), .B(n_347), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_148), .B(n_332), .Y(n_382) );
BUFx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g281 ( .A(n_149), .B(n_205), .Y(n_281) );
AND2x2_ASAP7_75t_L g330 ( .A(n_149), .B(n_176), .Y(n_330) );
INVx1_ASAP7_75t_L g376 ( .A(n_149), .Y(n_376) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_150), .Y(n_189) );
AND2x2_ASAP7_75t_L g231 ( .A(n_150), .B(n_205), .Y(n_231) );
INVx1_ASAP7_75t_L g248 ( .A(n_150), .Y(n_248) );
AND2x2_ASAP7_75t_L g254 ( .A(n_150), .B(n_169), .Y(n_254) );
AND2x2_ASAP7_75t_L g322 ( .A(n_157), .B(n_230), .Y(n_322) );
INVx2_ASAP7_75t_L g387 ( .A(n_157), .Y(n_387) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_169), .Y(n_157) );
AND2x2_ASAP7_75t_L g204 ( .A(n_158), .B(n_205), .Y(n_204) );
OR2x2_ASAP7_75t_L g217 ( .A(n_158), .B(n_177), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_158), .B(n_176), .Y(n_245) );
INVx1_ASAP7_75t_L g251 ( .A(n_158), .Y(n_251) );
INVx1_ASAP7_75t_L g268 ( .A(n_158), .Y(n_268) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_158), .Y(n_280) );
INVx2_ASAP7_75t_L g348 ( .A(n_158), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g205 ( .A(n_169), .Y(n_205) );
BUFx2_ASAP7_75t_L g302 ( .A(n_169), .Y(n_302) );
AND2x2_ASAP7_75t_L g347 ( .A(n_169), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_188), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_175), .B(n_284), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_175), .A2(n_346), .B(n_360), .Y(n_370) );
AND2x2_ASAP7_75t_L g395 ( .A(n_175), .B(n_281), .Y(n_395) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx1_ASAP7_75t_L g317 ( .A(n_177), .Y(n_317) );
AND2x2_ASAP7_75t_L g346 ( .A(n_177), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_178), .Y(n_230) );
INVx2_ASAP7_75t_L g249 ( .A(n_178), .Y(n_249) );
OR2x2_ASAP7_75t_L g250 ( .A(n_178), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx2_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
OR2x2_ASAP7_75t_L g216 ( .A(n_189), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g284 ( .A(n_189), .B(n_280), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_189), .B(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g385 ( .A(n_189), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_189), .B(n_322), .Y(n_397) );
AND2x2_ASAP7_75t_L g276 ( .A(n_190), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g299 ( .A(n_190), .B(n_192), .Y(n_299) );
INVx2_ASAP7_75t_L g211 ( .A(n_191), .Y(n_211) );
AND2x2_ASAP7_75t_L g239 ( .A(n_191), .B(n_212), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_191), .B(n_264), .Y(n_320) );
AND2x2_ASAP7_75t_L g234 ( .A(n_192), .B(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g381 ( .A(n_192), .Y(n_381) );
AND2x2_ASAP7_75t_L g393 ( .A(n_192), .B(n_256), .Y(n_393) );
AND2x2_ASAP7_75t_L g219 ( .A(n_193), .B(n_209), .Y(n_219) );
INVx1_ASAP7_75t_L g314 ( .A(n_193), .Y(n_314) );
AO21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_198), .Y(n_193) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x4_ASAP7_75t_L g212 ( .A(n_199), .B(n_213), .Y(n_212) );
INVxp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_206), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_203), .B(n_250), .Y(n_259) );
OR2x2_ASAP7_75t_L g391 ( .A(n_203), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g308 ( .A(n_204), .B(n_249), .Y(n_308) );
AND2x2_ASAP7_75t_L g316 ( .A(n_204), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g375 ( .A(n_204), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g399 ( .A(n_204), .B(n_246), .Y(n_399) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_205), .B(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g386 ( .A(n_205), .B(n_249), .Y(n_386) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
AND2x2_ASAP7_75t_L g238 ( .A(n_208), .B(n_239), .Y(n_238) );
INVxp67_ASAP7_75t_L g400 ( .A(n_208), .Y(n_400) );
NOR2x1_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx1_ASAP7_75t_L g235 ( .A(n_211), .Y(n_235) );
AND2x2_ASAP7_75t_L g286 ( .A(n_211), .B(n_219), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_211), .B(n_354), .Y(n_380) );
INVx2_ASAP7_75t_L g225 ( .A(n_212), .Y(n_225) );
INVx3_ASAP7_75t_L g277 ( .A(n_212), .Y(n_277) );
OR2x2_ASAP7_75t_L g305 ( .A(n_212), .B(n_306), .Y(n_305) );
AOI311xp33_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_218), .A3(n_220), .B(n_221), .C(n_232), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_215), .A2(n_253), .B(n_255), .C(n_257), .Y(n_252) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_SL g237 ( .A(n_217), .Y(n_237) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g255 ( .A(n_219), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_219), .B(n_235), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_219), .B(n_220), .Y(n_388) );
AND2x2_ASAP7_75t_L g310 ( .A(n_220), .B(n_224), .Y(n_310) );
AOI21xp33_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_226), .B(n_227), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g368 ( .A(n_224), .B(n_256), .Y(n_368) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_225), .B(n_242), .Y(n_241) );
INVx1_ASAP7_75t_L g262 ( .A(n_225), .Y(n_262) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
AND2x2_ASAP7_75t_L g253 ( .A(n_229), .B(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g298 ( .A(n_231), .Y(n_298) );
AND2x4_ASAP7_75t_L g360 ( .A(n_231), .B(n_329), .Y(n_360) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AOI222xp33_ASAP7_75t_L g311 ( .A1(n_234), .A2(n_300), .B1(n_312), .B2(n_316), .C1(n_318), .C2(n_322), .Y(n_311) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .C(n_243), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_237), .B(n_281), .Y(n_304) );
INVx1_ASAP7_75t_L g326 ( .A(n_239), .Y(n_326) );
INVx1_ASAP7_75t_L g260 ( .A(n_241), .Y(n_260) );
OR2x2_ASAP7_75t_L g325 ( .A(n_242), .B(n_326), .Y(n_325) );
OAI21xp33_ASAP7_75t_SL g243 ( .A1(n_244), .A2(n_246), .B(n_250), .Y(n_243) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_244), .B(n_262), .C(n_263), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_244), .A2(n_281), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_248), .Y(n_301) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_249), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g358 ( .A(n_249), .Y(n_358) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_249), .Y(n_374) );
INVx2_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_254), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g306 ( .A(n_256), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_260), .B1(n_261), .B2(n_265), .C(n_266), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_260), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g394 ( .A(n_260), .Y(n_394) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g275 ( .A(n_267), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_267), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g333 ( .A(n_267), .B(n_281), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_267), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g366 ( .A(n_267), .B(n_301), .Y(n_366) );
BUFx3_ASAP7_75t_L g329 ( .A(n_268), .Y(n_329) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND5xp2_ASAP7_75t_L g271 ( .A(n_272), .B(n_290), .C(n_311), .D(n_323), .E(n_338), .Y(n_271) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI32xp33_ASAP7_75t_L g363 ( .A1(n_275), .A2(n_302), .A3(n_318), .B1(n_364), .B2(n_366), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_277), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_SL g287 ( .A(n_281), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_285), .B1(n_287), .B2(n_288), .Y(n_282) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_299), .B2(n_300), .C(n_303), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g362 ( .A(n_294), .B(n_313), .Y(n_362) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_299), .A2(n_360), .B1(n_378), .B2(n_383), .C(n_384), .Y(n_377) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx2_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_304), .A2(n_305), .B1(n_307), .B2(n_309), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g321 ( .A(n_313), .Y(n_321) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B1(n_331), .B2(n_332), .C1(n_333), .C2(n_334), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_332), .A2(n_379), .B1(n_381), .B2(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B(n_344), .Y(n_338) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_349), .B(n_351), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B(n_361), .C(n_363), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI211xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_371), .C(n_396), .Y(n_367) );
CKINVDCx16_ASAP7_75t_R g372 ( .A(n_368), .Y(n_372) );
INVxp67_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI211xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B(n_377), .C(n_389), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_388), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_393), .B1(n_394), .B2(n_395), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_402), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_403), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_406), .A2(n_532), .B(n_545), .Y(n_544) );
XNOR2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_423), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_413), .B2(n_414), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_416), .Y(n_422) );
INVx1_ASAP7_75t_L g421 ( .A(n_417), .Y(n_421) );
INVx2_ASAP7_75t_L g523 ( .A(n_424), .Y(n_523) );
AND2x2_ASAP7_75t_SL g424 ( .A(n_425), .B(n_481), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_461), .Y(n_425) );
OAI221xp5_ASAP7_75t_SL g426 ( .A1(n_427), .A2(n_444), .B1(n_445), .B2(n_450), .C(n_451), .Y(n_426) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_439), .Y(n_429) );
AND2x6_ASAP7_75t_L g454 ( .A(n_430), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_L g464 ( .A(n_430), .B(n_465), .Y(n_464) );
AND2x6_ASAP7_75t_L g494 ( .A(n_430), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_436), .Y(n_430) );
AND2x2_ASAP7_75t_L g449 ( .A(n_431), .B(n_437), .Y(n_449) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_432), .B(n_437), .Y(n_460) );
AND2x2_ASAP7_75t_L g470 ( .A(n_432), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g502 ( .A(n_432), .B(n_441), .Y(n_502) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_435), .Y(n_438) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g471 ( .A(n_437), .Y(n_471) );
INVx1_ASAP7_75t_L g501 ( .A(n_437), .Y(n_501) );
AND2x4_ASAP7_75t_L g448 ( .A(n_439), .B(n_449), .Y(n_448) );
AND2x4_ASAP7_75t_L g458 ( .A(n_439), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_439), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_442), .Y(n_439) );
OR2x2_ASAP7_75t_L g456 ( .A(n_440), .B(n_443), .Y(n_456) );
AND2x2_ASAP7_75t_L g465 ( .A(n_440), .B(n_443), .Y(n_465) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g495 ( .A(n_441), .B(n_443), .Y(n_495) );
AND2x2_ASAP7_75t_L g500 ( .A(n_442), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g514 ( .A(n_442), .Y(n_514) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g487 ( .A(n_449), .Y(n_487) );
NAND2x1p5_ASAP7_75t_L g491 ( .A(n_449), .B(n_465), .Y(n_491) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx11_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g486 ( .A(n_456), .B(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x6_ASAP7_75t_L g479 ( .A(n_460), .B(n_480), .Y(n_479) );
OAI221xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_466), .B1(n_467), .B2(n_472), .C(n_473), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx3_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g477 ( .A(n_465), .B(n_470), .Y(n_477) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g521 ( .A(n_471), .Y(n_521) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx8_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .C(n_509), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_488), .B2(n_489), .Y(n_482) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_496), .B1(n_497), .B2(n_503), .C(n_504), .Y(n_492) );
INVx2_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g519 ( .A(n_495), .Y(n_519) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx4f_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g508 ( .A(n_501), .Y(n_508) );
AND2x4_ASAP7_75t_L g507 ( .A(n_502), .B(n_508), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g513 ( .A(n_502), .B(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_515), .B2(n_516), .Y(n_509) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
AND3x1_ASAP7_75t_SL g526 ( .A(n_527), .B(n_532), .C(n_534), .Y(n_526) );
INVxp67_ASAP7_75t_L g540 ( .A(n_527), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g541 ( .A(n_532), .Y(n_541) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_533), .B(n_535), .Y(n_545) );
OR2x2_ASAP7_75t_SL g551 ( .A(n_534), .B(n_541), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
OAI322xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_539), .A3(n_541), .B1(n_542), .B2(n_546), .C1(n_547), .C2(n_549), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_543), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_551), .Y(n_550) );
endmodule