module fake_jpeg_30388_n_185 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_185);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_16),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_3),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_11),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_41),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_0),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_0),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_86),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_74),
.B(n_1),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_1),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_56),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_68),
.B1(n_54),
.B2(n_57),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_102),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_65),
.B1(n_68),
.B2(n_54),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_57),
.B1(n_77),
.B2(n_58),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_80),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_111),
.B(n_6),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_57),
.B1(n_84),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_107),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_97),
.A2(n_75),
.B1(n_71),
.B2(n_55),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_115),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_65),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_69),
.B1(n_67),
.B2(n_66),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_121),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_118),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_61),
.B1(n_60),
.B2(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_2),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_2),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_5),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_113),
.A2(n_70),
.B1(n_24),
.B2(n_25),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_132),
.B1(n_143),
.B2(n_21),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_70),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_13),
.C(n_14),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_3),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_134),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_12),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_7),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_141),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_32),
.A3(n_52),
.B1(n_51),
.B2(n_49),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_15),
.Y(n_154)
);

INVxp67_ASAP7_75t_SL g140 ( 
.A(n_107),
.Y(n_140)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_8),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_104),
.B(n_12),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_20),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_155),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_150),
.B1(n_40),
.B2(n_42),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_124),
.Y(n_149)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_133),
.B(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_157),
.C(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_34),
.C(n_35),
.D(n_38),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_136),
.C(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_22),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_26),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

OAI321xp33_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_46),
.A3(n_48),
.B1(n_53),
.B2(n_145),
.C(n_150),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_172),
.A2(n_147),
.B1(n_161),
.B2(n_157),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_174),
.B(n_175),
.C(n_163),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_164),
.C(n_151),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_179),
.B(n_176),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_169),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_165),
.C(n_166),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_182),
.A2(n_170),
.B(n_178),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_175),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_161),
.Y(n_185)
);


endmodule