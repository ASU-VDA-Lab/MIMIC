module fake_jpeg_10017_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx11_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_41),
.Y(n_45)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_52),
.Y(n_72)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_33),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_21),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_71),
.B(n_80),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_30),
.B(n_33),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_81),
.B(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_66),
.B(n_85),
.Y(n_106)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_70),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_21),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_34),
.B1(n_26),
.B2(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_73),
.A2(n_75),
.B1(n_89),
.B2(n_38),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_26),
.B1(n_41),
.B2(n_38),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_85),
.B1(n_25),
.B2(n_33),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_79),
.B(n_82),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_21),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_25),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_86),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_29),
.B(n_31),
.C(n_28),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_87),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_31),
.B1(n_29),
.B2(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_50),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_95),
.A2(n_118),
.B1(n_74),
.B2(n_32),
.Y(n_133)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_104),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_68),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_97),
.B(n_99),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_18),
.B(n_32),
.Y(n_135)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_100),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_30),
.B1(n_23),
.B2(n_28),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_88),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_67),
.B1(n_74),
.B2(n_78),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_16),
.B1(n_20),
.B2(n_22),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_64),
.B(n_63),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_81),
.Y(n_130)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_66),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_133),
.B1(n_117),
.B2(n_120),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_18),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_121),
.C(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_104),
.C(n_16),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_64),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_128),
.B(n_131),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_71),
.B(n_80),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_130),
.B(n_152),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_72),
.B(n_81),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_92),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_59),
.B1(n_73),
.B2(n_91),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_134),
.B1(n_136),
.B2(n_117),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_116),
.A2(n_76),
.B1(n_90),
.B2(n_37),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_135),
.A2(n_17),
.B(n_16),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_42),
.B1(n_37),
.B2(n_40),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_113),
.A2(n_19),
.B(n_24),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_139),
.A2(n_146),
.B(n_148),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_98),
.A2(n_42),
.B1(n_87),
.B2(n_40),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_145),
.B1(n_112),
.B2(n_94),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_96),
.A2(n_42),
.B1(n_40),
.B2(n_93),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_0),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_22),
.B(n_24),
.C(n_19),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_110),
.A2(n_24),
.B(n_19),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_105),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_169),
.C(n_177),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_147),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_156),
.B(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_111),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_159),
.Y(n_199)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_182),
.B(n_1),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_146),
.B(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_161),
.B(n_163),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_99),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_167),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_0),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_184),
.B(n_1),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_138),
.B(n_94),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_171),
.Y(n_215)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_176),
.B(n_149),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_100),
.B1(n_117),
.B2(n_107),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_148),
.B1(n_20),
.B2(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_16),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_129),
.A2(n_22),
.B1(n_20),
.B2(n_16),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_20),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_183),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_149),
.B(n_107),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_130),
.A2(n_24),
.B(n_19),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_183),
.A2(n_186),
.B1(n_148),
.B2(n_20),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_129),
.A2(n_24),
.B(n_19),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_139),
.C(n_152),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_148),
.C(n_20),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_134),
.A2(n_107),
.B1(n_24),
.B2(n_19),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_131),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_204),
.C(n_182),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_189),
.A2(n_191),
.B1(n_193),
.B2(n_197),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_141),
.B1(n_150),
.B2(n_123),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_195),
.A2(n_211),
.B(n_213),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_126),
.B(n_144),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_196),
.A2(n_202),
.B(n_210),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_150),
.B1(n_126),
.B2(n_148),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_203),
.B1(n_158),
.B2(n_176),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_164),
.B(n_185),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_207),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_153),
.B(n_8),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_172),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_221),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_239),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_187),
.A2(n_186),
.B1(n_155),
.B2(n_156),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_219),
.A2(n_227),
.B1(n_234),
.B2(n_203),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_169),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_224),
.C(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_192),
.Y(n_226)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_153),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_211),
.B(n_206),
.Y(n_257)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_187),
.A2(n_184),
.B1(n_168),
.B2(n_2),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_9),
.B(n_4),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_210),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_9),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_209),
.C(n_189),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_202),
.B(n_8),
.Y(n_239)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_205),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_198),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_190),
.B1(n_195),
.B2(n_214),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_247),
.A2(n_194),
.B1(n_2),
.B2(n_5),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_220),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_251),
.B(n_256),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_190),
.C(n_197),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_233),
.C(n_239),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_205),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_259),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_222),
.B(n_207),
.Y(n_262)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_262),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.C(n_271),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_241),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_267),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_238),
.C(n_217),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_214),
.B1(n_234),
.B2(n_215),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_269),
.B1(n_270),
.B2(n_245),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_229),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_256),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_2),
.C(n_4),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_2),
.C(n_5),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_265),
.C(n_267),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_5),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_242),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_244),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_279),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_247),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_281),
.B1(n_6),
.B2(n_11),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_249),
.B1(n_240),
.B2(n_253),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_287),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_258),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_285),
.B(n_289),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_257),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_6),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_255),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_246),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_272),
.C(n_7),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_283),
.A2(n_273),
.B(n_264),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_290),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_295),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_296),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_6),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_11),
.C(n_12),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_12),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_291),
.B1(n_292),
.B2(n_294),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_284),
.B1(n_289),
.B2(n_278),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_304),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_284),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_305),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_15),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_300),
.C(n_303),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_310),
.B(n_311),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_300),
.B(n_15),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_305),
.B(n_302),
.Y(n_314)
);

OAI31xp33_ASAP7_75t_SL g316 ( 
.A1(n_314),
.A2(n_312),
.A3(n_309),
.B(n_306),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_303),
.C(n_315),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_308),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);


endmodule