module fake_netlist_5_1414_n_778 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_778);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_778;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_696;
wire n_255;
wire n_550;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_113),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_88),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_62),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_6),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_3),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_82),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_33),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_65),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_42),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_109),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_99),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_59),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_29),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_103),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_125),
.Y(n_180)
);

NOR2xp67_ASAP7_75t_L g181 ( 
.A(n_70),
.B(n_120),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_30),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_93),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_101),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_107),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_40),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_25),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_63),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_52),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_57),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_3),
.B(n_1),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_124),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_127),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_13),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_20),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_68),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_138),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_75),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_193),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_0),
.B(n_2),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_23),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_4),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_26),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_8),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_162),
.B(n_9),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_213),
.Y(n_241)
);

OA21x2_ASAP7_75t_L g242 ( 
.A1(n_178),
.A2(n_9),
.B(n_10),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_186),
.B(n_10),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_192),
.B(n_195),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_173),
.Y(n_250)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_158),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_204),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_159),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_163),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_158),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_215),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_237),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_166),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_253),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_218),
.Y(n_267)
);

AND2x6_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_200),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_210),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_167),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_210),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_251),
.B(n_168),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_169),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_228),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_225),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g281 ( 
.A1(n_219),
.A2(n_208),
.B1(n_207),
.B2(n_163),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_227),
.B(n_170),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_171),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_222),
.B(n_176),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_225),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

AND2x6_ASAP7_75t_L g289 ( 
.A(n_222),
.B(n_181),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

BUFx6f_ASAP7_75t_SL g291 ( 
.A(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_231),
.Y(n_292)
);

CKINVDCx6p67_ASAP7_75t_R g293 ( 
.A(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_234),
.B(n_177),
.Y(n_294)
);

OR2x6_ASAP7_75t_L g295 ( 
.A(n_256),
.B(n_187),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_250),
.B(n_179),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_237),
.Y(n_297)
);

AO21x2_ASAP7_75t_L g298 ( 
.A1(n_220),
.A2(n_182),
.B(n_205),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_224),
.B(n_183),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_231),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_221),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_250),
.B(n_189),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_224),
.B(n_196),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_221),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_260),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_246),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_246),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_266),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_260),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_236),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_244),
.C(n_238),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_222),
.Y(n_315)
);

NOR3xp33_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_233),
.C(n_254),
.Y(n_316)
);

NAND2xp33_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_199),
.Y(n_317)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_257),
.B(n_228),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

O2A1O1Ixp5_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_246),
.B(n_228),
.C(n_248),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_271),
.B(n_228),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_246),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_293),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_259),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_294),
.B(n_235),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_257),
.B(n_235),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_269),
.B(n_240),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_262),
.B(n_297),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_254),
.C(n_207),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_262),
.B(n_202),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_270),
.A2(n_248),
.B(n_249),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_297),
.B(n_203),
.Y(n_332)
);

NOR2x1p5_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_208),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_265),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_240),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_272),
.A2(n_217),
.B1(n_243),
.B2(n_249),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_259),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_268),
.B(n_283),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_243),
.Y(n_339)
);

OR2x6_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_220),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_232),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g342 ( 
.A1(n_296),
.A2(n_217),
.B(n_303),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_273),
.B(n_252),
.Y(n_343)
);

O2A1O1Ixp33_ASAP7_75t_L g344 ( 
.A1(n_285),
.A2(n_230),
.B(n_229),
.C(n_226),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_299),
.B(n_252),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_265),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_261),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_268),
.B(n_232),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_241),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_264),
.Y(n_352)
);

BUFx6f_ASAP7_75t_SL g353 ( 
.A(n_295),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_288),
.B(n_214),
.Y(n_354)
);

A2O1A1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_230),
.B(n_229),
.C(n_226),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g356 ( 
.A1(n_295),
.A2(n_242),
.B1(n_214),
.B2(n_216),
.Y(n_356)
);

OAI21x1_ASAP7_75t_L g357 ( 
.A1(n_264),
.A2(n_221),
.B(n_242),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_267),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_268),
.A2(n_242),
.B1(n_245),
.B2(n_239),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

OAI22xp33_ASAP7_75t_L g362 ( 
.A1(n_295),
.A2(n_242),
.B1(n_216),
.B2(n_245),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_275),
.B(n_252),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_268),
.B(n_232),
.Y(n_366)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_291),
.B(n_232),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_288),
.B(n_232),
.Y(n_369)
);

O2A1O1Ixp5_ASAP7_75t_L g370 ( 
.A1(n_275),
.A2(n_245),
.B(n_239),
.C(n_84),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_287),
.B(n_282),
.Y(n_371)
);

O2A1O1Ixp5_ASAP7_75t_L g372 ( 
.A1(n_320),
.A2(n_277),
.B(n_279),
.C(n_280),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_321),
.A2(n_291),
.B1(n_277),
.B2(n_280),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g375 ( 
.A1(n_312),
.A2(n_301),
.B(n_290),
.C(n_287),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_349),
.A2(n_282),
.B(n_279),
.Y(n_376)
);

O2A1O1Ixp33_ASAP7_75t_L g377 ( 
.A1(n_326),
.A2(n_301),
.B(n_290),
.C(n_298),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_305),
.B(n_302),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_366),
.A2(n_305),
.B(n_302),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_315),
.A2(n_298),
.B(n_245),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_340),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_352),
.Y(n_383)
);

AND2x6_ASAP7_75t_L g384 ( 
.A(n_307),
.B(n_298),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_239),
.Y(n_386)
);

NOR2xp67_ASAP7_75t_L g387 ( 
.A(n_308),
.B(n_27),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_339),
.A2(n_245),
.B(n_239),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_239),
.B1(n_83),
.B2(n_85),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_322),
.B(n_28),
.Y(n_390)
);

BUFx4f_ASAP7_75t_L g391 ( 
.A(n_340),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_323),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_327),
.B(n_11),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_360),
.A2(n_80),
.B(n_155),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_342),
.B(n_11),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_308),
.A2(n_89),
.B(n_153),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_310),
.A2(n_335),
.B1(n_309),
.B2(n_325),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_310),
.A2(n_309),
.B(n_359),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_317),
.A2(n_79),
.B(n_152),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_368),
.A2(n_77),
.B(n_151),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_331),
.A2(n_369),
.B(n_346),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_319),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_330),
.B(n_12),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_365),
.Y(n_405)
);

NAND2x1p5_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_31),
.Y(n_406)
);

AOI21xp33_ASAP7_75t_L g407 ( 
.A1(n_356),
.A2(n_12),
.B(n_13),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_332),
.B(n_345),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_L g409 ( 
.A1(n_313),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_306),
.Y(n_410)
);

O2A1O1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_362),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_369),
.A2(n_94),
.B(n_150),
.Y(n_412)
);

AO21x1_ASAP7_75t_L g413 ( 
.A1(n_336),
.A2(n_17),
.B(n_18),
.Y(n_413)
);

O2A1O1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_336),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

NAND2x1p5_ASAP7_75t_L g416 ( 
.A(n_351),
.B(n_32),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_311),
.A2(n_95),
.B(n_148),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_329),
.B(n_334),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_350),
.A2(n_91),
.B1(n_146),
.B2(n_145),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_361),
.B(n_19),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

O2A1O1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_355),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_318),
.B(n_34),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_363),
.B(n_21),
.Y(n_424)
);

AOI21x1_ASAP7_75t_L g425 ( 
.A1(n_358),
.A2(n_97),
.B(n_35),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_357),
.A2(n_98),
.B(n_36),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_316),
.A2(n_22),
.B(n_37),
.C(n_38),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_318),
.B(n_39),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_324),
.Y(n_430)
);

CKINVDCx8_ASAP7_75t_R g431 ( 
.A(n_353),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_324),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_318),
.A2(n_45),
.B(n_47),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_348),
.A2(n_48),
.B(n_49),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

AO32x2_ASAP7_75t_L g436 ( 
.A1(n_318),
.A2(n_50),
.A3(n_51),
.B1(n_53),
.B2(n_54),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_348),
.B(n_55),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_370),
.A2(n_56),
.B(n_58),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_353),
.B(n_60),
.Y(n_439)
);

AO22x1_ASAP7_75t_L g440 ( 
.A1(n_333),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_398),
.B(n_367),
.Y(n_441)
);

NAND3xp33_ASAP7_75t_SL g442 ( 
.A(n_404),
.B(n_344),
.C(n_72),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_392),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_372),
.A2(n_376),
.B(n_402),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_371),
.A2(n_367),
.B(n_73),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_399),
.A2(n_367),
.B(n_74),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_395),
.B(n_367),
.Y(n_447)
);

AO31x2_ASAP7_75t_L g448 ( 
.A1(n_380),
.A2(n_367),
.A3(n_76),
.B(n_90),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_378),
.A2(n_390),
.B(n_423),
.Y(n_449)
);

AOI21x1_ASAP7_75t_L g450 ( 
.A1(n_379),
.A2(n_367),
.B(n_96),
.Y(n_450)
);

NAND3x1_ASAP7_75t_L g451 ( 
.A(n_408),
.B(n_69),
.C(n_100),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_425),
.A2(n_102),
.B(n_104),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_105),
.B(n_108),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_382),
.B(n_110),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_418),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_373),
.B(n_115),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_405),
.B(n_116),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_374),
.A2(n_117),
.B(n_118),
.Y(n_459)
);

AO31x2_ASAP7_75t_L g460 ( 
.A1(n_375),
.A2(n_119),
.A3(n_121),
.B(n_122),
.Y(n_460)
);

OA22x2_ASAP7_75t_L g461 ( 
.A1(n_381),
.A2(n_123),
.B1(n_128),
.B2(n_130),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_383),
.A2(n_131),
.B(n_132),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_396),
.B(n_394),
.Y(n_464)
);

CKINVDCx11_ASAP7_75t_R g465 ( 
.A(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_384),
.B(n_134),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_384),
.B(n_135),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_136),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_391),
.B(n_137),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_430),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_433),
.A2(n_427),
.B(n_397),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_377),
.A2(n_407),
.B(n_411),
.C(n_387),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_393),
.B(n_386),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_391),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_383),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_387),
.A2(n_140),
.B(n_143),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_439),
.B(n_406),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_416),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_384),
.A2(n_388),
.B(n_400),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_420),
.B(n_144),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_424),
.B(n_426),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_426),
.B(n_157),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_435),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

NOR3xp33_ASAP7_75t_L g488 ( 
.A(n_440),
.B(n_414),
.C(n_409),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_438),
.A2(n_434),
.B(n_401),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_428),
.A2(n_389),
.B(n_437),
.Y(n_490)
);

NOR2x1_ASAP7_75t_SL g491 ( 
.A(n_432),
.B(n_419),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_413),
.B(n_417),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_412),
.B(n_422),
.Y(n_493)
);

NAND2x1_ASAP7_75t_L g494 ( 
.A(n_436),
.B(n_383),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_436),
.B(n_418),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_436),
.A2(n_396),
.B(n_312),
.C(n_395),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_392),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_382),
.B(n_405),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_496),
.B(n_464),
.Y(n_499)
);

NAND2x1p5_ASAP7_75t_L g500 ( 
.A(n_477),
.B(n_472),
.Y(n_500)
);

AO21x1_ASAP7_75t_L g501 ( 
.A1(n_495),
.A2(n_490),
.B(n_492),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_498),
.B(n_455),
.Y(n_502)
);

OAI21x1_ASAP7_75t_L g503 ( 
.A1(n_444),
.A2(n_489),
.B(n_445),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_498),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_458),
.B(n_457),
.Y(n_506)
);

AOI221xp5_ASAP7_75t_L g507 ( 
.A1(n_488),
.A2(n_483),
.B1(n_474),
.B2(n_480),
.C(n_458),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_461),
.A2(n_490),
.B1(n_442),
.B2(n_492),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_SL g509 ( 
.A(n_481),
.B(n_466),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_462),
.Y(n_510)
);

BUFx2_ASAP7_75t_R g511 ( 
.A(n_497),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_443),
.B(n_461),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_475),
.A2(n_441),
.B(n_447),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_467),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_487),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_482),
.A2(n_450),
.B(n_446),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_447),
.A2(n_441),
.B1(n_494),
.B2(n_484),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_466),
.A2(n_469),
.B(n_470),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_476),
.B(n_468),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_465),
.Y(n_520)
);

AOI22x1_ASAP7_75t_L g521 ( 
.A1(n_449),
.A2(n_482),
.B1(n_486),
.B2(n_471),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_452),
.A2(n_485),
.B(n_459),
.Y(n_522)
);

OAI21x1_ASAP7_75t_SL g523 ( 
.A1(n_491),
.A2(n_469),
.B(n_470),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_493),
.A2(n_454),
.B(n_484),
.Y(n_524)
);

OA21x2_ASAP7_75t_L g525 ( 
.A1(n_493),
.A2(n_463),
.B(n_485),
.Y(n_525)
);

O2A1O1Ixp33_ASAP7_75t_SL g526 ( 
.A1(n_456),
.A2(n_479),
.B(n_453),
.C(n_451),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_448),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_448),
.A2(n_474),
.B(n_496),
.Y(n_529)
);

O2A1O1Ixp33_ASAP7_75t_SL g530 ( 
.A1(n_460),
.A2(n_496),
.B(n_495),
.C(n_428),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_460),
.B(n_455),
.Y(n_531)
);

O2A1O1Ixp33_ASAP7_75t_L g532 ( 
.A1(n_460),
.A2(n_496),
.B(n_409),
.C(n_495),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_464),
.B(n_498),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_464),
.B(n_312),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_464),
.A2(n_316),
.B(n_408),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_495),
.A2(n_407),
.B1(n_488),
.B2(n_461),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_496),
.B(n_312),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_444),
.A2(n_372),
.B(n_489),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_464),
.B(n_498),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_497),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

A2O1A1Ixp33_ASAP7_75t_L g542 ( 
.A1(n_496),
.A2(n_395),
.B(n_396),
.C(n_483),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_455),
.B(n_477),
.Y(n_543)
);

OAI22xp33_ASAP7_75t_SL g544 ( 
.A1(n_480),
.A2(n_439),
.B1(n_343),
.B2(n_345),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_455),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_521),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_535),
.Y(n_547)
);

INVxp33_ASAP7_75t_L g548 ( 
.A(n_533),
.Y(n_548)
);

OR2x6_ASAP7_75t_L g549 ( 
.A(n_518),
.B(n_523),
.Y(n_549)
);

AOI21x1_ASAP7_75t_SL g550 ( 
.A1(n_537),
.A2(n_531),
.B(n_499),
.Y(n_550)
);

BUFx2_ASAP7_75t_SL g551 ( 
.A(n_539),
.Y(n_551)
);

AO21x2_ASAP7_75t_L g552 ( 
.A1(n_542),
.A2(n_513),
.B(n_516),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_536),
.A2(n_508),
.B1(n_542),
.B2(n_512),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_505),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_514),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_528),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_536),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_531),
.Y(n_558)
);

AOI21x1_ASAP7_75t_L g559 ( 
.A1(n_524),
.A2(n_517),
.B(n_503),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_514),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_538),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_531),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_529),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g565 ( 
.A1(n_530),
.A2(n_501),
.B(n_527),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_504),
.Y(n_566)
);

AO21x2_ASAP7_75t_L g567 ( 
.A1(n_530),
.A2(n_532),
.B(n_522),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g568 ( 
.A1(n_526),
.A2(n_525),
.B(n_510),
.Y(n_568)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_525),
.A2(n_508),
.B(n_507),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_519),
.B(n_506),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_525),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_541),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_502),
.B(n_545),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_515),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_502),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_512),
.B(n_504),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_515),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_543),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_543),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_543),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_512),
.B(n_500),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_500),
.B(n_509),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_540),
.B(n_511),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_556),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_570),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_557),
.B(n_520),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_556),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_557),
.B(n_562),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_557),
.B(n_544),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_562),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_547),
.B(n_575),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_562),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_559),
.A2(n_546),
.B(n_569),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_554),
.B(n_576),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_554),
.B(n_576),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_563),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_558),
.Y(n_599)
);

OR2x2_ASAP7_75t_L g600 ( 
.A(n_552),
.B(n_553),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_558),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_563),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_566),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_555),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_568),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_553),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_555),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_576),
.B(n_575),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_566),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_560),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_573),
.B(n_548),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_560),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_578),
.Y(n_615)
);

BUFx2_ASAP7_75t_SL g616 ( 
.A(n_582),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_564),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_561),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_572),
.B(n_581),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_581),
.B(n_580),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_552),
.B(n_573),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_552),
.B(n_565),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_551),
.B(n_579),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_568),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_590),
.B(n_619),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_605),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_618),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_L g628 ( 
.A1(n_590),
.A2(n_551),
.B1(n_581),
.B2(n_582),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_593),
.B(n_549),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_619),
.B(n_565),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_592),
.B(n_582),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_609),
.B(n_565),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_598),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_621),
.B(n_565),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_601),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_609),
.B(n_569),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_618),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_569),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_568),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_621),
.B(n_571),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_596),
.B(n_568),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_596),
.B(n_567),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_620),
.B(n_567),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_589),
.B(n_583),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_601),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_598),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_589),
.B(n_583),
.Y(n_647)
);

BUFx3_ASAP7_75t_L g648 ( 
.A(n_611),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_602),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_620),
.B(n_593),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_593),
.B(n_591),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_567),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_610),
.B(n_600),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_600),
.B(n_571),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_610),
.B(n_567),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_654),
.B(n_607),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_654),
.B(n_607),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_629),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_653),
.B(n_636),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_653),
.B(n_610),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_633),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_648),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_R g663 ( 
.A(n_648),
.B(n_584),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_627),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_640),
.B(n_622),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_636),
.B(n_622),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_627),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_603),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_633),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_629),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_648),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_627),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_646),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_629),
.B(n_638),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_638),
.B(n_617),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_640),
.B(n_587),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_637),
.Y(n_678)
);

NAND2x1p5_ASAP7_75t_L g679 ( 
.A(n_626),
.B(n_605),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_625),
.B(n_630),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_650),
.B(n_611),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_649),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_629),
.B(n_616),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_630),
.B(n_617),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_661),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_677),
.B(n_632),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_662),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_680),
.B(n_643),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_SL g689 ( 
.A1(n_658),
.A2(n_628),
.B(n_584),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_668),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_680),
.B(n_659),
.Y(n_691)
);

OR2x2_ASAP7_75t_L g692 ( 
.A(n_656),
.B(n_634),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_659),
.B(n_643),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_656),
.B(n_634),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_683),
.A2(n_631),
.B1(n_586),
.B2(n_587),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_677),
.B(n_632),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_674),
.B(n_639),
.Y(n_697)
);

OAI31xp33_ASAP7_75t_L g698 ( 
.A1(n_679),
.A2(n_613),
.A3(n_584),
.B(n_579),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_661),
.Y(n_699)
);

AND3x2_ASAP7_75t_L g700 ( 
.A(n_671),
.B(n_645),
.C(n_635),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_674),
.B(n_635),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_674),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_673),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_673),
.Y(n_704)
);

OAI32xp33_ASAP7_75t_L g705 ( 
.A1(n_694),
.A2(n_657),
.A3(n_681),
.B1(n_665),
.B2(n_682),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_689),
.A2(n_683),
.B1(n_670),
.B2(n_658),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_698),
.B(n_663),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_697),
.B(n_674),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_697),
.B(n_666),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_695),
.A2(n_690),
.B1(n_683),
.B2(n_670),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_704),
.B(n_666),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_701),
.A2(n_683),
.B1(n_658),
.B2(n_670),
.Y(n_712)
);

O2A1O1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_687),
.A2(n_623),
.B(n_657),
.C(n_615),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_701),
.A2(n_702),
.B1(n_660),
.B2(n_616),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_685),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_699),
.A2(n_549),
.B(n_682),
.C(n_676),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_691),
.B(n_660),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_708),
.B(n_702),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_707),
.A2(n_694),
.B1(n_701),
.B2(n_692),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_711),
.B(n_686),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_SL g721 ( 
.A1(n_705),
.A2(n_691),
.B1(n_655),
.B2(n_642),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_715),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_709),
.B(n_688),
.Y(n_723)
);

AOI311xp33_ASAP7_75t_L g724 ( 
.A1(n_719),
.A2(n_711),
.A3(n_703),
.B(n_696),
.C(n_676),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_718),
.Y(n_725)
);

AOI221xp5_ASAP7_75t_L g726 ( 
.A1(n_721),
.A2(n_713),
.B1(n_716),
.B2(n_710),
.C(n_706),
.Y(n_726)
);

A2O1A1O1Ixp25_ASAP7_75t_L g727 ( 
.A1(n_721),
.A2(n_700),
.B(n_714),
.C(n_712),
.D(n_669),
.Y(n_727)
);

OAI221xp5_ASAP7_75t_SL g728 ( 
.A1(n_720),
.A2(n_665),
.B1(n_549),
.B2(n_717),
.C(n_688),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_722),
.A2(n_655),
.B1(n_642),
.B2(n_693),
.Y(n_729)
);

AND4x1_ASAP7_75t_L g730 ( 
.A(n_724),
.B(n_723),
.C(n_693),
.D(n_578),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_725),
.Y(n_731)
);

AND4x1_ASAP7_75t_L g732 ( 
.A(n_726),
.B(n_580),
.C(n_577),
.D(n_639),
.Y(n_732)
);

AOI211xp5_ASAP7_75t_L g733 ( 
.A1(n_727),
.A2(n_647),
.B(n_644),
.C(n_577),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_732),
.B(n_730),
.Y(n_734)
);

NOR2x1_ASAP7_75t_L g735 ( 
.A(n_731),
.B(n_728),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_734),
.A2(n_733),
.B1(n_729),
.B2(n_684),
.Y(n_736)
);

NOR2x1_ASAP7_75t_L g737 ( 
.A(n_735),
.B(n_608),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_734),
.A2(n_675),
.B1(n_684),
.B2(n_650),
.Y(n_738)
);

XOR2xp5_ASAP7_75t_L g739 ( 
.A(n_736),
.B(n_679),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_737),
.Y(n_740)
);

NAND3xp33_ASAP7_75t_L g741 ( 
.A(n_738),
.B(n_574),
.C(n_599),
.Y(n_741)
);

NAND2x1p5_ASAP7_75t_L g742 ( 
.A(n_737),
.B(n_574),
.Y(n_742)
);

NAND4xp75_ASAP7_75t_L g743 ( 
.A(n_737),
.B(n_614),
.C(n_612),
.D(n_675),
.Y(n_743)
);

NAND2xp33_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_679),
.Y(n_744)
);

XNOR2x1_ASAP7_75t_L g745 ( 
.A(n_737),
.B(n_549),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_742),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_739),
.A2(n_641),
.B1(n_645),
.B2(n_672),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_740),
.B(n_678),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_741),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_744),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_745),
.Y(n_751)
);

OR2x6_ASAP7_75t_L g752 ( 
.A(n_751),
.B(n_743),
.Y(n_752)
);

AO22x2_ASAP7_75t_L g753 ( 
.A1(n_749),
.A2(n_574),
.B1(n_604),
.B2(n_608),
.Y(n_753)
);

BUFx2_ASAP7_75t_SL g754 ( 
.A(n_746),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_748),
.Y(n_755)
);

AO22x2_ASAP7_75t_L g756 ( 
.A1(n_750),
.A2(n_604),
.B1(n_626),
.B2(n_597),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_752),
.A2(n_747),
.B1(n_647),
.B2(n_644),
.Y(n_757)
);

XNOR2xp5_ASAP7_75t_L g758 ( 
.A(n_754),
.B(n_549),
.Y(n_758)
);

OAI22x1_ASAP7_75t_L g759 ( 
.A1(n_755),
.A2(n_626),
.B1(n_605),
.B2(n_599),
.Y(n_759)
);

XOR2x2_ASAP7_75t_L g760 ( 
.A(n_756),
.B(n_614),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_753),
.A2(n_641),
.B1(n_549),
.B2(n_597),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_754),
.B(n_678),
.Y(n_762)
);

OA21x2_ASAP7_75t_L g763 ( 
.A1(n_755),
.A2(n_546),
.B(n_672),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_762),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_SL g765 ( 
.A1(n_758),
.A2(n_626),
.B1(n_612),
.B2(n_546),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_763),
.A2(n_550),
.B(n_559),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_757),
.A2(n_605),
.B1(n_664),
.B2(n_667),
.Y(n_767)
);

AO221x1_ASAP7_75t_L g768 ( 
.A1(n_759),
.A2(n_624),
.B1(n_606),
.B2(n_588),
.C(n_585),
.Y(n_768)
);

OAI21x1_ASAP7_75t_L g769 ( 
.A1(n_761),
.A2(n_550),
.B(n_667),
.Y(n_769)
);

OAI21xp33_ASAP7_75t_L g770 ( 
.A1(n_760),
.A2(n_652),
.B(n_664),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_770),
.A2(n_652),
.B1(n_594),
.B2(n_651),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_764),
.A2(n_594),
.B1(n_651),
.B2(n_585),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_768),
.Y(n_773)
);

OAI21xp33_ASAP7_75t_L g774 ( 
.A1(n_767),
.A2(n_769),
.B(n_766),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_773),
.B(n_765),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_774),
.Y(n_776)
);

OA21x2_ASAP7_75t_L g777 ( 
.A1(n_775),
.A2(n_771),
.B(n_772),
.Y(n_777)
);

AOI21xp33_ASAP7_75t_L g778 ( 
.A1(n_777),
.A2(n_776),
.B(n_594),
.Y(n_778)
);


endmodule