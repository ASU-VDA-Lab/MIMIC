module fake_jpeg_482_n_686 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_686);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_686;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_4),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_61),
.B(n_62),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_65),
.Y(n_179)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_67),
.B(n_76),
.Y(n_177)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_70),
.B(n_71),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_8),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_72),
.Y(n_203)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_74),
.Y(n_220)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_75),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_30),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g142 ( 
.A(n_77),
.Y(n_142)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_27),
.B(n_11),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_80),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_81),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_82),
.Y(n_225)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_84),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_85),
.B(n_94),
.Y(n_181)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_86),
.Y(n_169)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_20),
.Y(n_87)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_88),
.Y(n_195)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_90),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_91),
.Y(n_136)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g223 ( 
.A(n_92),
.Y(n_223)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_93),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_99),
.Y(n_193)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_100),
.Y(n_172)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_102),
.B(n_103),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_48),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_104),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_37),
.A2(n_11),
.B(n_18),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g186 ( 
.A1(n_105),
.A2(n_14),
.B(n_19),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_108),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_40),
.B(n_11),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_129),
.Y(n_199)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_11),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_52),
.Y(n_113)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_40),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_115),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_117),
.Y(n_214)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_118),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_120),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_29),
.Y(n_121)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_124),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx2_ASAP7_75t_SL g166 ( 
.A(n_126),
.Y(n_166)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_44),
.Y(n_127)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_127),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_44),
.B(n_13),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_32),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_48),
.Y(n_130)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_29),
.Y(n_132)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_60),
.A2(n_58),
.B1(n_25),
.B2(n_35),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_134),
.A2(n_147),
.B1(n_150),
.B2(n_154),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_143),
.B(n_159),
.C(n_188),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_87),
.A2(n_31),
.B1(n_25),
.B2(n_58),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_31),
.B1(n_35),
.B2(n_41),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_61),
.B(n_56),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_151),
.B(n_156),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_109),
.B(n_56),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_152),
.B(n_211),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_63),
.A2(n_31),
.B1(n_41),
.B2(n_45),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_59),
.B(n_45),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_54),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_75),
.A2(n_54),
.B1(n_21),
.B2(n_26),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_162),
.A2(n_198),
.B1(n_148),
.B2(n_161),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_110),
.B(n_21),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_171),
.B(n_191),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_73),
.A2(n_33),
.B1(n_28),
.B2(n_26),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_173),
.A2(n_175),
.B1(n_187),
.B2(n_197),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_98),
.A2(n_33),
.B1(n_28),
.B2(n_20),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_81),
.B(n_20),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_178),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_186),
.A2(n_213),
.B(n_175),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_116),
.A2(n_20),
.B1(n_53),
.B2(n_39),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_82),
.B(n_14),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_114),
.B(n_15),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_106),
.B1(n_95),
.B2(n_90),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_84),
.A2(n_20),
.B1(n_53),
.B2(n_39),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_101),
.A2(n_53),
.B1(n_7),
.B2(n_13),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_118),
.A2(n_53),
.B1(n_7),
.B2(n_16),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_207),
.A2(n_210),
.B1(n_213),
.B2(n_217),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_105),
.B(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_208),
.B(n_212),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_107),
.A2(n_66),
.B1(n_69),
.B2(n_96),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_78),
.B(n_6),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_108),
.B(n_6),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_77),
.A2(n_53),
.B1(n_7),
.B2(n_17),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_64),
.B(n_5),
.Y(n_215)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_215),
.B(n_216),
.C(n_230),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_65),
.B(n_5),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_72),
.A2(n_5),
.B1(n_18),
.B2(n_17),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_78),
.B(n_19),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_77),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_117),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_222),
.Y(n_297)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_130),
.Y(n_226)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_74),
.A2(n_125),
.B1(n_119),
.B2(n_111),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_229),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_91),
.B(n_5),
.Y(n_230)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_145),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_233),
.Y(n_343)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_225),
.Y(n_234)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_235),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_126),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_236),
.B(n_237),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_1),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_96),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_238),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_231),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_239),
.Y(n_323)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_241),
.Y(n_319)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_243),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_244),
.B(n_245),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_177),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_246),
.A2(n_250),
.B1(n_187),
.B2(n_197),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_189),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_248),
.B(n_284),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_170),
.B(n_1),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_249),
.B(n_260),
.Y(n_342)
);

AOI22x1_ASAP7_75t_L g250 ( 
.A1(n_188),
.A2(n_88),
.B1(n_115),
.B2(n_92),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_251),
.B(n_252),
.Y(n_335)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

BUFx4f_ASAP7_75t_SL g254 ( 
.A(n_165),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_254),
.Y(n_325)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_255),
.Y(n_346)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_185),
.Y(n_256)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_214),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_257),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_140),
.B(n_120),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_135),
.Y(n_259)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_259),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_141),
.B(n_2),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_172),
.Y(n_261)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_180),
.Y(n_262)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_262),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_263),
.A2(n_310),
.B1(n_316),
.B2(n_318),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_159),
.B(n_4),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_264),
.B(n_278),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_265),
.B(n_274),
.Y(n_345)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_163),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_267),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_268),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_219),
.A2(n_4),
.B1(n_17),
.B2(n_204),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_269),
.Y(n_337)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_190),
.Y(n_271)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_271),
.Y(n_349)
);

OR2x2_ASAP7_75t_SL g272 ( 
.A(n_178),
.B(n_17),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_272),
.B(n_312),
.C(n_313),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_4),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_273),
.Y(n_353)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_164),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_275),
.Y(n_354)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_135),
.Y(n_276)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_276),
.Y(n_366)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_139),
.Y(n_277)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_277),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_169),
.B(n_193),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_178),
.B(n_153),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g348 ( 
.A(n_279),
.B(n_287),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_281),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_139),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_282),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_283),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_181),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_176),
.B(n_146),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_286),
.B(n_309),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g287 ( 
.A(n_149),
.B(n_144),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_155),
.B(n_174),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_290),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_196),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_160),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_163),
.Y(n_291)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_291),
.Y(n_370)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_200),
.Y(n_292)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_293),
.B(n_295),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_157),
.B(n_192),
.Y(n_295)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_179),
.Y(n_296)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_296),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_206),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_301),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_218),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_183),
.A2(n_168),
.B1(n_202),
.B2(n_206),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_302),
.A2(n_305),
.B1(n_307),
.B2(n_308),
.Y(n_332)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_227),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_304),
.B(n_306),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_168),
.A2(n_202),
.B1(n_166),
.B2(n_165),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_142),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_161),
.B(n_182),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_195),
.Y(n_308)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_173),
.A2(n_134),
.B(n_147),
.C(n_201),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_218),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_136),
.B(n_138),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_227),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_136),
.B(n_138),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_314),
.B(n_315),
.C(n_317),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_142),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_167),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_167),
.B(n_224),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_224),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_294),
.A2(n_229),
.B1(n_154),
.B2(n_150),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_322),
.A2(n_327),
.B1(n_331),
.B2(n_356),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_303),
.A2(n_207),
.B1(n_220),
.B2(n_203),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_242),
.A2(n_223),
.B1(n_203),
.B2(n_220),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_336),
.A2(n_347),
.B1(n_361),
.B2(n_369),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_309),
.A2(n_223),
.B1(n_195),
.B2(n_205),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g352 ( 
.A1(n_283),
.A2(n_210),
.B(n_182),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_352),
.A2(n_360),
.B(n_377),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_246),
.A2(n_205),
.B1(n_184),
.B2(n_158),
.Y(n_356)
);

AOI32xp33_ASAP7_75t_L g358 ( 
.A1(n_236),
.A2(n_264),
.A3(n_266),
.B1(n_260),
.B2(n_249),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_285),
.Y(n_383)
);

OAI22x1_ASAP7_75t_L g360 ( 
.A1(n_281),
.A2(n_184),
.B1(n_142),
.B2(n_158),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_311),
.A2(n_263),
.B1(n_247),
.B2(n_279),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_279),
.A2(n_286),
.B1(n_250),
.B2(n_280),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_250),
.A2(n_317),
.B1(n_314),
.B2(n_312),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_374),
.A2(n_369),
.B1(n_361),
.B2(n_334),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_270),
.A2(n_278),
.B1(n_272),
.B2(n_237),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_376),
.A2(n_380),
.B1(n_287),
.B2(n_254),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_238),
.A2(n_268),
.B(n_257),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_300),
.A2(n_241),
.B1(n_316),
.B2(n_318),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_335),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_382),
.B(n_391),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_383),
.A2(n_386),
.B(n_389),
.Y(n_436)
);

NOR2x1_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_381),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_341),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_337),
.A2(n_233),
.B1(n_243),
.B2(n_255),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_287),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_387),
.B(n_426),
.C(n_329),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_333),
.B(n_287),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_392),
.Y(n_439)
);

AOI21xp33_ASAP7_75t_SL g389 ( 
.A1(n_326),
.A2(n_238),
.B(n_297),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_390),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_335),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_253),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_393),
.B(n_395),
.Y(n_469)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_394),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_397),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_352),
.A2(n_265),
.B(n_239),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_398),
.A2(n_408),
.B(n_417),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_400),
.B1(n_414),
.B2(n_429),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_374),
.A2(n_296),
.B1(n_277),
.B2(n_310),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_402),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_364),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_403),
.B(n_406),
.Y(n_445)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_324),
.Y(n_404)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_324),
.Y(n_405)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_344),
.B(n_275),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_344),
.B(n_292),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_415),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_SL g408 ( 
.A1(n_371),
.A2(n_304),
.B1(n_267),
.B2(n_291),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_332),
.A2(n_253),
.B(n_240),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_409),
.A2(n_412),
.B(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_410),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_332),
.A2(n_240),
.B(n_234),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_320),
.B(n_301),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_413),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_336),
.A2(n_299),
.B1(n_282),
.B2(n_259),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_261),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_353),
.B(n_262),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_416),
.B(n_421),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_340),
.A2(n_271),
.B(n_256),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_362),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_418),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_327),
.A2(n_322),
.B1(n_331),
.B2(n_356),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_419),
.A2(n_427),
.B(n_379),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_347),
.A2(n_254),
.B1(n_276),
.B2(n_297),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_423),
.B1(n_428),
.B2(n_431),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_345),
.B(n_362),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_340),
.A2(n_350),
.B1(n_330),
.B2(n_360),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_363),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_424),
.Y(n_438)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_348),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_425),
.B(n_430),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_326),
.C(n_320),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_363),
.A2(n_377),
.B(n_348),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_330),
.A2(n_360),
.B1(n_380),
.B2(n_348),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_358),
.A2(n_342),
.B1(n_376),
.B2(n_338),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_342),
.A2(n_338),
.B1(n_375),
.B2(n_367),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_434),
.A2(n_435),
.B(n_446),
.Y(n_491)
);

A2O1A1O1Ixp25_ASAP7_75t_L g435 ( 
.A1(n_384),
.A2(n_379),
.B(n_341),
.C(n_349),
.D(n_339),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_441),
.B(n_442),
.C(n_449),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_426),
.B(n_387),
.C(n_425),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_426),
.B(n_349),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_454),
.A2(n_458),
.B(n_459),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_339),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_455),
.B(n_462),
.C(n_472),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_392),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_466),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_411),
.A2(n_375),
.B1(n_367),
.B2(n_355),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_457),
.A2(n_464),
.B1(n_394),
.B2(n_390),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_398),
.A2(n_355),
.B(n_325),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_384),
.A2(n_325),
.B(n_359),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_329),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_422),
.A2(n_409),
.B(n_412),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_465),
.B(n_388),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_411),
.A2(n_328),
.B1(n_366),
.B2(n_378),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_422),
.A2(n_359),
.B(n_323),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_416),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_415),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_382),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_427),
.B(n_372),
.C(n_365),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_444),
.Y(n_474)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_474),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_451),
.A2(n_399),
.B1(n_385),
.B2(n_409),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_475),
.A2(n_476),
.B1(n_483),
.B2(n_505),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_451),
.A2(n_385),
.B1(n_412),
.B2(n_423),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_465),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_478),
.B(n_490),
.Y(n_540)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_444),
.Y(n_479)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_479),
.Y(n_525)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_447),
.Y(n_480)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_480),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_389),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_507),
.Y(n_517)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_447),
.Y(n_482)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_482),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_437),
.A2(n_385),
.B1(n_423),
.B2(n_400),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_484),
.A2(n_509),
.B1(n_452),
.B2(n_473),
.Y(n_533)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_453),
.Y(n_486)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_486),
.Y(n_546)
);

MAJx2_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_424),
.C(n_418),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_487),
.B(n_470),
.Y(n_527)
);

OA22x2_ASAP7_75t_L g488 ( 
.A1(n_432),
.A2(n_419),
.B1(n_428),
.B2(n_396),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_488),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_458),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_433),
.B(n_391),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_492),
.B(n_497),
.Y(n_514)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_453),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_493),
.B(n_494),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_495),
.A2(n_499),
.B(n_503),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_433),
.B(n_403),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_502),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_438),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_437),
.A2(n_428),
.B1(n_396),
.B2(n_431),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_498),
.A2(n_512),
.B1(n_478),
.B2(n_503),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_446),
.A2(n_401),
.B(n_383),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_500),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_449),
.B(n_407),
.C(n_406),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_513),
.C(n_448),
.Y(n_526)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_460),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_413),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_467),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_508),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_434),
.A2(n_400),
.B1(n_414),
.B2(n_431),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_455),
.B(n_417),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_468),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_463),
.A2(n_464),
.B1(n_457),
.B2(n_462),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_467),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_510),
.B(n_469),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_439),
.B(n_421),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_511),
.B(n_487),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_454),
.A2(n_420),
.B1(n_408),
.B2(n_413),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_439),
.B(n_413),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_454),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_524),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_498),
.A2(n_438),
.B1(n_445),
.B2(n_448),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_518),
.A2(n_521),
.B1(n_528),
.B2(n_530),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_483),
.A2(n_475),
.B1(n_476),
.B2(n_509),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_485),
.B(n_472),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_526),
.B(n_491),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_527),
.B(n_534),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_490),
.A2(n_445),
.B1(n_471),
.B2(n_456),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_505),
.A2(n_443),
.B1(n_452),
.B2(n_466),
.Y(n_530)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_531),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_485),
.B(n_470),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_532),
.B(n_536),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_548),
.B1(n_495),
.B2(n_503),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_496),
.A2(n_469),
.B1(n_443),
.B2(n_450),
.Y(n_535)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_489),
.B(n_450),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_489),
.B(n_436),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_537),
.B(n_539),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_512),
.A2(n_414),
.B1(n_436),
.B2(n_440),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_538),
.A2(n_551),
.B1(n_397),
.B2(n_343),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_507),
.B(n_435),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g541 ( 
.A(n_500),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_541),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_511),
.B(n_435),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_549),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_499),
.A2(n_440),
.B1(n_473),
.B2(n_420),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_501),
.B(n_513),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_477),
.B(n_404),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_550),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_547),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_552),
.B(n_565),
.C(n_523),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_553),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_514),
.B(n_365),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_554),
.B(n_555),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_536),
.B(n_430),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_579),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_524),
.B(n_532),
.C(n_517),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_558),
.B(n_569),
.C(n_573),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_540),
.A2(n_491),
.B(n_506),
.Y(n_563)
);

INVxp33_ASAP7_75t_L g609 ( 
.A(n_563),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_520),
.A2(n_506),
.B(n_488),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_529),
.A2(n_488),
.B(n_508),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_567),
.B(n_568),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_551),
.A2(n_488),
.B(n_386),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_517),
.B(n_405),
.C(n_410),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_519),
.Y(n_570)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_570),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_370),
.C(n_468),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_537),
.B(n_370),
.C(n_343),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_575),
.B(n_516),
.C(n_523),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_518),
.Y(n_576)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_576),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_526),
.B(n_372),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_577),
.B(n_569),
.Y(n_596)
);

FAx1_ASAP7_75t_SL g578 ( 
.A(n_527),
.B(n_323),
.CI(n_343),
.CON(n_578),
.SN(n_578)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_578),
.B(n_580),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_534),
.B(n_366),
.Y(n_579)
);

INVxp33_ASAP7_75t_L g580 ( 
.A(n_528),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_522),
.Y(n_581)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_581),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_520),
.B(n_548),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_546),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_583),
.A2(n_515),
.B1(n_521),
.B2(n_538),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_570),
.Y(n_584)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_584),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_585),
.A2(n_586),
.B1(n_583),
.B2(n_568),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_559),
.A2(n_530),
.B1(n_543),
.B2(n_539),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_574),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_587),
.B(n_604),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_560),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_593),
.B(n_608),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_594),
.A2(n_567),
.B(n_565),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_595),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_596),
.B(n_558),
.Y(n_610)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_599),
.B(n_603),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_602),
.A2(n_582),
.B(n_556),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_562),
.B(n_573),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_576),
.B(n_541),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_564),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_605),
.B(n_606),
.Y(n_620)
);

MAJx2_ASAP7_75t_L g606 ( 
.A(n_566),
.B(n_542),
.C(n_525),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_562),
.B(n_544),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_607),
.B(n_579),
.C(n_575),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_580),
.B(n_346),
.Y(n_608)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_610),
.Y(n_639)
);

NOR2xp67_ASAP7_75t_SL g638 ( 
.A(n_612),
.B(n_614),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_613),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_561),
.C(n_572),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g632 ( 
.A1(n_615),
.A2(n_616),
.B1(n_626),
.B2(n_590),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_588),
.A2(n_582),
.B1(n_553),
.B2(n_563),
.Y(n_616)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_617),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_584),
.B(n_572),
.Y(n_621)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_621),
.Y(n_642)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_591),
.A2(n_578),
.B(n_571),
.C(n_566),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_622),
.A2(n_625),
.B(n_617),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_589),
.B(n_561),
.C(n_571),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_623),
.B(n_630),
.C(n_606),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_597),
.B(n_578),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_624),
.B(n_601),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_591),
.A2(n_397),
.B(n_328),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_588),
.A2(n_378),
.B1(n_373),
.B2(n_346),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g629 ( 
.A1(n_609),
.A2(n_321),
.B(n_590),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_629),
.A2(n_611),
.B(n_626),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_603),
.B(n_321),
.C(n_599),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_632),
.A2(n_640),
.B1(n_645),
.B2(n_618),
.Y(n_655)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_612),
.B(n_607),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_633),
.B(n_635),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_615),
.A2(n_598),
.B1(n_585),
.B2(n_602),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_634),
.B(n_643),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_610),
.B(n_592),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_641),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_616),
.A2(n_586),
.B1(n_609),
.B2(n_604),
.Y(n_640)
);

INVxp67_ASAP7_75t_L g641 ( 
.A(n_620),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_SL g644 ( 
.A1(n_624),
.A2(n_595),
.B(n_601),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_644),
.A2(n_647),
.B(n_629),
.Y(n_651)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_613),
.A2(n_321),
.B1(n_600),
.B2(n_620),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_646),
.B(n_622),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_619),
.B(n_627),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_648),
.B(n_643),
.Y(n_660)
);

AOI221xp5_ASAP7_75t_L g649 ( 
.A1(n_639),
.A2(n_611),
.B1(n_628),
.B2(n_625),
.C(n_619),
.Y(n_649)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_649),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_637),
.B(n_627),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_650),
.B(n_654),
.Y(n_665)
);

XOR2x2_ASAP7_75t_L g666 ( 
.A(n_651),
.B(n_655),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_633),
.B(n_630),
.C(n_614),
.Y(n_654)
);

NOR2xp67_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_623),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_656),
.A2(n_658),
.B(n_645),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_631),
.A2(n_621),
.B(n_618),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_635),
.B(n_632),
.C(n_640),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_659),
.B(n_660),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_641),
.B(n_628),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_661),
.B(n_642),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_662),
.A2(n_646),
.B(n_631),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_654),
.B(n_644),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_663),
.B(n_671),
.Y(n_676)
);

AOI21xp33_ASAP7_75t_L g673 ( 
.A1(n_664),
.A2(n_667),
.B(n_651),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_669),
.Y(n_674)
);

BUFx24_ASAP7_75t_SL g671 ( 
.A(n_652),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g672 ( 
.A(n_657),
.B(n_642),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_672),
.B(n_658),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_673),
.A2(n_675),
.B(n_677),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_665),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_670),
.B(n_659),
.C(n_653),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_678),
.B(n_675),
.C(n_676),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_SL g679 ( 
.A1(n_674),
.A2(n_668),
.B(n_666),
.C(n_662),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_679),
.B(n_680),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_681),
.B(n_653),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g684 ( 
.A(n_683),
.B(n_666),
.C(n_655),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_684),
.A2(n_682),
.B1(n_634),
.B2(n_647),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_685),
.Y(n_686)
);


endmodule