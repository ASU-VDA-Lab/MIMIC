module fake_ariane_505_n_94 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_10, n_94);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_10;

output n_94;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_92;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_88;
wire n_68;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_35;
wire n_54;
wire n_25;

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_21),
.B1(n_22),
.B2(n_14),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AND2x6_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_18),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx6p67_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_5),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AND2x4_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_17),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_8),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_23),
.A2(n_31),
.B1(n_36),
.B2(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_25),
.B(n_28),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_24),
.B(n_40),
.Y(n_51)
);

NAND2x1_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

OAI21x1_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_24),
.B(n_32),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_26),
.B(n_29),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_41),
.B(n_46),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_42),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_45),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_35),
.B(n_29),
.C(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_66),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_59),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_64),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_71),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_71),
.B1(n_38),
.B2(n_64),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_62),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

NOR4xp25_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_68),
.C(n_74),
.D(n_75),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_43),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_80),
.C(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_81),
.Y(n_85)
);

NAND4xp75_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_27),
.C(n_33),
.D(n_34),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_45),
.Y(n_87)
);

OAI211xp5_ASAP7_75t_SL g88 ( 
.A1(n_84),
.A2(n_82),
.B(n_27),
.C(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_27),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_33),
.B1(n_34),
.B2(n_27),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_34),
.B(n_48),
.C(n_49),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_90),
.B(n_89),
.Y(n_93)
);

AOI221xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_48),
.B1(n_49),
.B2(n_92),
.C(n_56),
.Y(n_94)
);


endmodule