module fake_jpeg_11836_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_20),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_0),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_52),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_72),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_81),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_60),
.B1(n_50),
.B2(n_55),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_80),
.A2(n_62),
.B1(n_54),
.B2(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_57),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_51),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_67),
.B1(n_50),
.B2(n_55),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_100),
.B1(n_47),
.B2(n_2),
.Y(n_106)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_53),
.C(n_26),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_91),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_65),
.B1(n_49),
.B2(n_51),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_76),
.A2(n_49),
.B1(n_59),
.B2(n_56),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_75),
.B(n_0),
.C(n_1),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_4),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_119)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_101),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_114),
.B1(n_90),
.B2(n_12),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_119),
.Y(n_135)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_122),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_100),
.A2(n_9),
.B(n_10),
.Y(n_118)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_43),
.B(n_21),
.C(n_22),
.D(n_24),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_125),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_120),
.B1(n_111),
.B2(n_118),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_16),
.C(n_18),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_131),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_42),
.C(n_25),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_19),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_145),
.B1(n_134),
.B2(n_113),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_133),
.C(n_136),
.Y(n_143)
);

AOI321xp33_ASAP7_75t_L g146 ( 
.A1(n_143),
.A2(n_144),
.A3(n_138),
.B1(n_136),
.B2(n_113),
.C(n_134),
.Y(n_146)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_141),
.B(n_135),
.C(n_123),
.Y(n_144)
);

AOI322xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_135),
.A3(n_130),
.B1(n_120),
.B2(n_108),
.C1(n_112),
.C2(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_28),
.B(n_29),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_30),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_32),
.B(n_35),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_37),
.C(n_39),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_41),
.Y(n_154)
);


endmodule