module fake_jpeg_8658_n_173 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_31),
.A2(n_20),
.B1(n_24),
.B2(n_23),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_20),
.B1(n_31),
.B2(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_65),
.B1(n_41),
.B2(n_38),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_62),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_61),
.Y(n_81)
);

INVxp67_ASAP7_75t_SL g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_68),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_35),
.B1(n_32),
.B2(n_37),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_20),
.B1(n_31),
.B2(n_35),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_37),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_16),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_86),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_67),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_75),
.Y(n_91)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_29),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_51),
.B1(n_37),
.B2(n_30),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_30),
.B(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_29),
.B1(n_19),
.B2(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_64),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_98),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_48),
.C(n_32),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_101),
.C(n_94),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_96),
.B(n_84),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_76),
.B(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_36),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

AO221x1_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_75),
.B1(n_81),
.B2(n_64),
.C(n_82),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_30),
.C(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_102),
.B(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_108),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_116),
.B(n_101),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_89),
.B(n_17),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_109),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_113),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_15),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_39),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_117),
.C(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_15),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_16),
.Y(n_126)
);

AOI22x1_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_36),
.B1(n_26),
.B2(n_22),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_57),
.C(n_17),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_88),
.C(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_125),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_95),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_120),
.A2(n_123),
.B(n_131),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_127),
.A2(n_28),
.B1(n_14),
.B2(n_23),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_117),
.B(n_114),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_100),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_142),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_92),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_26),
.C(n_27),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_129),
.A2(n_120),
.B1(n_123),
.B2(n_121),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_26),
.B1(n_27),
.B2(n_8),
.Y(n_147)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_28),
.B1(n_24),
.B2(n_18),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_130),
.B(n_128),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_139),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_SL g141 ( 
.A(n_119),
.B(n_14),
.C(n_18),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_6),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_57),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_142),
.C(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_147),
.B(n_150),
.Y(n_156)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_0),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_154),
.Y(n_159)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_145),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_157),
.B1(n_156),
.B2(n_158),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_141),
.B1(n_140),
.B2(n_8),
.Y(n_157)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_5),
.C(n_12),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_9),
.B(n_1),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_149),
.A3(n_151),
.B1(n_143),
.B2(n_9),
.C1(n_10),
.C2(n_6),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_152),
.B(n_2),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_162),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_163),
.B(n_1),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_167),
.C(n_160),
.Y(n_168)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_3),
.B(n_4),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_159),
.A2(n_2),
.B(n_3),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_165),
.B(n_3),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_169),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_171),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.Y(n_173)
);


endmodule