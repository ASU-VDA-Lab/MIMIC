module fake_aes_3207_n_573 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_573);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_573;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_64), .Y(n_80) );
NOR2xp33_ASAP7_75t_L g81 ( .A(n_69), .B(n_57), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_78), .Y(n_82) );
INVx1_ASAP7_75t_SL g83 ( .A(n_59), .Y(n_83) );
CKINVDCx14_ASAP7_75t_R g84 ( .A(n_5), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_66), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
INVxp67_ASAP7_75t_L g87 ( .A(n_79), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_10), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_41), .Y(n_90) );
XOR2xp5_ASAP7_75t_L g91 ( .A(n_74), .B(n_23), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_1), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_11), .Y(n_94) );
CKINVDCx14_ASAP7_75t_R g95 ( .A(n_71), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_7), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_77), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_26), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_13), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_17), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_48), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_37), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_63), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_1), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_32), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_22), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_31), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_33), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_35), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_21), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_8), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_90), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_82), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_96), .B(n_0), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_115), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_92), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_102), .B(n_0), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_115), .B(n_2), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g127 ( .A(n_103), .B(n_40), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_80), .B(n_2), .Y(n_128) );
AND2x2_ASAP7_75t_L g129 ( .A(n_95), .B(n_3), .Y(n_129) );
AND2x2_ASAP7_75t_L g130 ( .A(n_102), .B(n_3), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_92), .B(n_4), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_89), .B(n_4), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_89), .B(n_5), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_98), .Y(n_137) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_91), .A2(n_6), .B1(n_8), .B2(n_9), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_103), .Y(n_139) );
NOR2xp67_ASAP7_75t_L g140 ( .A(n_87), .B(n_6), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_124), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_139), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_124), .B(n_94), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx3_ASAP7_75t_L g146 ( .A(n_124), .Y(n_146) );
INVx4_ASAP7_75t_SL g147 ( .A(n_124), .Y(n_147) );
BUFx10_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
AND2x2_ASAP7_75t_L g149 ( .A(n_139), .B(n_105), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_118), .B(n_113), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
BUFx2_ASAP7_75t_L g152 ( .A(n_129), .Y(n_152) );
OR2x2_ASAP7_75t_L g153 ( .A(n_120), .B(n_106), .Y(n_153) );
INVxp67_ASAP7_75t_SL g154 ( .A(n_129), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_118), .B(n_122), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_137), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_137), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_137), .Y(n_158) );
INVx5_ASAP7_75t_L g159 ( .A(n_116), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_116), .Y(n_160) );
OR2x2_ASAP7_75t_L g161 ( .A(n_119), .B(n_99), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_121), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_122), .B(n_97), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_121), .Y(n_165) );
INVx5_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
OR2x6_ASAP7_75t_L g168 ( .A(n_138), .B(n_91), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_155), .A2(n_134), .B(n_131), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_162), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_149), .B(n_127), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_162), .B(n_125), .Y(n_172) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_162), .B(n_133), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_166), .B(n_125), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_167), .Y(n_176) );
NOR2xp67_ASAP7_75t_L g177 ( .A(n_153), .B(n_126), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_167), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_167), .B(n_105), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_166), .B(n_131), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_167), .B(n_136), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_166), .B(n_134), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_152), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_143), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_147), .B(n_136), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_166), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_147), .B(n_140), .Y(n_189) );
NOR2xp33_ASAP7_75t_R g190 ( .A(n_148), .B(n_111), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_152), .B(n_135), .Y(n_191) );
NOR3xp33_ASAP7_75t_SL g192 ( .A(n_164), .B(n_138), .C(n_110), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_144), .A2(n_135), .B(n_132), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_142), .B(n_140), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_154), .B(n_123), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g196 ( .A1(n_150), .A2(n_88), .B(n_114), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_166), .B(n_128), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_148), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_142), .B(n_110), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_143), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_141), .B(n_113), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_141), .B(n_144), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_141), .B(n_123), .Y(n_204) );
NOR2x2_ASAP7_75t_L g205 ( .A(n_168), .B(n_98), .Y(n_205) );
AO22x1_ASAP7_75t_L g206 ( .A1(n_199), .A2(n_144), .B1(n_146), .B2(n_141), .Y(n_206) );
INVx4_ASAP7_75t_L g207 ( .A(n_173), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_173), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_180), .B(n_148), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_173), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_204), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_185), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_177), .B(n_161), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_183), .B(n_161), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_186), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_183), .B(n_144), .Y(n_216) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_203), .A2(n_169), .B(n_174), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_178), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_183), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_199), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_191), .B(n_153), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_172), .A2(n_146), .B(n_165), .C(n_163), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_180), .B(n_147), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_187), .B(n_148), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_201), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_187), .Y(n_227) );
O2A1O1Ixp5_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_151), .B(n_160), .C(n_163), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_201), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_178), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_187), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_191), .B(n_147), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_170), .B(n_146), .Y(n_233) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_189), .B(n_88), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_195), .B(n_165), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_170), .A2(n_168), .B1(n_163), .B2(n_160), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_176), .Y(n_237) );
NAND2x1p5_ASAP7_75t_L g238 ( .A(n_179), .B(n_151), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_195), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_196), .A2(n_168), .B1(n_160), .B2(n_151), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_202), .A2(n_145), .B(n_157), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_222), .B(n_185), .Y(n_242) );
INVxp67_ASAP7_75t_SL g243 ( .A(n_220), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_228), .A2(n_198), .B(n_193), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_241), .A2(n_143), .B(n_101), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_223), .A2(n_101), .B(n_160), .Y(n_246) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_210), .Y(n_247) );
INVx4_ASAP7_75t_L g248 ( .A(n_207), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_211), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_217), .A2(n_182), .B(n_184), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_236), .A2(n_168), .B1(n_194), .B2(n_181), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
BUFx12f_ASAP7_75t_L g253 ( .A(n_207), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_SL g254 ( .A1(n_220), .A2(n_175), .B(n_197), .C(n_188), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_207), .B(n_189), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_236), .A2(n_168), .B1(n_190), .B2(n_194), .Y(n_256) );
OAI21x1_ASAP7_75t_L g257 ( .A1(n_217), .A2(n_151), .B(n_114), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_240), .A2(n_112), .B(n_157), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_215), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_214), .B(n_194), .Y(n_261) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_240), .A2(n_112), .B(n_145), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_207), .B(n_189), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_210), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_215), .A2(n_156), .B(n_100), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_218), .A2(n_194), .B(n_200), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_216), .A2(n_156), .B(n_104), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_237), .Y(n_268) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_232), .A2(n_109), .B(n_107), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_210), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_243), .A2(n_234), .B1(n_239), .B2(n_208), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_212), .B1(n_234), .B2(n_209), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_213), .B1(n_192), .B2(n_239), .C(n_212), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_266), .A2(n_226), .B(n_218), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_243), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_251), .A2(n_234), .B1(n_210), .B2(n_221), .Y(n_276) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_257), .A2(n_108), .B(n_218), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_249), .B(n_208), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_251), .A2(n_210), .B1(n_224), .B2(n_231), .Y(n_279) );
OR2x2_ASAP7_75t_L g280 ( .A(n_261), .B(n_210), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_266), .A2(n_229), .B(n_226), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_253), .A2(n_224), .B1(n_227), .B2(n_237), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_253), .A2(n_227), .B1(n_225), .B2(n_235), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_249), .A2(n_238), .B1(n_226), .B2(n_229), .Y(n_284) );
AOI21xp33_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_230), .B(n_219), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_252), .B(n_229), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_252), .B(n_238), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_261), .A2(n_205), .B(n_93), .Y(n_288) );
OAI21xp33_ASAP7_75t_L g289 ( .A1(n_250), .A2(n_233), .B(n_238), .Y(n_289) );
AOI222xp33_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_205), .B1(n_206), .B2(n_83), .C1(n_230), .C2(n_219), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_257), .A2(n_81), .B(n_206), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_248), .Y(n_292) );
AO21x2_ASAP7_75t_L g293 ( .A1(n_257), .A2(n_230), .B(n_219), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_248), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_292), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_277), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_292), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_273), .A2(n_248), .B1(n_255), .B2(n_268), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_286), .B(n_248), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_286), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_273), .A2(n_255), .B1(n_268), .B2(n_269), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_260), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_280), .B(n_258), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_271), .A2(n_258), .B1(n_260), .B2(n_255), .Y(n_307) );
AO31x2_ASAP7_75t_L g308 ( .A1(n_284), .A2(n_258), .A3(n_260), .B(n_262), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
INVx4_ASAP7_75t_L g311 ( .A(n_294), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_287), .B(n_270), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_277), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_293), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_280), .B(n_270), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_271), .B(n_247), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_284), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_293), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_297), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_303), .B(n_287), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_297), .Y(n_322) );
NAND4xp25_ASAP7_75t_L g323 ( .A(n_300), .B(n_290), .C(n_288), .D(n_272), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_309), .Y(n_324) );
OAI33xp33_ASAP7_75t_L g325 ( .A1(n_307), .A2(n_289), .A3(n_10), .B1(n_11), .B2(n_12), .B3(n_13), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_304), .A2(n_288), .B1(n_290), .B2(n_276), .C(n_283), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_303), .B(n_279), .C(n_282), .D(n_285), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_296), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_311), .B(n_263), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_307), .A2(n_285), .B1(n_289), .B2(n_291), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_309), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_310), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_298), .B(n_293), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_305), .B(n_293), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_318), .A2(n_250), .B1(n_281), .B2(n_274), .C(n_269), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_298), .B(n_247), .Y(n_339) );
AND2x4_ASAP7_75t_SL g340 ( .A(n_301), .B(n_255), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_310), .Y(n_341) );
BUFx3_ASAP7_75t_L g342 ( .A(n_295), .Y(n_342) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_295), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_316), .B(n_291), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_305), .B(n_291), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_313), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_313), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_313), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_314), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_323), .B(n_299), .C(n_311), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_337), .B(n_316), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_337), .B(n_318), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_321), .B(n_302), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_336), .B(n_302), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_324), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_320), .Y(n_357) );
OAI31xp33_ASAP7_75t_L g358 ( .A1(n_323), .A2(n_301), .A3(n_263), .B(n_317), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_345), .B(n_314), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_345), .B(n_314), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g362 ( .A(n_325), .B(n_311), .C(n_299), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_320), .B(n_317), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_333), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_320), .B(n_308), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_320), .B(n_308), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_328), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_341), .B(n_308), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_328), .B(n_299), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_341), .B(n_347), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_350), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_343), .B(n_306), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_347), .B(n_308), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_348), .B(n_308), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_350), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_348), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_328), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_319), .B(n_308), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_319), .B(n_312), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_322), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_322), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_339), .B(n_306), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_334), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_334), .B(n_312), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_335), .B(n_315), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_339), .B(n_315), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_346), .B(n_315), .Y(n_388) );
NAND2x1_ASAP7_75t_L g389 ( .A(n_328), .B(n_301), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_346), .B(n_315), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_342), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_349), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_326), .B(n_301), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_342), .B(n_311), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_335), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_330), .B(n_269), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_356), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_353), .B(n_344), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_396), .B(n_342), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_396), .B(n_344), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_355), .B(n_340), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_358), .A2(n_327), .B1(n_329), .B2(n_340), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_384), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_384), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_361), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_358), .A2(n_331), .B1(n_329), .B2(n_332), .C(n_338), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_364), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_367), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_389), .B(n_259), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_367), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_372), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_391), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_351), .A2(n_340), .B1(n_254), .B2(n_269), .C(n_270), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_353), .B(n_291), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_354), .B(n_9), .Y(n_420) );
NOR3xp33_ASAP7_75t_SL g421 ( .A(n_351), .B(n_12), .C(n_14), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_359), .B(n_262), .Y(n_422) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_368), .B(n_267), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_352), .B(n_259), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_352), .B(n_259), .Y(n_425) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_368), .B(n_267), .Y(n_426) );
INVxp67_ASAP7_75t_L g427 ( .A(n_378), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_359), .B(n_262), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_360), .B(n_14), .Y(n_429) );
INVxp33_ASAP7_75t_L g430 ( .A(n_389), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_386), .B(n_15), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_392), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_392), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_360), .B(n_15), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_372), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_388), .B(n_246), .Y(n_436) );
INVxp67_ASAP7_75t_SL g437 ( .A(n_370), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_376), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_388), .B(n_246), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_376), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_373), .B(n_16), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_393), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_377), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_380), .B(n_16), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_395), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_380), .B(n_385), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_386), .B(n_267), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_385), .B(n_267), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_371), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_393), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_390), .B(n_246), .Y(n_451) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_406), .A2(n_362), .B1(n_370), .B2(n_368), .C(n_394), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_430), .A2(n_368), .B(n_395), .C(n_383), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_399), .B(n_390), .Y(n_454) );
OAI222xp33_ASAP7_75t_L g455 ( .A1(n_437), .A2(n_370), .B1(n_395), .B2(n_387), .C1(n_397), .C2(n_377), .Y(n_455) );
NOR2x1_ASAP7_75t_L g456 ( .A(n_417), .B(n_395), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_449), .B(n_371), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_446), .B(n_374), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_406), .A2(n_382), .B1(n_381), .B2(n_375), .Y(n_459) );
INVxp67_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_430), .A2(n_374), .B(n_369), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_407), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_411), .A2(n_375), .B1(n_369), .B2(n_363), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_399), .B(n_363), .Y(n_464) );
OAI21xp33_ASAP7_75t_L g465 ( .A1(n_421), .A2(n_365), .B(n_366), .Y(n_465) );
AOI32xp33_ASAP7_75t_L g466 ( .A1(n_418), .A2(n_366), .A3(n_365), .B1(n_379), .B2(n_382), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_398), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_407), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_401), .Y(n_469) );
AOI322xp5_ASAP7_75t_L g470 ( .A1(n_420), .A2(n_379), .A3(n_381), .B1(n_357), .B2(n_264), .C1(n_270), .C2(n_159), .Y(n_470) );
NOR4xp25_ASAP7_75t_SL g471 ( .A(n_416), .B(n_357), .C(n_255), .D(n_264), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_404), .B(n_264), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_403), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_409), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_445), .B(n_245), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_400), .A2(n_265), .B(n_245), .C(n_244), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g477 ( .A1(n_431), .A2(n_255), .B1(n_263), .B2(n_159), .Y(n_477) );
OAI22x1_ASAP7_75t_L g478 ( .A1(n_427), .A2(n_263), .B1(n_159), .B2(n_24), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_410), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_405), .B(n_245), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_441), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_435), .B(n_244), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_431), .B(n_18), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_408), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_412), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_413), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_415), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_422), .B(n_244), .Y(n_488) );
AOI21xp5_ASAP7_75t_SL g489 ( .A1(n_414), .A2(n_265), .B(n_25), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_419), .A2(n_159), .B1(n_265), .B2(n_158), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_424), .B(n_159), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_438), .Y(n_492) );
NOR4xp25_ASAP7_75t_SL g493 ( .A(n_440), .B(n_19), .C(n_27), .D(n_28), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_419), .B(n_159), .Y(n_494) );
AND2x2_ASAP7_75t_SL g495 ( .A(n_424), .B(n_29), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_423), .A2(n_158), .B(n_38), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_444), .B(n_36), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_425), .A2(n_158), .B1(n_42), .B2(n_43), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_454), .B(n_422), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_466), .B(n_429), .C(n_434), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_463), .B(n_443), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_457), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g503 ( .A1(n_456), .A2(n_414), .B1(n_425), .B2(n_448), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_461), .B(n_428), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_457), .B(n_428), .Y(n_505) );
OAI222xp33_ASAP7_75t_L g506 ( .A1(n_459), .A2(n_426), .B1(n_447), .B2(n_448), .C1(n_436), .C2(n_451), .Y(n_506) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_459), .A2(n_408), .B1(n_450), .B2(n_432), .C(n_442), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_458), .B(n_447), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_460), .B(n_451), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_467), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_465), .B(n_450), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_469), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_481), .B(n_442), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_453), .A2(n_433), .B(n_432), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_464), .B(n_433), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_473), .B(n_439), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_474), .Y(n_518) );
AOI21xp33_ASAP7_75t_SL g519 ( .A1(n_495), .A2(n_439), .B(n_436), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_479), .B(n_158), .Y(n_520) );
NOR2xp67_ASAP7_75t_L g521 ( .A(n_478), .B(n_39), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_452), .B(n_455), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_485), .Y(n_523) );
XNOR2xp5_ASAP7_75t_L g524 ( .A(n_477), .B(n_44), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_486), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_487), .Y(n_526) );
OAI211xp5_ASAP7_75t_L g527 ( .A1(n_471), .A2(n_158), .B(n_46), .C(n_47), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_496), .A2(n_158), .B(n_49), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_477), .A2(n_45), .B(n_50), .C(n_51), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_522), .A2(n_491), .B1(n_496), .B2(n_498), .Y(n_530) );
XNOR2xp5_ASAP7_75t_L g531 ( .A(n_500), .B(n_492), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_522), .B(n_498), .Y(n_532) );
OAI211xp5_ASAP7_75t_L g533 ( .A1(n_521), .A2(n_470), .B(n_483), .C(n_497), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_501), .B(n_488), .Y(n_534) );
XNOR2xp5_ASAP7_75t_L g535 ( .A(n_524), .B(n_472), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_503), .Y(n_536) );
OAI21xp33_ASAP7_75t_L g537 ( .A1(n_504), .A2(n_494), .B(n_480), .Y(n_537) );
NOR2xp33_ASAP7_75t_SL g538 ( .A(n_506), .B(n_475), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_510), .Y(n_540) );
AOI32xp33_ASAP7_75t_L g541 ( .A1(n_507), .A2(n_484), .A3(n_468), .B1(n_490), .B2(n_482), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_512), .Y(n_542) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_527), .A2(n_489), .B(n_476), .Y(n_543) );
AOI211xp5_ASAP7_75t_L g544 ( .A1(n_519), .A2(n_482), .B(n_493), .C(n_55), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_513), .A2(n_52), .B1(n_54), .B2(n_56), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_518), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_513), .B(n_60), .Y(n_547) );
NAND4xp25_ASAP7_75t_L g548 ( .A(n_532), .B(n_544), .C(n_538), .D(n_543), .Y(n_548) );
AOI22xp5_ASAP7_75t_SL g549 ( .A1(n_536), .A2(n_511), .B1(n_528), .B2(n_514), .Y(n_549) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_530), .A2(n_529), .B(n_520), .C(n_508), .Y(n_550) );
OAI211xp5_ASAP7_75t_SL g551 ( .A1(n_541), .A2(n_526), .B(n_525), .C(n_523), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_540), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_539), .B(n_509), .Y(n_553) );
AOI211x1_ASAP7_75t_SL g554 ( .A1(n_534), .A2(n_516), .B(n_515), .C(n_505), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_542), .Y(n_555) );
NAND4xp75_ASAP7_75t_L g556 ( .A(n_547), .B(n_499), .C(n_517), .D(n_529), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_546), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_553), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_552), .B(n_537), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_555), .Y(n_560) );
OAI21xp33_ASAP7_75t_L g561 ( .A1(n_548), .A2(n_538), .B(n_531), .Y(n_561) );
NOR4xp25_ASAP7_75t_L g562 ( .A(n_551), .B(n_533), .C(n_517), .D(n_499), .Y(n_562) );
OR4x2_ASAP7_75t_L g563 ( .A(n_561), .B(n_562), .C(n_549), .D(n_556), .Y(n_563) );
NOR2x2_ASAP7_75t_L g564 ( .A(n_558), .B(n_550), .Y(n_564) );
OAI22xp5_ASAP7_75t_SL g565 ( .A1(n_559), .A2(n_535), .B1(n_554), .B2(n_545), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_563), .Y(n_566) );
AOI21xp33_ASAP7_75t_L g567 ( .A1(n_565), .A2(n_560), .B(n_557), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_566), .A2(n_564), .B1(n_553), .B2(n_65), .Y(n_568) );
OAI22xp5_ASAP7_75t_SL g569 ( .A1(n_567), .A2(n_61), .B1(n_62), .B2(n_67), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_569), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g571 ( .A1(n_570), .A2(n_568), .B1(n_70), .B2(n_73), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_571), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_572), .A2(n_68), .B1(n_75), .B2(n_76), .Y(n_573) );
endmodule