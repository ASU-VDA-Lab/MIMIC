module fake_jpeg_9560_n_295 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_48),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_29),
.B1(n_19),
.B2(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_35),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_26),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_35),
.C(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_19),
.B1(n_30),
.B2(n_28),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_27),
.B1(n_26),
.B2(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_70),
.Y(n_113)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_71),
.B(n_87),
.Y(n_130)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_77),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_79),
.Y(n_120)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_80),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_94),
.B1(n_101),
.B2(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_18),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_98),
.Y(n_105)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_96),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_27),
.B1(n_22),
.B2(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_57),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_26),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_55),
.B(n_18),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_25),
.B1(n_22),
.B2(n_24),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_70),
.B1(n_49),
.B2(n_53),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_48),
.C(n_43),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_114),
.C(n_101),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_98),
.A2(n_28),
.B(n_20),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_20),
.B(n_30),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_121),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_43),
.C(n_53),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_91),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_68),
.B1(n_20),
.B2(n_83),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_65),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_71),
.B(n_103),
.C(n_97),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_128),
.Y(n_158)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_65),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_129),
.B(n_131),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_33),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_130),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g134 ( 
.A(n_111),
.B(n_86),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_151),
.B(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_139),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_79),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_137),
.B(n_147),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_144),
.B1(n_145),
.B2(n_152),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_32),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_23),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_149),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_49),
.B1(n_53),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_100),
.B1(n_83),
.B2(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_146),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_157),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_99),
.B(n_23),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_69),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_119),
.A2(n_69),
.B1(n_33),
.B2(n_31),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_33),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_161),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_115),
.A2(n_105),
.B1(n_123),
.B2(n_121),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_156),
.B1(n_138),
.B2(n_153),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_33),
.B1(n_31),
.B2(n_21),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_107),
.A2(n_23),
.B(n_31),
.C(n_21),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_159),
.A2(n_129),
.B(n_110),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_31),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_1),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_177),
.C(n_132),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_184),
.B(n_148),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_150),
.A2(n_116),
.B1(n_129),
.B2(n_125),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_178),
.B(n_10),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_182),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_176),
.A2(n_187),
.B1(n_159),
.B2(n_21),
.Y(n_204)
);

NOR2x1_ASAP7_75t_R g178 ( 
.A(n_134),
.B(n_23),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_118),
.Y(n_179)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_145),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_124),
.B(n_117),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_185),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_134),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_11),
.Y(n_214)
);

AO21x2_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_104),
.B(n_106),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_127),
.B1(n_125),
.B2(n_106),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_191),
.A2(n_135),
.B1(n_157),
.B2(n_124),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_197),
.C(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_196),
.B(n_190),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_137),
.C(n_140),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_204),
.B(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_158),
.C(n_155),
.Y(n_200)
);

OAI322xp33_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_151),
.A3(n_148),
.B1(n_147),
.B2(n_159),
.C1(n_149),
.C2(n_156),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_SL g227 ( 
.A(n_202),
.B(n_209),
.C(n_184),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_159),
.B1(n_117),
.B2(n_21),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_186),
.A2(n_187),
.B1(n_179),
.B2(n_174),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_206),
.B1(n_167),
.B2(n_164),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_159),
.B1(n_18),
.B2(n_23),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_2),
.Y(n_207)
);

AOI221xp5_ASAP7_75t_L g209 ( 
.A1(n_170),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_210),
.B(n_215),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_211)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_169),
.B(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_11),
.Y(n_216)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_216),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_183),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_217),
.B(n_226),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_205),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_227),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_231),
.B(n_207),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_216),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_163),
.C(n_177),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_200),
.C(n_198),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_230),
.A2(n_232),
.B1(n_234),
.B2(n_204),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_170),
.B(n_167),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_175),
.B1(n_166),
.B2(n_168),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_215),
.B(n_171),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_233),
.B(n_212),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_194),
.A2(n_168),
.B1(n_190),
.B2(n_172),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_201),
.Y(n_251)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_236),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_221),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_197),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_242),
.C(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_222),
.A2(n_199),
.B(n_207),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_248),
.B(n_250),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_228),
.C(n_198),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_210),
.C(n_206),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_230),
.C(n_220),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_195),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_231),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_212),
.B1(n_201),
.B2(n_13),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_217),
.Y(n_260)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_264),
.C(n_241),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_263),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_218),
.B1(n_219),
.B2(n_236),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_245),
.B1(n_218),
.B2(n_252),
.Y(n_271)
);

NOR2x1p5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_227),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_262),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_260),
.B(n_224),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_232),
.C(n_223),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_242),
.C(n_239),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_270),
.C(n_274),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_272),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_238),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_262),
.A2(n_223),
.B1(n_224),
.B2(n_237),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_256),
.B1(n_258),
.B2(n_14),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_11),
.B(n_12),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_258),
.B(n_13),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_282),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_280),
.B(n_281),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_16),
.Y(n_281)
);

AOI31xp33_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_12),
.A3(n_13),
.B(n_14),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_270),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_287),
.B(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_283),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_266),
.C(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_291),
.C(n_286),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_15),
.B(n_289),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_15),
.Y(n_295)
);


endmodule