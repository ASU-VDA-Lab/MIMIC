module fake_jpeg_7720_n_208 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_82;
wire n_96;

BUFx24_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_11),
.B(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_47),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_40),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_0),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_55),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_44),
.A2(n_32),
.B1(n_34),
.B2(n_21),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_35),
.B1(n_43),
.B2(n_18),
.Y(n_77)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_20),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_59),
.B(n_65),
.Y(n_82)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g63 ( 
.A(n_35),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_18),
.Y(n_74)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_69),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_20),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_72),
.Y(n_99)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_22),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_95),
.B(n_71),
.Y(n_113)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_81),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_77),
.A2(n_88),
.B1(n_49),
.B2(n_68),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_38),
.B1(n_36),
.B2(n_43),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_49),
.B1(n_62),
.B2(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_70),
.A2(n_22),
.B1(n_25),
.B2(n_29),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_83),
.A2(n_76),
.B1(n_85),
.B2(n_97),
.Y(n_118)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_87),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_30),
.B1(n_28),
.B2(n_21),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g89 ( 
.A(n_55),
.B(n_38),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_27),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_23),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_36),
.Y(n_106)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_29),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_71),
.B1(n_64),
.B2(n_24),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_100),
.B(n_26),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_113),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_36),
.B(n_47),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_89),
.C(n_100),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_107),
.B1(n_111),
.B2(n_91),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_81),
.B(n_16),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_114),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_74),
.A2(n_52),
.B(n_50),
.C(n_23),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_73),
.A2(n_2),
.B(n_3),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_94),
.B1(n_79),
.B2(n_31),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_24),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_50),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_93),
.B1(n_98),
.B2(n_84),
.Y(n_125)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_76),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_133),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_131),
.A2(n_120),
.B(n_101),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_85),
.B1(n_80),
.B2(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_75),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_78),
.B1(n_86),
.B2(n_91),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_106),
.B(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_144),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_142),
.B1(n_79),
.B2(n_123),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_122),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_143),
.A2(n_79),
.B1(n_103),
.B2(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_82),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.C(n_154),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_101),
.C(n_103),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_150),
.A2(n_157),
.B1(n_9),
.B2(n_5),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_138),
.A2(n_114),
.B(n_105),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_2),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_138),
.A2(n_121),
.B(n_112),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_158),
.B(n_160),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_112),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_121),
.B(n_116),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_156),
.A2(n_137),
.B1(n_139),
.B2(n_130),
.C(n_124),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_108),
.B(n_119),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_123),
.B(n_3),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_134),
.B1(n_143),
.B2(n_125),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_164),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_144),
.C(n_137),
.Y(n_167)
);

OAI321xp33_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_124),
.A3(n_132),
.B1(n_128),
.B2(n_135),
.C(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_152),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_158),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_161),
.A2(n_128),
.B1(n_16),
.B2(n_15),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_12),
.Y(n_172)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_172),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_171),
.B(n_162),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_154),
.C(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_182),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_145),
.C(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_183),
.B(n_184),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

OA21x2_ASAP7_75t_SL g187 ( 
.A1(n_177),
.A2(n_171),
.B(n_173),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_188),
.B(n_180),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_168),
.CI(n_160),
.CON(n_189),
.SN(n_189)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_189),
.A2(n_191),
.B1(n_181),
.B2(n_149),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_149),
.B1(n_166),
.B2(n_157),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_190),
.B(n_179),
.C(n_175),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_193),
.C(n_4),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_175),
.C(n_176),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_196),
.B(n_189),
.C(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_185),
.A2(n_151),
.B1(n_5),
.B2(n_7),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

OAI221xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_199),
.B1(n_4),
.B2(n_7),
.C(n_8),
.Y(n_204)
);

AOI31xp33_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_189),
.A3(n_151),
.B(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_4),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_194),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_202),
.A2(n_203),
.B(n_204),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_7),
.B(n_9),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_9),
.Y(n_207)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_207),
.B(n_205),
.CI(n_197),
.CON(n_208),
.SN(n_208)
);


endmodule