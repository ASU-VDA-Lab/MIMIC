module real_jpeg_30947_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_0),
.Y(n_397)
);

BUFx12f_ASAP7_75t_L g488 ( 
.A(n_0),
.Y(n_488)
);

NAND2x1p5_ASAP7_75t_L g177 ( 
.A(n_1),
.B(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_1),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_R g398 ( 
.A(n_1),
.B(n_399),
.Y(n_398)
);

NAND2x1_ASAP7_75t_L g404 ( 
.A(n_1),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_1),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_1),
.B(n_497),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_1),
.B(n_333),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_1),
.B(n_525),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_1),
.B(n_396),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

NAND2x1p5_ASAP7_75t_L g43 ( 
.A(n_2),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_2),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_2),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_2),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_2),
.B(n_155),
.Y(n_154)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_2),
.B(n_224),
.Y(n_223)
);

NAND2x1_ASAP7_75t_L g133 ( 
.A(n_3),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g318 ( 
.A(n_3),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_3),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_3),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_3),
.B(n_437),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_3),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_3),
.B(n_502),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_3),
.B(n_530),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_4),
.A2(n_19),
.B(n_570),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_4),
.B(n_571),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_5),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_5),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_5),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_5),
.B(n_506),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_5),
.B(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_5),
.B(n_540),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_5),
.B(n_544),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_8),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_8),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_8),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_168),
.Y(n_172)
);

NAND2x1_ASAP7_75t_L g183 ( 
.A(n_9),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_9),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_9),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_9),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_9),
.B(n_396),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_10),
.Y(n_571)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_11),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_11),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_12),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_49),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_13),
.B(n_60),
.Y(n_59)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_13),
.B(n_96),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_13),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_13),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_13),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_13),
.B(n_155),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_74),
.Y(n_73)
);

NAND2x1_ASAP7_75t_SL g85 ( 
.A(n_14),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_14),
.B(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_14),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_14),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_14),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_14),
.B(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_15),
.Y(n_226)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_16),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

NAND2x1_ASAP7_75t_L g150 ( 
.A(n_17),
.B(n_44),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_17),
.B(n_189),
.Y(n_188)
);

AND2x4_ASAP7_75t_SL g228 ( 
.A(n_17),
.B(n_88),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_17),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_17),
.B(n_367),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_17),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_17),
.B(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_17),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_105),
.B(n_118),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_21),
.B(n_105),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_80),
.C(n_83),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_22),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_R g22 ( 
.A(n_23),
.B(n_41),
.C(n_57),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_23),
.B(n_42),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.C(n_35),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_24),
.A2(n_25),
.B1(n_30),
.B2(n_161),
.Y(n_266)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_28),
.Y(n_435)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_29),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_31),
.A2(n_152),
.B1(n_161),
.B2(n_162),
.Y(n_151)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_31),
.B(n_154),
.C(n_157),
.Y(n_165)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_33),
.Y(n_212)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_33),
.Y(n_365)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_33),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_35),
.Y(n_265)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_40),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_43),
.A2(n_90),
.B1(n_207),
.B2(n_208),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_45),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_55),
.B2(n_56),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_55),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_56),
.B1(n_95),
.B2(n_100),
.Y(n_94)
);

MAJx2_ASAP7_75t_L g108 ( 
.A(n_47),
.B(n_100),
.C(n_101),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_47),
.Y(n_353)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_48),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_50),
.Y(n_309)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_51),
.A2(n_55),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_51),
.B(n_315),
.C(n_318),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_51),
.B(n_318),
.Y(n_357)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_53),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_54),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_59),
.C(n_63),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_56),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_57),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_67),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_59),
.A2(n_195),
.B1(n_196),
.B2(n_203),
.Y(n_194)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_59),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_59),
.A2(n_63),
.B1(n_110),
.B2(n_203),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_59),
.A2(n_203),
.B1(n_363),
.B2(n_428),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_60),
.Y(n_467)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_61),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_67)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_71),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_77),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_81),
.C(n_82),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_80),
.B(n_83),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_91),
.B2(n_92),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_91),
.C(n_93),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_90),
.B(n_201),
.C(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_101),
.Y(n_93)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_95),
.A2(n_100),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_129),
.Y(n_128)
);

OAI22x1_ASAP7_75t_L g243 ( 
.A1(n_95),
.A2(n_133),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_102),
.B(n_145),
.C(n_211),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_103),
.A2(n_146),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_103),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_117),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_116),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_113),
.A2(n_114),
.B1(n_167),
.B2(n_172),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_113),
.A2(n_114),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_113),
.B(n_167),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_113),
.B(n_221),
.C(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_114),
.A2(n_165),
.B(n_236),
.C(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_291),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_283),
.B(n_289),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_271),
.B(n_282),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_250),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_124),
.B(n_250),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_191),
.B(n_249),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_125),
.B(n_381),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_163),
.C(n_173),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_126),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.C(n_151),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_127),
.A2(n_128),
.B1(n_137),
.B2(n_138),
.Y(n_375)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2x1_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_130),
.B(n_133),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_130),
.Y(n_245)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_132),
.Y(n_504)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.C(n_150),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2x2_ASAP7_75t_L g320 ( 
.A(n_140),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_141),
.A2(n_342),
.B1(n_344),
.B2(n_345),
.Y(n_341)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_142),
.Y(n_546)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_144),
.Y(n_317)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_146),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_149),
.Y(n_209)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_150),
.Y(n_322)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_151),
.Y(n_374)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_160),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g358 ( 
.A(n_153),
.B(n_359),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_153),
.A2(n_154),
.B1(n_359),
.B2(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_157),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_157),
.A2(n_160),
.B1(n_227),
.B2(n_228),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_157),
.B(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_157),
.B(n_470),
.Y(n_494)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_159),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_160),
.B(n_222),
.C(n_227),
.Y(n_221)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_164),
.B(n_173),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_171),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_182),
.C(n_186),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2x1_ASAP7_75t_L g324 ( 
.A(n_175),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_179),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g352 ( 
.A(n_177),
.B(n_179),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_178),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_179),
.B(n_201),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_179),
.A2(n_202),
.B(n_475),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_179),
.B(n_476),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_183),
.A2(n_188),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_183),
.Y(n_326)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_185),
.Y(n_499)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_188),
.Y(n_327)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_190),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_217),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_217),
.Y(n_249)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_193),
.B(n_218),
.Y(n_381)
);

XOR2x2_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_204),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_194),
.B(n_205),
.C(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_261)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_201),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_201),
.Y(n_476)
);

XNOR2x1_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_203),
.B(n_363),
.C(n_366),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_210),
.B2(n_216),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

INVxp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_238),
.B1(n_239),
.B2(n_248),
.Y(n_218)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

XNOR2x1_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_235),
.Y(n_219)
);

INVxp33_ASAP7_75t_SL g253 ( 
.A(n_220),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_229),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_223),
.Y(n_310)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_226),
.Y(n_541)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx8_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_253),
.C(n_254),
.Y(n_252)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.C(n_246),
.Y(n_239)
);

XOR2x2_ASAP7_75t_L g346 ( 
.A(n_240),
.B(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_241),
.B(n_308),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_243),
.B(n_246),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_262),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_255),
.C(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_260),
.C(n_261),
.Y(n_281)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_269),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_267),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_269),
.C(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_281),
.C(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVxp33_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_287),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_287),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_449),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_386),
.B(n_445),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_298),
.B(n_450),
.C(n_452),
.Y(n_449)
);

AOI22x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_348),
.B1(n_379),
.B2(n_382),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_300),
.B(n_349),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

MAJx2_ASAP7_75t_L g383 ( 
.A(n_301),
.B(n_384),
.C(n_385),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_346),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_323),
.C(n_328),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_305),
.B(n_323),
.C(n_328),
.Y(n_384)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_306),
.B(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_314),
.C(n_320),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_307),
.B(n_320),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.C(n_311),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_311),
.B(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_314),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_315),
.B(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_324),
.B(n_329),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_334),
.C(n_341),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_331),
.B1(n_334),
.B2(n_335),
.Y(n_371)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_371),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_341),
.A2(n_395),
.B(n_398),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_345),
.Y(n_399)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_346),
.Y(n_385)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_372),
.C(n_376),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.C(n_369),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_370),
.Y(n_390)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

XOR2x2_ASAP7_75t_SL g389 ( 
.A(n_355),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.C(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_358),
.B(n_362),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_363),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_366),
.B(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_373),
.B(n_377),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_380),
.B(n_383),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_380),
.B(n_383),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_413),
.B(n_444),
.Y(n_386)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_387),
.B(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_411),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_388),
.B(n_411),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.C(n_408),
.Y(n_388)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_408),
.Y(n_415)
);

MAJx2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.C(n_400),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_392),
.B(n_419),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_394),
.B(n_400),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_403),
.C(n_404),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g462 ( 
.A(n_402),
.B(n_463),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_403),
.B(n_404),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XNOR2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_414),
.B(n_416),
.Y(n_451)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_424),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_418),
.B(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_425),
.Y(n_455)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_429),
.C(n_432),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_426),
.B(n_459),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_429),
.A2(n_430),
.B1(n_432),
.B2(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_432),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_436),
.C(n_439),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_433),
.A2(n_434),
.B1(n_439),
.B2(n_440),
.Y(n_560)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_436),
.B(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx5_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B(n_448),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_453),
.A2(n_477),
.B(n_568),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.Y(n_453)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_454),
.Y(n_569)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_457),
.B(n_569),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_461),
.C(n_464),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_458),
.B(n_564),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_461),
.A2(n_462),
.B1(n_464),
.B2(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_464),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.C(n_474),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_465),
.A2(n_466),
.B1(n_474),
.B2(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_468),
.B(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g556 ( 
.A(n_474),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_562),
.B(n_567),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_479),
.A2(n_551),
.B(n_561),
.Y(n_478)
);

AOI21x1_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_521),
.B(n_550),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_513),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_495),
.B1(n_511),
.B2(n_512),
.Y(n_481)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_482),
.Y(n_511)
);

AOI221xp5_ASAP7_75t_L g550 ( 
.A1(n_482),
.A2(n_495),
.B1(n_511),
.B2(n_512),
.C(n_513),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_484),
.B1(n_493),
.B2(n_494),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_483),
.B(n_494),
.C(n_512),
.Y(n_552)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_489),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_489),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_487),
.Y(n_485)
);

INVx8_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx8_ASAP7_75t_L g531 ( 
.A(n_488),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx6_ASAP7_75t_L g528 ( 
.A(n_492),
.Y(n_528)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_500),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_496),
.B(n_501),
.C(n_505),
.Y(n_558)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_505),
.B1(n_509),
.B2(n_510),
.Y(n_500)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_505),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_507),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_516),
.C(n_517),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_514),
.A2(n_515),
.B1(n_533),
.B2(n_534),
.Y(n_532)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_516),
.A2(n_517),
.B1(n_518),
.B2(n_535),
.Y(n_534)
);

CKINVDCx12_ASAP7_75t_R g535 ( 
.A(n_516),
.Y(n_535)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_522),
.A2(n_536),
.B(n_549),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_532),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_523),
.B(n_532),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_529),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_529),
.Y(n_538)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_537),
.A2(n_542),
.B(n_548),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_538),
.B(n_539),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_538),
.B(n_539),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_547),
.Y(n_542)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_553),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_552),
.B(n_553),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_554),
.B(n_557),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_558),
.C(n_559),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_559),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_563),
.B(n_566),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_SL g567 ( 
.A(n_563),
.B(n_566),
.Y(n_567)
);


endmodule