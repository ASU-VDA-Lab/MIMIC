module fake_jpeg_19635_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx4_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_20),
.B(n_27),
.C(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_28),
.B(n_16),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_16),
.B1(n_24),
.B2(n_31),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_48),
.B1(n_54),
.B2(n_35),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_46),
.B(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_39),
.B1(n_24),
.B2(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_28),
.B1(n_19),
.B2(n_18),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_37),
.C(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_51),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_60),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_63),
.B(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_72),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_66),
.B(n_73),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_71),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_37),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_53),
.C(n_44),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_34),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_40),
.B(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_36),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_31),
.B1(n_40),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_52),
.B1(n_20),
.B2(n_25),
.Y(n_102)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_37),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_32),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_52),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_105),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_77),
.B(n_67),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_106),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_94),
.B1(n_80),
.B2(n_64),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_29),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_75),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_65),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_111),
.B(n_112),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_127),
.B1(n_95),
.B2(n_93),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_20),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_97),
.B(n_94),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_125),
.B(n_129),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_61),
.C(n_59),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_87),
.C(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_120),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_83),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_68),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_60),
.B(n_68),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_105),
.A2(n_84),
.B1(n_82),
.B2(n_62),
.Y(n_127)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_66),
.B(n_71),
.C(n_65),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_133),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_131),
.B(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_120),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_112),
.B1(n_132),
.B2(n_122),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_139),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_99),
.B1(n_128),
.B2(n_110),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_144),
.B1(n_146),
.B2(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_154),
.Y(n_161)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_109),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_92),
.B1(n_107),
.B2(n_103),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_113),
.A2(n_87),
.B1(n_108),
.B2(n_30),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_157),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_156),
.C(n_115),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_116),
.B(n_23),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_151),
.B(n_134),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_152),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_129),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_19),
.C(n_26),
.Y(n_156)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_26),
.A3(n_22),
.B1(n_20),
.B2(n_25),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_172),
.C(n_156),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_115),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_168),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_166),
.B1(n_146),
.B2(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_122),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_167),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_142),
.A2(n_123),
.B1(n_126),
.B2(n_118),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_22),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_125),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_174),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_118),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_137),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_176),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_126),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_181),
.C(n_185),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_187),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_144),
.C(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_188),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_153),
.C(n_145),
.Y(n_185)
);

OAI322xp33_ASAP7_75t_L g186 ( 
.A1(n_168),
.A2(n_157),
.A3(n_135),
.B1(n_152),
.B2(n_21),
.C1(n_23),
.C2(n_13),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_186),
.B(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_135),
.B1(n_2),
.B2(n_3),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_21),
.C(n_13),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_172),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_196),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_195),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_175),
.C(n_169),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_194),
.A2(n_1),
.B(n_4),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_177),
.B(n_174),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_200),
.Y(n_208)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_175),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_21),
.C(n_2),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_5),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_197),
.A2(n_166),
.B1(n_181),
.B2(n_185),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_206),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_190),
.B1(n_11),
.B2(n_3),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_196),
.B1(n_190),
.B2(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_5),
.C(n_7),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_210),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_208),
.B(n_209),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.Y(n_220)
);

OA21x2_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_1),
.B(n_4),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_215),
.B(n_7),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_202),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_7),
.C(n_8),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_219),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_9),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_221),
.B(n_222),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_212),
.B(n_214),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_217),
.B(n_8),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_226),
.B(n_227),
.C(n_223),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_9),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_229),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_9),
.Y(n_231)
);


endmodule