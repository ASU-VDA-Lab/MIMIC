module real_jpeg_23509_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_221;
wire n_300;
wire n_292;
wire n_288;
wire n_249;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_299;
wire n_105;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_293;
wire n_275;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_240;
wire n_55;
wire n_185;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_1),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_300),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_2),
.B(n_301),
.Y(n_300)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_3),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g301 ( 
.A(n_5),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_6),
.A2(n_10),
.B1(n_22),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_6),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_6),
.A2(n_52),
.B1(n_81),
.B2(n_82),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_30),
.C(n_32),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_6),
.B(n_29),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_6),
.B(n_59),
.C(n_62),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_6),
.B(n_78),
.C(n_81),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_6),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_6),
.B(n_108),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_6),
.B(n_71),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_24),
.B1(n_26),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_8),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_68),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_8),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_20),
.B1(n_31),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_20),
.B1(n_62),
.B2(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_20),
.B1(n_81),
.B2(n_82),
.Y(n_94)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_41),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_11),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_11),
.A2(n_41),
.B1(n_81),
.B2(n_82),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_13),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_44),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_42),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_37),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_27),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_19),
.A2(n_29),
.B1(n_35),
.B2(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_24),
.B1(n_30),
.B2(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_23),
.B(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_28),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_29),
.A2(n_35),
.B1(n_51),
.B2(n_66),
.Y(n_65)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_29)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_32),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_32),
.B(n_227),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_38),
.B(n_46),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_49),
.B(n_50),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_84),
.B(n_299),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_47),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_47),
.B(n_297),
.Y(n_298)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.CI(n_64),
.CON(n_47),
.SN(n_47)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_49),
.A2(n_50),
.B(n_67),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_56),
.A2(n_61),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_71),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_57),
.B(n_113),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_61),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OA22x2_ASAP7_75t_SL g61 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_61),
.A2(n_122),
.B(n_123),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_61),
.A2(n_112),
.B(n_123),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_63),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_62),
.B(n_240),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.C(n_72),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_65),
.B(n_131),
.C(n_138),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_65),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_65),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_65),
.A2(n_138),
.B1(n_139),
.B2(n_152),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_65),
.A2(n_110),
.B1(n_152),
.B2(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_65),
.B(n_110),
.C(n_190),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_69),
.A2(n_72),
.B1(n_120),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_69),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_72),
.A2(n_120),
.B1(n_121),
.B2(n_124),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_72),
.B(n_116),
.C(n_121),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_83),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_74),
.B(n_99),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_76),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_76),
.A2(n_99),
.B1(n_108),
.B2(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_80),
.A2(n_98),
.B(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_81),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_81),
.B(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_296),
.B(n_298),
.Y(n_84)
);

OAI211xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_140),
.B(n_154),
.C(n_295),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_125),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_87),
.B(n_125),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_103),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_88),
.B(n_105),
.C(n_114),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_95),
.B(n_100),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_89),
.A2(n_100),
.B1(n_101),
.B2(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_89),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_89),
.A2(n_96),
.B1(n_128),
.B2(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_91),
.B(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_92),
.A2(n_94),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_92),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_93),
.A2(n_133),
.B(n_167),
.Y(n_166)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_96),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_114),
.B2(n_115),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_106),
.B(n_110),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.Y(n_105)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_110),
.B(n_211),
.C(n_213),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_110),
.A2(n_201),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_117),
.B1(n_148),
.B2(n_153),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_116),
.B(n_138),
.C(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_116),
.A2(n_117),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_116),
.A2(n_117),
.B1(n_172),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_164),
.C(n_172),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_117),
.B(n_144),
.C(n_148),
.Y(n_297)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_121),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.C(n_130),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_126),
.B(n_129),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_132),
.Y(n_286)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_134),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_135),
.A2(n_136),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_135),
.A2(n_136),
.B1(n_224),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_136),
.B(n_218),
.C(n_224),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_195),
.C(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_138),
.A2(n_139),
.B1(n_186),
.B2(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_138),
.A2(n_139),
.B1(n_170),
.B2(n_183),
.Y(n_263)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_139),
.B(n_170),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_SL g154 ( 
.A(n_141),
.B(n_155),
.C(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_142),
.B(n_143),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_176),
.B(n_294),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_174),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_158),
.B(n_174),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_159),
.B(n_161),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_163),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_164),
.A2(n_165),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_170),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_166),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_197),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_170),
.A2(n_183),
.B1(n_239),
.B2(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_170),
.B(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_289),
.B(n_293),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_214),
.B(n_275),
.C(n_288),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_203),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_179),
.B(n_203),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_189),
.B2(n_202),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_182),
.B(n_188),
.C(n_202),
.Y(n_276)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_185),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_191),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_194),
.A2(n_195),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_249),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_195),
.B(n_249),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.C(n_210),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_204),
.A2(n_205),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_209),
.B(n_210),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_213),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_211),
.B(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_213),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_274),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_233),
.B(n_273),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_230),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_217),
.B(n_230),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_218),
.A2(n_219),
.B1(n_269),
.B2(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_223),
.B(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_266),
.B(n_272),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_260),
.B(n_265),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_252),
.B(n_259),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_242),
.B(n_251),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_239),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_248),
.B(n_250),
.Y(n_242)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_254),
.Y(n_259)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_257),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_287),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_284),
.B2(n_285),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_285),
.C(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);


endmodule