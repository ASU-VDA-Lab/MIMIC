module fake_jpeg_26130_n_102 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_102);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_4),
.B(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_28),
.Y(n_34)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_16),
.B(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_18),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_29),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_19),
.B1(n_16),
.B2(n_21),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_19),
.B1(n_14),
.B2(n_12),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_27),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_49),
.B1(n_34),
.B2(n_13),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_20),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_47),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_12),
.A3(n_14),
.B1(n_13),
.B2(n_15),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_34),
.Y(n_53)
);

NAND2x1p5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_30),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_60),
.B(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_5),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_15),
.B1(n_12),
.B2(n_27),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_39),
.C(n_24),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_39),
.C(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_13),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_1),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_20),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_65),
.Y(n_76)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_69),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_56),
.B1(n_54),
.B2(n_50),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_58),
.B1(n_39),
.B2(n_37),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_60),
.A2(n_3),
.B(n_4),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_77),
.B1(n_69),
.B2(n_6),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_75),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_24),
.C(n_25),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_63),
.A2(n_22),
.B(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_79),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_70),
.B1(n_71),
.B2(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_67),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_6),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_85),
.A2(n_86),
.B(n_9),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_78),
.B(n_76),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_89),
.B(n_91),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_77),
.B(n_8),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_94),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_81),
.B(n_10),
.Y(n_94)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_3),
.C(n_36),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_36),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g99 ( 
.A(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_36),
.Y(n_98)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_22),
.A3(n_24),
.B1(n_25),
.B2(n_32),
.C1(n_36),
.C2(n_96),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_32),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_99),
.Y(n_102)
);


endmodule