module fake_jpeg_1622_n_649 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_649);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_649;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_539;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_9),
.B(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_58),
.Y(n_160)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_59),
.Y(n_182)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_25),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_61),
.B(n_80),
.Y(n_144)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_64),
.Y(n_154)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_68),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_76),
.Y(n_133)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_70),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_72),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_73),
.Y(n_159)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_39),
.B(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_77),
.Y(n_184)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_1),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_82),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_39),
.B(n_56),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_83),
.B(n_56),
.Y(n_146)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_85),
.B(n_7),
.Y(n_175)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_87),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_26),
.B(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_88),
.B(n_98),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_92),
.Y(n_181)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_93),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_95),
.Y(n_204)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_26),
.B(n_2),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_33),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_100),
.A2(n_41),
.B1(n_126),
.B2(n_127),
.Y(n_208)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_20),
.B(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_105),
.B(n_106),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g106 ( 
.A1(n_36),
.A2(n_5),
.B(n_7),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

BUFx24_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_111),
.Y(n_221)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_117),
.Y(n_135)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_113),
.Y(n_231)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_31),
.Y(n_114)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_20),
.B(n_5),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_115),
.B(n_10),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_116),
.Y(n_233)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_36),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_37),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_123),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_119),
.Y(n_229)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_120),
.B(n_122),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_30),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_130),
.Y(n_142)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_126),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_52),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_128),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx2_ASAP7_75t_R g202 ( 
.A(n_129),
.Y(n_202)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_54),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_30),
.Y(n_132)
);

CKINVDCx12_ASAP7_75t_R g234 ( 
.A(n_132),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_69),
.A2(n_40),
.B1(n_54),
.B2(n_34),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_140),
.A2(n_171),
.B1(n_228),
.B2(n_178),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_145),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_146),
.B(n_147),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_61),
.B(n_32),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_80),
.A2(n_32),
.B1(n_51),
.B2(n_50),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_152),
.A2(n_168),
.B1(n_208),
.B2(n_217),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_105),
.B(n_27),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_163),
.B(n_164),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_27),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_88),
.A2(n_41),
.B1(n_54),
.B2(n_34),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_167),
.A2(n_215),
.B1(n_203),
.B2(n_168),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_70),
.A2(n_21),
.B1(n_50),
.B2(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_98),
.B(n_51),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_183),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_67),
.A2(n_45),
.B1(n_40),
.B2(n_38),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_178),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_68),
.A2(n_38),
.B1(n_44),
.B2(n_35),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_90),
.B(n_35),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_110),
.A2(n_21),
.B(n_40),
.C(n_45),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g295 ( 
.A1(n_190),
.A2(n_200),
.B(n_234),
.C(n_217),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_84),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_191),
.B(n_194),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_87),
.B(n_45),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_192),
.B(n_209),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_124),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_131),
.B(n_8),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_196),
.B(n_197),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_131),
.B(n_8),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_79),
.B(n_8),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_199),
.B(n_210),
.Y(n_319)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_82),
.A2(n_37),
.B(n_41),
.C(n_11),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_89),
.B(n_9),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_79),
.B(n_10),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_212),
.B(n_213),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_10),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_116),
.B(n_11),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_SL g316 ( 
.A1(n_214),
.A2(n_219),
.B(n_207),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_99),
.A2(n_37),
.B1(n_12),
.B2(n_13),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_94),
.A2(n_37),
.B1(n_12),
.B2(n_13),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_218),
.B1(n_226),
.B2(n_134),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_97),
.A2(n_129),
.B1(n_121),
.B2(n_119),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_103),
.A2(n_37),
.B1(n_12),
.B2(n_13),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_130),
.B(n_11),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_82),
.A2(n_37),
.B1(n_15),
.B2(n_17),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_222),
.A2(n_224),
.B1(n_230),
.B2(n_177),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_80),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_228),
.B1(n_140),
.B2(n_232),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_69),
.A2(n_17),
.B1(n_80),
.B2(n_61),
.Y(n_224)
);

OA22x2_ASAP7_75t_L g227 ( 
.A1(n_111),
.A2(n_17),
.B1(n_113),
.B2(n_108),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_227),
.A2(n_190),
.B(n_230),
.C(n_134),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_100),
.A2(n_69),
.B1(n_61),
.B2(n_85),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_L g230 ( 
.A1(n_111),
.A2(n_109),
.B1(n_84),
.B2(n_70),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_76),
.B(n_61),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_133),
.Y(n_244)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_142),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_236),
.B(n_253),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_237),
.Y(n_359)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_239),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_161),
.A2(n_200),
.B1(n_204),
.B2(n_137),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_240),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_241),
.A2(n_250),
.B1(n_312),
.B2(n_244),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_242),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_361)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_244),
.B(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_181),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_245),
.B(n_249),
.Y(n_331)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_246),
.Y(n_372)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_227),
.A2(n_171),
.B1(n_223),
.B2(n_136),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_170),
.B(n_135),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_144),
.A2(n_227),
.B1(n_172),
.B2(n_231),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_139),
.B(n_182),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_255),
.B(n_265),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_203),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_257),
.B(n_294),
.Y(n_345)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_259),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_205),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_260),
.B(n_271),
.Y(n_328)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_261),
.Y(n_358)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_211),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_263),
.Y(n_339)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_139),
.B(n_204),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_157),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_267),
.B(n_303),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_201),
.B(n_161),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_268),
.B(n_285),
.C(n_296),
.Y(n_326)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_205),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_270),
.B(n_273),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_201),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_206),
.A2(n_155),
.B1(n_201),
.B2(n_165),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_272),
.A2(n_277),
.B1(n_293),
.B2(n_301),
.Y(n_370)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_275),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_187),
.A2(n_188),
.B1(n_155),
.B2(n_198),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_141),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_287),
.Y(n_347)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_279),
.Y(n_364)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_154),
.Y(n_280)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_280),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_154),
.B(n_157),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_281),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_176),
.B(n_184),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_282),
.Y(n_362)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_283),
.Y(n_383)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_176),
.Y(n_284)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_284),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_184),
.B(n_195),
.C(n_151),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_226),
.A2(n_179),
.B1(n_162),
.B2(n_198),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_286),
.A2(n_276),
.B1(n_294),
.B2(n_265),
.Y(n_353)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_151),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_162),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_289),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_179),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_156),
.Y(n_290)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_290),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_150),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_292),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_187),
.A2(n_188),
.B1(n_150),
.B2(n_165),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_226),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_295),
.A2(n_313),
.B(n_256),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g296 ( 
.A(n_156),
.B(n_186),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_195),
.A2(n_159),
.B1(n_153),
.B2(n_186),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_298),
.A2(n_315),
.B1(n_318),
.B2(n_321),
.Y(n_338)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_299),
.B(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_185),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_305),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_143),
.A2(n_158),
.B1(n_173),
.B2(n_153),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_143),
.B(n_159),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_173),
.B(n_229),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_149),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_306),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_148),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_149),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_202),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_307),
.Y(n_367)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_308),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_229),
.B(n_233),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_229),
.B(n_189),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_158),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_311),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_SL g313 ( 
.A(n_202),
.B(n_189),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_177),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_314),
.Y(n_380)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_193),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_207),
.B(n_193),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_317),
.B(n_322),
.Y(n_354)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_166),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_166),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_174),
.B(n_209),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_174),
.B(n_209),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_323),
.B(n_238),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_295),
.A2(n_242),
.B(n_302),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_330),
.A2(n_335),
.B(n_347),
.Y(n_421)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_322),
.A2(n_323),
.B(n_236),
.C(n_267),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_334),
.B(n_360),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_276),
.A2(n_312),
.B1(n_256),
.B2(n_266),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_337),
.A2(n_353),
.B1(n_376),
.B2(n_382),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_301),
.A2(n_241),
.B1(n_251),
.B2(n_293),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_244),
.A2(n_277),
.B1(n_320),
.B2(n_291),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

AOI32xp33_ASAP7_75t_L g349 ( 
.A1(n_313),
.A2(n_319),
.A3(n_253),
.B1(n_247),
.B2(n_268),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_349),
.B(n_282),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_352),
.B(n_356),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_257),
.Y(n_398)
);

AO22x1_ASAP7_75t_SL g356 ( 
.A1(n_282),
.A2(n_281),
.B1(n_266),
.B2(n_248),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g363 ( 
.A1(n_297),
.A2(n_317),
.B(n_269),
.C(n_255),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_363),
.B(n_375),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_283),
.A2(n_274),
.B1(n_262),
.B2(n_261),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_368),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_282),
.A2(n_303),
.B(n_309),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_369),
.A2(n_299),
.B(n_304),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_285),
.B(n_281),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_310),
.A2(n_296),
.B1(n_243),
.B2(n_235),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_296),
.A2(n_258),
.B1(n_292),
.B2(n_311),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_387),
.B(n_399),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_280),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_401),
.Y(n_439)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_389),
.Y(n_435)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_284),
.Y(n_391)
);

XNOR2x1_ASAP7_75t_L g463 ( 
.A(n_391),
.B(n_422),
.Y(n_463)
);

OR2x2_ASAP7_75t_SL g392 ( 
.A(n_362),
.B(n_246),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_392),
.A2(n_419),
.B(n_325),
.Y(n_457)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_382),
.Y(n_396)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_397),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_398),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_367),
.B(n_315),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_352),
.A2(n_308),
.B1(n_264),
.B2(n_275),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_400),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_367),
.B(n_279),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_361),
.A2(n_263),
.B1(n_337),
.B2(n_365),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_402),
.A2(n_408),
.B1(n_414),
.B2(n_416),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_361),
.A2(n_330),
.B1(n_355),
.B2(n_354),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_384),
.A2(n_359),
.B1(n_333),
.B2(n_370),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_384),
.A2(n_359),
.B1(n_333),
.B2(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_406),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_353),
.A2(n_371),
.B1(n_363),
.B2(n_369),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_345),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_409),
.B(n_429),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_357),
.A2(n_371),
.B1(n_362),
.B2(n_334),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_410),
.A2(n_415),
.B1(n_418),
.B2(n_341),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_360),
.B(n_375),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_412),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_331),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_350),
.B1(n_376),
.B2(n_346),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_357),
.A2(n_350),
.B1(n_346),
.B2(n_326),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_328),
.A2(n_356),
.B1(n_326),
.B2(n_349),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_417),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_326),
.A2(n_356),
.B1(n_329),
.B2(n_338),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_351),
.A2(n_336),
.B(n_329),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_356),
.A2(n_327),
.B1(n_335),
.B2(n_366),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_420),
.A2(n_364),
.B1(n_372),
.B2(n_339),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_421),
.A2(n_423),
.B(n_372),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_331),
.B(n_347),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_345),
.A2(n_377),
.B(n_383),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_424),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_378),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_427),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_380),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_385),
.B(n_373),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_431),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_345),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_343),
.B(n_377),
.C(n_383),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g432 ( 
.A(n_377),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_432),
.B(n_341),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_373),
.Y(n_436)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_436),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_396),
.A2(n_366),
.B1(n_378),
.B2(n_379),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx13_ASAP7_75t_L g438 ( 
.A(n_392),
.Y(n_438)
);

INVx11_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_418),
.B(n_379),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_444),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_446),
.B(n_447),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_425),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_448),
.A2(n_457),
.B(n_468),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_427),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_449),
.B(n_450),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_358),
.Y(n_450)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_394),
.Y(n_455)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_404),
.A2(n_342),
.B1(n_340),
.B2(n_325),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_456),
.A2(n_386),
.B1(n_441),
.B2(n_454),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_412),
.B(n_358),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_458),
.B(n_459),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_422),
.B(n_340),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_398),
.B(n_342),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_461),
.B(n_423),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_428),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_462),
.B(n_388),
.Y(n_480)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_389),
.Y(n_465)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

CKINVDCx12_ASAP7_75t_R g467 ( 
.A(n_392),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_467),
.Y(n_475)
);

INVx13_ASAP7_75t_L g469 ( 
.A(n_409),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g472 ( 
.A(n_469),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_470),
.A2(n_400),
.B1(n_405),
.B2(n_429),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_426),
.A2(n_339),
.B1(n_364),
.B2(n_413),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_471),
.A2(n_430),
.B(n_423),
.Y(n_501)
);

OAI221xp5_ASAP7_75t_L g473 ( 
.A1(n_448),
.A2(n_407),
.B1(n_416),
.B2(n_387),
.C(n_395),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_491),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_463),
.B(n_415),
.C(n_391),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_486),
.C(n_489),
.Y(n_520)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_435),
.Y(n_479)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_479),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_480),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_451),
.B(n_411),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_493),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_492),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_463),
.B(n_403),
.C(n_407),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_487),
.A2(n_436),
.B1(n_445),
.B2(n_456),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_414),
.C(n_421),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g492 ( 
.A1(n_468),
.A2(n_393),
.B(n_420),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_464),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_433),
.A2(n_457),
.B(n_466),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g538 ( 
.A1(n_495),
.A2(n_505),
.B(n_438),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_434),
.A2(n_402),
.B1(n_393),
.B2(n_386),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_497),
.A2(n_507),
.B1(n_462),
.B2(n_447),
.Y(n_517)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_498),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_440),
.B(n_466),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_499),
.B(n_503),
.C(n_504),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_451),
.B(n_395),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_502),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g513 ( 
.A(n_501),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_450),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_410),
.C(n_393),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_408),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_457),
.A2(n_397),
.B(n_432),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_465),
.Y(n_506)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_506),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_434),
.A2(n_401),
.B1(n_399),
.B2(n_417),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_449),
.B(n_431),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_499),
.Y(n_523)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_442),
.Y(n_509)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_509),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_484),
.A2(n_444),
.B1(n_452),
.B2(n_441),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_519),
.B(n_522),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_436),
.Y(n_522)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_483),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_526),
.B1(n_530),
.B2(n_536),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_483),
.B(n_464),
.Y(n_525)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_525),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_490),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_507),
.Y(n_527)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_490),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_493),
.B(n_439),
.Y(n_531)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_531),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_494),
.A2(n_452),
.B(n_467),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_532),
.A2(n_535),
.B(n_537),
.Y(n_557)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_482),
.Y(n_533)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_533),
.Y(n_547)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_534),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_494),
.A2(n_505),
.B(n_475),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_492),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_538),
.A2(n_540),
.B(n_484),
.Y(n_563)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_478),
.Y(n_539)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_539),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_497),
.A2(n_470),
.B1(n_439),
.B2(n_444),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_492),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_541),
.B(n_542),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_491),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_474),
.B(n_458),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_543),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_474),
.B(n_446),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_544),
.B(n_502),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_489),
.C(n_477),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_549),
.B(n_554),
.C(n_559),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_503),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_551),
.B(n_561),
.Y(n_579)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_552),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_545),
.B(n_486),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_556),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_504),
.C(n_444),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_523),
.B(n_473),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_520),
.B(n_488),
.C(n_510),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_520),
.B(n_510),
.C(n_460),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_560),
.B(n_572),
.C(n_573),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_516),
.B(n_495),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_516),
.B(n_460),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g594 ( 
.A(n_562),
.B(n_565),
.Y(n_594)
);

AO21x1_ASAP7_75t_L g581 ( 
.A1(n_563),
.A2(n_515),
.B(n_535),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_515),
.A2(n_475),
.B(n_501),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g586 ( 
.A1(n_564),
.A2(n_515),
.B(n_522),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_517),
.B(n_521),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_538),
.B(n_472),
.C(n_487),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_538),
.B(n_472),
.C(n_506),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_514),
.B(n_453),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_511),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_568),
.A2(n_527),
.B1(n_511),
.B2(n_524),
.Y(n_577)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_577),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_573),
.Y(n_578)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_578),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_550),
.A2(n_542),
.B1(n_530),
.B2(n_526),
.Y(n_580)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_569),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_582),
.B(n_585),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_555),
.A2(n_521),
.B1(n_540),
.B2(n_532),
.Y(n_585)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_571),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_589),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_588),
.B(n_509),
.Y(n_607)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_567),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_551),
.B(n_522),
.C(n_537),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_590),
.B(n_593),
.C(n_595),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_566),
.A2(n_525),
.B1(n_531),
.B2(n_476),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_591),
.B(n_597),
.Y(n_606)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_570),
.A2(n_519),
.B1(n_541),
.B2(n_536),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_554),
.B(n_560),
.C(n_559),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_553),
.B(n_513),
.C(n_544),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_557),
.A2(n_513),
.B(n_496),
.Y(n_596)
);

OAI321xp33_ASAP7_75t_L g599 ( 
.A1(n_596),
.A2(n_564),
.A3(n_570),
.B1(n_557),
.B2(n_563),
.C(n_548),
.Y(n_599)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_599),
.A2(n_585),
.B(n_586),
.Y(n_616)
);

AOI31xp33_ASAP7_75t_L g603 ( 
.A1(n_576),
.A2(n_549),
.A3(n_546),
.B(n_556),
.Y(n_603)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_603),
.Y(n_617)
);

A2O1A1O1Ixp25_ASAP7_75t_L g604 ( 
.A1(n_595),
.A2(n_561),
.B(n_565),
.C(n_496),
.D(n_562),
.Y(n_604)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_604),
.A2(n_596),
.B(n_581),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_543),
.C(n_547),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_605),
.B(n_608),
.C(n_612),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_607),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_583),
.C(n_579),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_580),
.A2(n_471),
.B1(n_512),
.B2(n_529),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_610),
.A2(n_597),
.B1(n_592),
.B2(n_518),
.Y(n_618)
);

BUFx24_ASAP7_75t_SL g611 ( 
.A(n_589),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_611),
.B(n_584),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_575),
.B(n_583),
.C(n_579),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_578),
.B(n_547),
.C(n_529),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_613),
.B(n_614),
.C(n_443),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_590),
.B(n_528),
.C(n_518),
.Y(n_614)
);

AOI21x1_ASAP7_75t_SL g627 ( 
.A1(n_615),
.A2(n_616),
.B(n_621),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_618),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g619 ( 
.A1(n_609),
.A2(n_594),
.B1(n_584),
.B2(n_528),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_619),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_620),
.B(n_624),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_600),
.A2(n_594),
.B(n_498),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_606),
.A2(n_479),
.B1(n_533),
.B2(n_453),
.Y(n_622)
);

INVxp33_ASAP7_75t_L g630 ( 
.A(n_622),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_602),
.B(n_482),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_626),
.B(n_602),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_629),
.B(n_633),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_625),
.B(n_605),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_SL g634 ( 
.A(n_623),
.B(n_601),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_634),
.B(n_635),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_625),
.B(n_608),
.C(n_612),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_627),
.A2(n_617),
.B(n_616),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_636),
.A2(n_638),
.B(n_639),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_628),
.B(n_624),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g642 ( 
.A(n_637),
.B(n_626),
.Y(n_642)
);

AOI31xp67_ASAP7_75t_L g638 ( 
.A1(n_630),
.A2(n_598),
.A3(n_614),
.B(n_613),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_631),
.B(n_620),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_642),
.A2(n_621),
.B(n_619),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_641),
.B(n_631),
.Y(n_644)
);

AO21x2_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_640),
.B(n_615),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_645),
.B(n_646),
.C(n_643),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_SL g648 ( 
.A1(n_647),
.A2(n_632),
.B1(n_622),
.B2(n_610),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_648),
.Y(n_649)
);


endmodule