module fake_aes_10883_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
AOI22xp33_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_6), .B(n_3), .Y(n_7) );
AOI221xp5_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_3), .B1(n_4), .B2(n_0), .C(n_2), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_4), .Y(n_9) );
NOR2xp33_ASAP7_75t_L g10 ( .A(n_9), .B(n_8), .Y(n_10) );
NOR3xp33_ASAP7_75t_SL g11 ( .A(n_9), .B(n_1), .C(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
AOI222xp33_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_2), .C1(n_11), .C2(n_10), .Y(n_13) );
endmodule