module fake_jpeg_14109_n_569 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_569);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_569;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_57),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_58),
.B(n_64),
.Y(n_125)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_62),
.Y(n_173)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_38),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_38),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_75),
.Y(n_129)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_18),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_86),
.Y(n_131)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

BUFx16f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_79),
.Y(n_177)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_81),
.Y(n_156)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_82),
.Y(n_175)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_84),
.Y(n_152)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_85),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_19),
.B(n_15),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_19),
.B(n_15),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_89),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_25),
.B(n_15),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_92),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_25),
.B(n_1),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_1),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_99),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_32),
.Y(n_97)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_27),
.Y(n_98)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_31),
.B(n_2),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_110),
.Y(n_178)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_40),
.Y(n_111)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

BUFx24_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g233 ( 
.A(n_117),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_53),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_123),
.B(n_128),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_160),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g128 ( 
.A(n_83),
.B(n_30),
.Y(n_128)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_34),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_139),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_34),
.Y(n_139)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_58),
.A2(n_45),
.B(n_46),
.Y(n_144)
);

NAND2x1_ASAP7_75t_SL g229 ( 
.A(n_144),
.B(n_51),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_79),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_145),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_154),
.Y(n_197)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

NOR2x1_ASAP7_75t_R g154 ( 
.A(n_64),
.B(n_30),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_75),
.B(n_30),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_78),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_162),
.B(n_179),
.Y(n_203)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_60),
.B(n_39),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_169),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_93),
.B(n_39),
.Y(n_169)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_56),
.B(n_47),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_72),
.B(n_47),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_42),
.Y(n_212)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_127),
.Y(n_185)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_185),
.Y(n_296)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_187),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_118),
.A2(n_69),
.B1(n_17),
.B2(n_41),
.Y(n_189)
);

OAI22x1_ASAP7_75t_SL g288 ( 
.A1(n_189),
.A2(n_221),
.B1(n_243),
.B2(n_152),
.Y(n_288)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_135),
.Y(n_192)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_193),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_131),
.B(n_46),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_194),
.B(n_206),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_100),
.B1(n_57),
.B2(n_76),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_198),
.A2(n_208),
.B1(n_121),
.B2(n_116),
.Y(n_280)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_132),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_199),
.Y(n_301)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_204),
.Y(n_271)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_131),
.B(n_52),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_153),
.B(n_90),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_207),
.B(n_213),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_123),
.A2(n_104),
.B1(n_103),
.B2(n_96),
.Y(n_208)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g304 ( 
.A(n_211),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_212),
.B(n_245),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_95),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_33),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_217),
.Y(n_284)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_216),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_37),
.Y(n_217)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_173),
.Y(n_219)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_219),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_153),
.B(n_42),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_220),
.B(n_224),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_134),
.A2(n_17),
.B1(n_41),
.B2(n_43),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_222),
.Y(n_255)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_126),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_155),
.A2(n_111),
.B1(n_54),
.B2(n_51),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_231),
.B1(n_120),
.B2(n_112),
.Y(n_260)
);

CKINVDCx12_ASAP7_75t_R g226 ( 
.A(n_177),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_226),
.Y(n_264)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_126),
.B(n_36),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_228),
.B(n_230),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_156),
.B(n_148),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_129),
.B(n_41),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_155),
.A2(n_51),
.B1(n_44),
.B2(n_40),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_129),
.B(n_17),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_232),
.B(n_236),
.Y(n_302)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_128),
.B(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_130),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_125),
.B(n_40),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_239),
.B(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_130),
.Y(n_240)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_145),
.Y(n_241)
);

OA22x2_ASAP7_75t_L g242 ( 
.A1(n_144),
.A2(n_44),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

AND2x2_ASAP7_75t_SL g274 ( 
.A(n_242),
.B(n_6),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_133),
.A2(n_44),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_176),
.Y(n_244)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_170),
.Y(n_245)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_167),
.Y(n_246)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_175),
.Y(n_247)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_247),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_125),
.B(n_2),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_5),
.Y(n_268)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_246),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_172),
.B1(n_160),
.B2(n_170),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_251),
.A2(n_253),
.B1(n_265),
.B2(n_215),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_184),
.A2(n_122),
.B1(n_142),
.B2(n_120),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_184),
.B(n_163),
.C(n_159),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_256),
.B(n_258),
.C(n_272),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_184),
.B(n_121),
.C(n_156),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_260),
.B(n_274),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_196),
.A2(n_112),
.B1(n_167),
.B2(n_115),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g338 ( 
.A1(n_267),
.A2(n_294),
.B(n_299),
.Y(n_338)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_268),
.B(n_11),
.C(n_12),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g272 ( 
.A(n_218),
.B(n_156),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_203),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_279),
.B(n_281),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_280),
.A2(n_297),
.B1(n_235),
.B2(n_187),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_190),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g286 ( 
.A1(n_229),
.A2(n_148),
.B(n_141),
.C(n_151),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_238),
.B(n_195),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_197),
.B(n_161),
.C(n_158),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_291),
.C(n_211),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_288),
.A2(n_195),
.B1(n_188),
.B2(n_238),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_233),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_290),
.B(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_200),
.B(n_161),
.C(n_149),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_222),
.B(n_152),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_293),
.B(n_222),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_140),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_208),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_SL g299 ( 
.A(n_233),
.B(n_10),
.C(n_11),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_209),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx13_ASAP7_75t_L g309 ( 
.A(n_255),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_309),
.Y(n_363)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_310),
.Y(n_376)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_275),
.Y(n_311)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_242),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_313),
.B(n_317),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_314),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_252),
.B(n_204),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_315),
.B(n_316),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_205),
.Y(n_317)
);

OAI22x1_ASAP7_75t_SL g318 ( 
.A1(n_288),
.A2(n_189),
.B1(n_221),
.B2(n_243),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_318),
.A2(n_354),
.B1(n_274),
.B2(n_250),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_259),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_320),
.B(n_323),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_306),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_186),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_332),
.Y(n_372)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_264),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_335),
.Y(n_365)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_328),
.A2(n_265),
.B(n_285),
.Y(n_378)
);

INVx5_ASAP7_75t_L g329 ( 
.A(n_262),
.Y(n_329)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_329),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_330),
.A2(n_339),
.B1(n_344),
.B2(n_356),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_342),
.C(n_287),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_185),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_298),
.B(n_183),
.C(n_193),
.Y(n_333)
);

NOR3xp33_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_349),
.C(n_352),
.Y(n_364)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g336 ( 
.A(n_286),
.B(n_188),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_345),
.Y(n_370)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_340),
.B(n_346),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_256),
.B(n_219),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_343),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_258),
.B(n_216),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_307),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g344 ( 
.A1(n_280),
.A2(n_215),
.B1(n_249),
.B2(n_244),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_257),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_269),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_348),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_284),
.B(n_263),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_307),
.Y(n_381)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_271),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_353),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_266),
.B(n_227),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_271),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_273),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_12),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_294),
.A2(n_199),
.B1(n_247),
.B2(n_14),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_357),
.B(n_373),
.C(n_379),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_316),
.A2(n_274),
.B(n_291),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_361),
.A2(n_362),
.B(n_378),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_328),
.A2(n_250),
.B(n_255),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_366),
.A2(n_380),
.B1(n_384),
.B2(n_386),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_278),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_319),
.B(n_260),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_312),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_270),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_318),
.A2(n_297),
.B1(n_292),
.B2(n_262),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_292),
.B1(n_295),
.B2(n_282),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_296),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_389),
.C(n_394),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_347),
.A2(n_301),
.B1(n_254),
.B2(n_304),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_347),
.A2(n_304),
.B1(n_301),
.B2(n_285),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_341),
.B(n_273),
.C(n_289),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_321),
.B(n_289),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_393),
.B(n_308),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_313),
.B(n_254),
.C(n_202),
.Y(n_394)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_396),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_317),
.B(n_13),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_311),
.Y(n_409)
);

AND2x6_ASAP7_75t_L g398 ( 
.A(n_370),
.B(n_336),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_405),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_322),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_399),
.B(n_403),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_338),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_402),
.A2(n_431),
.B(n_394),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_372),
.B(n_324),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_380),
.A2(n_332),
.B1(n_354),
.B2(n_312),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_404),
.A2(n_329),
.B1(n_348),
.B2(n_309),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_358),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_408),
.B(n_418),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_409),
.B(n_429),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_410),
.B(n_416),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_310),
.Y(n_411)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_411),
.Y(n_441)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_412),
.Y(n_448)
);

INVx13_ASAP7_75t_L g413 ( 
.A(n_363),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_390),
.Y(n_414)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_414),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_358),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_421),
.Y(n_444)
);

BUFx12_ASAP7_75t_L g416 ( 
.A(n_363),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_362),
.A2(n_343),
.B(n_340),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_417),
.A2(n_371),
.B(n_358),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_368),
.B(n_350),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_419),
.B(n_427),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_355),
.Y(n_420)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_353),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_423),
.B(n_425),
.Y(n_447)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_351),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_428),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_325),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

NOR2x1_ASAP7_75t_L g429 ( 
.A(n_359),
.B(n_366),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_378),
.A2(n_337),
.B(n_327),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_389),
.B(n_346),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_432),
.B(n_379),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_433),
.A2(n_446),
.B(n_459),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_434),
.B(n_403),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_418),
.B(n_373),
.C(n_385),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_456),
.C(n_430),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g437 ( 
.A(n_402),
.B(n_359),
.CI(n_357),
.CON(n_437),
.SN(n_437)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_437),
.B(n_400),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_406),
.A2(n_386),
.B1(n_384),
.B2(n_361),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_438),
.A2(n_445),
.B1(n_458),
.B2(n_404),
.Y(n_470)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_412),
.A2(n_368),
.B1(n_395),
.B2(n_391),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_399),
.B(n_365),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_449),
.B(n_450),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_419),
.B(n_360),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_371),
.B(n_376),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_417),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_408),
.B(n_396),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_432),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_374),
.C(n_392),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_427),
.B(n_401),
.Y(n_457)
);

NOR2x1_ASAP7_75t_L g467 ( 
.A(n_457),
.B(n_410),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_405),
.A2(n_392),
.B1(n_374),
.B2(n_377),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_424),
.A2(n_377),
.B(n_364),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_461),
.A2(n_422),
.B1(n_423),
.B2(n_413),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_469),
.C(n_476),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_465),
.B(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_467),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_435),
.A2(n_424),
.B1(n_431),
.B2(n_429),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_468),
.B(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_415),
.C(n_421),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_470),
.A2(n_435),
.B1(n_440),
.B2(n_448),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_456),
.B(n_429),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_471),
.B(n_486),
.Y(n_498)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_444),
.Y(n_473)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_473),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_475),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_434),
.B(n_420),
.C(n_411),
.Y(n_476)
);

NOR2x1_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_401),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_444),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_478),
.B(n_482),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_409),
.C(n_426),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_479),
.B(n_483),
.C(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_460),
.B(n_407),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_480),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_481),
.A2(n_459),
.B(n_439),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_453),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_454),
.B(n_428),
.C(n_425),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_414),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_488),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_439),
.B(n_398),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_487),
.B(n_433),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_457),
.B(n_202),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g526 ( 
.A(n_489),
.B(n_495),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_491),
.B(n_496),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_492),
.A2(n_451),
.B1(n_468),
.B2(n_473),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_438),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_446),
.C(n_458),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_499),
.C(n_447),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_448),
.C(n_440),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_442),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_506),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_472),
.B(n_445),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_505),
.B(n_479),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_465),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_466),
.B(n_451),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_507),
.B(n_475),
.Y(n_515)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_510),
.Y(n_527)
);

AOI221xp5_ASAP7_75t_L g512 ( 
.A1(n_504),
.A2(n_480),
.B1(n_455),
.B2(n_485),
.C(n_463),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_512),
.B(n_520),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_494),
.A2(n_470),
.B1(n_474),
.B2(n_485),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_513),
.B(n_521),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_522),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_515),
.B(n_506),
.Y(n_536)
);

BUFx12_ASAP7_75t_L g517 ( 
.A(n_499),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_517),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_451),
.B1(n_487),
.B2(n_441),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_518),
.A2(n_523),
.B1(n_447),
.B2(n_462),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_509),
.A2(n_477),
.B(n_441),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_507),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_508),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_497),
.B(n_461),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_500),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_490),
.A2(n_455),
.B1(n_462),
.B2(n_460),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_498),
.C(n_493),
.Y(n_531)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_501),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_525),
.A2(n_437),
.B1(n_503),
.B2(n_453),
.Y(n_540)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_528),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_518),
.A2(n_510),
.B(n_489),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_529),
.A2(n_516),
.B1(n_526),
.B2(n_515),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_531),
.B(n_534),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_521),
.A2(n_496),
.B1(n_498),
.B2(n_495),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_536),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_519),
.A2(n_437),
.B1(n_398),
.B2(n_493),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_524),
.B(n_502),
.C(n_503),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_537),
.B(n_511),
.C(n_526),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_511),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_540),
.B(n_416),
.Y(n_550)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_541),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_467),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_542),
.B(n_543),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_544),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_531),
.B(n_517),
.C(n_416),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_546),
.B(n_536),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_517),
.B1(n_413),
.B2(n_416),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_529),
.C(n_528),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_550),
.A2(n_535),
.B(n_534),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_552),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_545),
.A2(n_538),
.B1(n_535),
.B2(n_527),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_553),
.B(n_546),
.C(n_543),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_554),
.A2(n_547),
.B1(n_544),
.B2(n_533),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_558),
.B(n_559),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_555),
.B(n_556),
.C(n_557),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_561),
.B(n_551),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_563),
.B(n_560),
.Y(n_564)
);

O2A1O1Ixp33_ASAP7_75t_SL g565 ( 
.A1(n_564),
.A2(n_562),
.B(n_548),
.C(n_537),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_548),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_566),
.A2(n_202),
.B(n_13),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_13),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_13),
.Y(n_569)
);


endmodule