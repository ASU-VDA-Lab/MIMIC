module fake_jpeg_31704_n_206 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_206);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_22),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_35),
.Y(n_58)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_31),
.Y(n_62)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_7),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_18),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_8),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_25),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_65),
.B1(n_68),
.B2(n_77),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_13),
.B1(n_26),
.B2(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_38),
.A2(n_28),
.B1(n_13),
.B2(n_21),
.Y(n_66)
);

OAI22x1_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_87),
.B1(n_69),
.B2(n_59),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_71),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_51),
.A2(n_20),
.B1(n_19),
.B2(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_33),
.B(n_20),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_57),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_76),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_14),
.B1(n_6),
.B2(n_5),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_14),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_6),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_48),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_104),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_36),
.B1(n_44),
.B2(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_91),
.B1(n_97),
.B2(n_61),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_93),
.A2(n_109),
.B1(n_98),
.B2(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_9),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_105),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_54),
.B(n_10),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_116),
.C(n_63),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_113),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_11),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_107),
.B(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_83),
.Y(n_110)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g127 ( 
.A(n_111),
.Y(n_127)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_60),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_86),
.Y(n_116)
);

AO22x1_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_82),
.B1(n_63),
.B2(n_56),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_116),
.B(n_96),
.Y(n_143)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_121),
.B1(n_90),
.B2(n_89),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_109),
.A2(n_61),
.B1(n_73),
.B2(n_82),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_122),
.B(n_125),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_79),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_99),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_99),
.B(n_55),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_55),
.A3(n_74),
.B1(n_107),
.B2(n_92),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_114),
.B(n_95),
.C(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_114),
.B1(n_98),
.B2(n_103),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_126),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_141),
.C(n_145),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_89),
.B(n_92),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_150),
.B1(n_117),
.B2(n_119),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_100),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_144),
.B(n_149),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_117),
.B(n_121),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_SL g163 ( 
.A(n_147),
.B(n_124),
.C(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_105),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_142),
.B(n_128),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_132),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_141),
.B1(n_101),
.B2(n_129),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_147),
.C(n_138),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_139),
.A2(n_136),
.B(n_129),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_166),
.B(n_101),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_136),
.C(n_104),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_140),
.B1(n_144),
.B2(n_143),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_173),
.B(n_178),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_163),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_133),
.C(n_111),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_177),
.C(n_165),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_133),
.C(n_112),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_179),
.B(n_180),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_171),
.B(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_183),
.B(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_159),
.C(n_154),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_160),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_161),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_172),
.B1(n_173),
.B2(n_169),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_137),
.C(n_115),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_169),
.B1(n_174),
.B2(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_180),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_167),
.B(n_153),
.Y(n_192)
);

OAI31xp33_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_184),
.A3(n_183),
.B(n_181),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_195),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_196),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_192),
.A2(n_179),
.B(n_127),
.C(n_137),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_187),
.B(n_189),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_120),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_198),
.B1(n_191),
.B2(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_191),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_202),
.B(n_120),
.Y(n_204)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_200),
.B(n_74),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_203),
.Y(n_206)
);


endmodule