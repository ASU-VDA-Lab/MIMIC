module fake_netlist_1_9108_n_1607 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1607);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1607;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1603;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1605;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_1595;
wire n_1604;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1600;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1602;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_1606;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_1537;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1601;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1335;
wire n_1239;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_167), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_267), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_178), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_79), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_294), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_210), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_347), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_50), .Y(n_360) );
BUFx6f_ASAP7_75t_L g361 ( .A(n_106), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_339), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_185), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_319), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_22), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g367 ( .A(n_211), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_133), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_104), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_221), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_298), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_158), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_27), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_82), .Y(n_374) );
INVxp33_ASAP7_75t_L g375 ( .A(n_255), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_193), .Y(n_376) );
INVx4_ASAP7_75t_R g377 ( .A(n_209), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_171), .Y(n_378) );
INVxp33_ASAP7_75t_L g379 ( .A(n_254), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_157), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_187), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_15), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_204), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_333), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_58), .B(n_199), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_256), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_217), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_344), .Y(n_388) );
CKINVDCx14_ASAP7_75t_R g389 ( .A(n_349), .Y(n_389) );
BUFx3_ASAP7_75t_L g390 ( .A(n_313), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_348), .Y(n_391) );
BUFx2_ASAP7_75t_L g392 ( .A(n_145), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_42), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
CKINVDCx16_ASAP7_75t_R g395 ( .A(n_250), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_295), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_149), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_342), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_277), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_230), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_12), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_123), .B(n_257), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_141), .Y(n_403) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_335), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_113), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_35), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_351), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_188), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_147), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_81), .B(n_144), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_142), .Y(n_411) );
INVx1_ASAP7_75t_SL g412 ( .A(n_21), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_181), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_29), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_300), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_284), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_28), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_43), .Y(n_418) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_233), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_266), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_8), .Y(n_421) );
BUFx10_ASAP7_75t_L g422 ( .A(n_82), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_15), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_53), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_263), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_151), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_60), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g428 ( .A(n_352), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_283), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_6), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_328), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_195), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_306), .Y(n_433) );
INVxp33_ASAP7_75t_L g434 ( .A(n_215), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_67), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_43), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_320), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_106), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_241), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_274), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_259), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_156), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_76), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_186), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_99), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_134), .Y(n_446) );
BUFx2_ASAP7_75t_SL g447 ( .A(n_173), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_275), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_293), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_120), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_97), .Y(n_451) );
INVxp33_ASAP7_75t_L g452 ( .A(n_94), .Y(n_452) );
CKINVDCx16_ASAP7_75t_R g453 ( .A(n_100), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_251), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_34), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_112), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_59), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_127), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_96), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_258), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_304), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_189), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_14), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_19), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_53), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_175), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_169), .Y(n_467) );
INVxp33_ASAP7_75t_SL g468 ( .A(n_176), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_60), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_252), .Y(n_470) );
INVxp33_ASAP7_75t_SL g471 ( .A(n_119), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_308), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_196), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_71), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_78), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_151), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_14), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_225), .Y(n_478) );
BUFx5_ASAP7_75t_L g479 ( .A(n_203), .Y(n_479) );
INVxp67_ASAP7_75t_L g480 ( .A(n_58), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_25), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_326), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_247), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_17), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_37), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_281), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_16), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_331), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_150), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_86), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_123), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_73), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_206), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_231), .Y(n_494) );
INVxp67_ASAP7_75t_L g495 ( .A(n_37), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_168), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_35), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_63), .Y(n_498) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_61), .B(n_68), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_321), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_329), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_46), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_71), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_177), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_144), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_48), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_63), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_288), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_101), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_297), .Y(n_510) );
BUFx3_ASAP7_75t_L g511 ( .A(n_261), .Y(n_511) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_180), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_120), .Y(n_513) );
BUFx3_ASAP7_75t_L g514 ( .A(n_279), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_246), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_138), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_74), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_346), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_202), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_184), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_6), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_240), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_86), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_23), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_228), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_208), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_216), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_45), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_3), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_124), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_198), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_243), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_245), .Y(n_533) );
INVx1_ASAP7_75t_SL g534 ( .A(n_55), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_269), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_174), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_341), .Y(n_537) );
INVxp67_ASAP7_75t_L g538 ( .A(n_146), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_280), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_183), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_9), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_338), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_46), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_375), .B(n_0), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_373), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_432), .B(n_0), .Y(n_547) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_404), .Y(n_548) );
INVx3_ASAP7_75t_L g549 ( .A(n_456), .Y(n_549) );
BUFx3_ASAP7_75t_L g550 ( .A(n_358), .Y(n_550) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_404), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_373), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_452), .B(n_375), .Y(n_553) );
OA21x2_ASAP7_75t_L g554 ( .A1(n_357), .A2(n_1), .B(n_2), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_456), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_382), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_382), .Y(n_557) );
INVx5_ASAP7_75t_L g558 ( .A(n_404), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_397), .Y(n_559) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_435), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_435), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_479), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_397), .Y(n_563) );
INVx6_ASAP7_75t_L g564 ( .A(n_479), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_479), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_479), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_403), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_479), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_403), .Y(n_569) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_357), .A2(n_155), .B(n_154), .Y(n_570) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_404), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_426), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_426), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_452), .B(n_4), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_443), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_443), .Y(n_576) );
INVx2_ASAP7_75t_SL g577 ( .A(n_415), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_446), .B(n_4), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_446), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_379), .B(n_5), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_479), .Y(n_581) );
OAI22xp5_ASAP7_75t_SL g582 ( .A1(n_427), .A2(n_8), .B1(n_5), .B2(n_7), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_450), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_450), .Y(n_584) );
INVx3_ASAP7_75t_L g585 ( .A(n_365), .Y(n_585) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_358), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_513), .B(n_7), .Y(n_587) );
INVx4_ASAP7_75t_L g588 ( .A(n_564), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_553), .B(n_561), .Y(n_589) );
BUFx2_ASAP7_75t_L g590 ( .A(n_561), .Y(n_590) );
INVx4_ASAP7_75t_L g591 ( .A(n_564), .Y(n_591) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_553), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_553), .B(n_379), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_548), .Y(n_594) );
NOR2xp33_ASAP7_75t_SL g595 ( .A(n_580), .B(n_367), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_549), .B(n_434), .Y(n_596) );
AND3x2_ASAP7_75t_L g597 ( .A(n_580), .B(n_411), .C(n_392), .Y(n_597) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_580), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_564), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_548), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_548), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_577), .B(n_434), .Y(n_602) );
AND2x6_ASAP7_75t_L g603 ( .A(n_578), .B(n_364), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_578), .A2(n_587), .B1(n_554), .B2(n_585), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_578), .B(n_365), .Y(n_605) );
BUFx4_ASAP7_75t_L g606 ( .A(n_574), .Y(n_606) );
BUFx8_ASAP7_75t_SL g607 ( .A(n_547), .Y(n_607) );
BUFx8_ASAP7_75t_SL g608 ( .A(n_547), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_545), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_578), .A2(n_368), .B1(n_369), .B2(n_356), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_549), .B(n_396), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_545), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_549), .B(n_396), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_545), .Y(n_614) );
INVx3_ASAP7_75t_L g615 ( .A(n_564), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_549), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_549), .B(n_408), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_545), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_562), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_562), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_555), .B(n_408), .Y(n_621) );
INVx5_ASAP7_75t_L g622 ( .A(n_564), .Y(n_622) );
INVx2_ASAP7_75t_SL g623 ( .A(n_564), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_578), .B(n_444), .Y(n_624) );
INVx3_ASAP7_75t_L g625 ( .A(n_587), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_562), .Y(n_626) );
INVxp33_ASAP7_75t_L g627 ( .A(n_574), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_577), .B(n_386), .Y(n_628) );
NOR2x1p5_ASAP7_75t_L g629 ( .A(n_547), .B(n_393), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_627), .B(n_577), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_625), .A2(n_587), .B(n_547), .C(n_565), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_593), .B(n_587), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_596), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_625), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_595), .B(n_395), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_592), .A2(n_544), .B1(n_587), .B2(n_471), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_595), .A2(n_453), .B1(n_560), .B2(n_498), .Y(n_638) );
BUFx2_ASAP7_75t_L g639 ( .A(n_607), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_610), .B(n_441), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_616), .Y(n_641) );
NAND2x1_ASAP7_75t_L g642 ( .A(n_603), .B(n_377), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_590), .B(n_544), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_550), .Y(n_644) );
AO22x1_ASAP7_75t_L g645 ( .A1(n_598), .A2(n_560), .B1(n_471), .B2(n_468), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_625), .Y(n_646) );
NAND2xp33_ASAP7_75t_SL g647 ( .A(n_629), .B(n_353), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_610), .B(n_532), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_629), .B(n_517), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_590), .B(n_422), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_602), .B(n_550), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_625), .Y(n_652) );
O2A1O1Ixp5_ASAP7_75t_L g653 ( .A1(n_605), .A2(n_555), .B(n_512), .C(n_388), .Y(n_653) );
BUFx3_ASAP7_75t_L g654 ( .A(n_590), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_602), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_589), .B(n_363), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_611), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_611), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_603), .B(n_555), .Y(n_659) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_589), .B(n_363), .Y(n_660) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_589), .A2(n_370), .B1(n_371), .B2(n_353), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_628), .B(n_468), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_603), .A2(n_554), .B1(n_566), .B2(n_565), .Y(n_663) );
INVx5_ASAP7_75t_L g664 ( .A(n_603), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g665 ( .A(n_588), .B(n_372), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_607), .B(n_391), .Y(n_666) );
NOR2x2_ASAP7_75t_L g667 ( .A(n_606), .B(n_427), .Y(n_667) );
NOR2x1p5_ASAP7_75t_L g668 ( .A(n_597), .B(n_393), .Y(n_668) );
AOI22xp5_ASAP7_75t_SL g669 ( .A1(n_606), .A2(n_523), .B1(n_498), .B2(n_371), .Y(n_669) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_608), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_603), .A2(n_429), .B1(n_454), .B2(n_370), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g672 ( .A1(n_606), .A2(n_582), .B1(n_523), .B2(n_429), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_624), .B(n_448), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_624), .B(n_448), .Y(n_674) );
INVx4_ASAP7_75t_L g675 ( .A(n_588), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_604), .B(n_478), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_597), .B(n_454), .Y(n_677) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_609), .A2(n_519), .B1(n_531), .B2(n_467), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_609), .B(n_510), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_608), .B(n_483), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_613), .B(n_467), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_612), .A2(n_554), .B1(n_566), .B2(n_565), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_613), .B(n_519), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_617), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_614), .B(n_539), .Y(n_685) );
INVxp67_ASAP7_75t_L g686 ( .A(n_617), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_621), .B(n_531), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_588), .B(n_362), .Y(n_688) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_588), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_621), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_619), .Y(n_691) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_619), .A2(n_581), .B(n_568), .C(n_570), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_620), .B(n_568), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_591), .B(n_546), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_620), .A2(n_582), .B1(n_455), .B2(n_464), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_626), .B(n_568), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_623), .A2(n_570), .B(n_568), .Y(n_697) );
OR2x6_ASAP7_75t_L g698 ( .A(n_591), .B(n_499), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_626), .B(n_581), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_618), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_623), .A2(n_457), .B1(n_464), .B2(n_455), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_591), .B(n_581), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_654), .Y(n_703) );
OR2x6_ASAP7_75t_SL g704 ( .A(n_670), .B(n_457), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_646), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_675), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_686), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_661), .B(n_507), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_697), .A2(n_591), .B(n_623), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_657), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_630), .B(n_591), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_SL g712 ( .A1(n_692), .A2(n_355), .B(n_359), .C(n_354), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_702), .A2(n_615), .B(n_599), .Y(n_713) );
NOR2xp33_ASAP7_75t_R g714 ( .A(n_647), .B(n_389), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g715 ( .A1(n_655), .A2(n_430), .B(n_495), .C(n_480), .Y(n_715) );
AND2x4_ASAP7_75t_L g716 ( .A(n_634), .B(n_374), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_658), .B(n_507), .Y(n_717) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_664), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_633), .A2(n_615), .B(n_599), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_649), .B(n_360), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_684), .B(n_538), .Y(n_721) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_664), .Y(n_722) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_633), .A2(n_622), .B(n_554), .Y(n_723) );
NOR2xp33_ASAP7_75t_SL g724 ( .A(n_664), .B(n_622), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_649), .B(n_366), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_635), .Y(n_726) );
BUFx2_ASAP7_75t_L g727 ( .A(n_667), .Y(n_727) );
OR2x6_ASAP7_75t_SL g728 ( .A(n_669), .B(n_405), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_681), .B(n_422), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_652), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_694), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_690), .B(n_554), .Y(n_732) );
INVx2_ASAP7_75t_L g733 ( .A(n_694), .Y(n_733) );
O2A1O1Ixp33_ASAP7_75t_L g734 ( .A1(n_638), .A2(n_410), .B(n_414), .C(n_401), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_644), .Y(n_735) );
BUFx12f_ASAP7_75t_L g736 ( .A(n_639), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_651), .Y(n_737) );
INVxp67_ASAP7_75t_L g738 ( .A(n_631), .Y(n_738) );
INVx2_ASAP7_75t_SL g739 ( .A(n_681), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_631), .B(n_585), .Y(n_740) );
INVx1_ASAP7_75t_L g741 ( .A(n_693), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_671), .A2(n_585), .B1(n_417), .B2(n_421), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_691), .B(n_406), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_683), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_683), .B(n_422), .Y(n_745) );
AND2x4_ASAP7_75t_L g746 ( .A(n_650), .B(n_418), .Y(n_746) );
INVx8_ASAP7_75t_L g747 ( .A(n_698), .Y(n_747) );
O2A1O1Ixp33_ASAP7_75t_L g748 ( .A1(n_640), .A2(n_423), .B(n_445), .C(n_438), .Y(n_748) );
CKINVDCx8_ASAP7_75t_R g749 ( .A(n_677), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_637), .B(n_409), .Y(n_750) );
INVxp67_ASAP7_75t_L g751 ( .A(n_687), .Y(n_751) );
OR2x6_ASAP7_75t_L g752 ( .A(n_677), .B(n_447), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_662), .A2(n_451), .B(n_459), .C(n_458), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_656), .B(n_463), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_693), .Y(n_755) );
O2A1O1Ixp33_ASAP7_75t_L g756 ( .A1(n_648), .A2(n_469), .B(n_475), .C(n_465), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_660), .B(n_528), .Y(n_757) );
INVx5_ASAP7_75t_L g758 ( .A(n_689), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g759 ( .A1(n_663), .A2(n_476), .B1(n_481), .B2(n_477), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_643), .B(n_530), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_653), .A2(n_484), .B(n_487), .C(n_485), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_641), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_643), .B(n_412), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_687), .B(n_436), .Y(n_764) );
OR2x6_ASAP7_75t_L g765 ( .A(n_645), .B(n_513), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_698), .B(n_489), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_636), .A2(n_534), .B1(n_474), .B2(n_402), .Y(n_767) );
INVx4_ASAP7_75t_L g768 ( .A(n_689), .Y(n_768) );
BUFx8_ASAP7_75t_SL g769 ( .A(n_698), .Y(n_769) );
O2A1O1Ixp5_ASAP7_75t_L g770 ( .A1(n_642), .A2(n_385), .B(n_462), .C(n_444), .Y(n_770) );
AND2x6_ASAP7_75t_L g771 ( .A(n_659), .B(n_364), .Y(n_771) );
BUFx2_ASAP7_75t_L g772 ( .A(n_678), .Y(n_772) );
AND2x6_ASAP7_75t_SL g773 ( .A(n_666), .B(n_385), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_696), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_699), .B(n_490), .Y(n_775) );
A2O1A1Ixp33_ASAP7_75t_L g776 ( .A1(n_699), .A2(n_492), .B(n_497), .C(n_491), .Y(n_776) );
INVxp67_ASAP7_75t_L g777 ( .A(n_701), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_676), .A2(n_503), .B1(n_505), .B2(n_502), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_679), .Y(n_779) );
OA21x2_ASAP7_75t_L g780 ( .A1(n_682), .A2(n_600), .B(n_594), .Y(n_780) );
NOR2xp33_ASAP7_75t_R g781 ( .A(n_680), .B(n_384), .Y(n_781) );
NAND2xp33_ASAP7_75t_SL g782 ( .A(n_668), .B(n_387), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_673), .B(n_506), .Y(n_783) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_685), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_674), .B(n_665), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_695), .A2(n_516), .B1(n_521), .B2(n_509), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_700), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_688), .B(n_524), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_672), .B(n_546), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_646), .Y(n_790) );
NOR3xp33_ASAP7_75t_SL g791 ( .A(n_638), .B(n_419), .C(n_416), .Y(n_791) );
INVx2_ASAP7_75t_SL g792 ( .A(n_654), .Y(n_792) );
NAND2xp5_ASAP7_75t_SL g793 ( .A(n_686), .B(n_428), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_686), .Y(n_794) );
INVxp67_ASAP7_75t_L g795 ( .A(n_654), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_686), .B(n_529), .Y(n_796) );
INVx3_ASAP7_75t_L g797 ( .A(n_675), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_675), .Y(n_798) );
BUFx3_ASAP7_75t_L g799 ( .A(n_639), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_632), .A2(n_543), .B(n_541), .C(n_552), .Y(n_800) );
AND2x2_ASAP7_75t_SL g801 ( .A(n_671), .B(n_361), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_630), .B(n_552), .Y(n_802) );
AND2x4_ASAP7_75t_L g803 ( .A(n_655), .B(n_556), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_630), .B(n_557), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_654), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_654), .B(n_376), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_686), .Y(n_807) );
INVx2_ASAP7_75t_L g808 ( .A(n_646), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_686), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_654), .B(n_381), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_657), .A2(n_559), .B1(n_563), .B2(n_557), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_646), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g813 ( .A1(n_697), .A2(n_601), .B(n_383), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_654), .B(n_559), .Y(n_814) );
AND2x4_ASAP7_75t_L g815 ( .A(n_655), .B(n_563), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_654), .Y(n_816) );
AND2x2_ASAP7_75t_SL g817 ( .A(n_671), .B(n_361), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_686), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_646), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_646), .Y(n_820) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_657), .A2(n_569), .B1(n_572), .B2(n_567), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_710), .Y(n_822) );
AND2x6_ASAP7_75t_L g823 ( .A(n_741), .B(n_466), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_707), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_755), .Y(n_825) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_786), .A2(n_567), .B1(n_573), .B2(n_572), .C(n_569), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_738), .B(n_573), .Y(n_827) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_732), .A2(n_394), .B(n_380), .Y(n_828) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_758), .Y(n_829) );
BUFx3_ASAP7_75t_L g830 ( .A(n_736), .Y(n_830) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_805), .Y(n_831) );
A2O1A1Ixp33_ASAP7_75t_L g832 ( .A1(n_779), .A2(n_399), .B(n_400), .C(n_398), .Y(n_832) );
AOI21xp5_ASAP7_75t_L g833 ( .A1(n_813), .A2(n_425), .B(n_420), .Y(n_833) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_786), .A2(n_579), .B1(n_583), .B2(n_576), .C(n_575), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_794), .Y(n_835) );
AOI221x1_ASAP7_75t_L g836 ( .A1(n_759), .A2(n_586), .B1(n_433), .B2(n_442), .C(n_440), .Y(n_836) );
AO31x2_ASAP7_75t_L g837 ( .A1(n_759), .A2(n_493), .A3(n_576), .B(n_575), .Y(n_837) );
CKINVDCx11_ASAP7_75t_R g838 ( .A(n_704), .Y(n_838) );
O2A1O1Ixp33_ASAP7_75t_L g839 ( .A1(n_753), .A2(n_583), .B(n_584), .C(n_579), .Y(n_839) );
INVx1_ASAP7_75t_SL g840 ( .A(n_703), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_807), .Y(n_841) );
O2A1O1Ixp33_ASAP7_75t_L g842 ( .A1(n_800), .A2(n_584), .B(n_449), .C(n_460), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g843 ( .A1(n_728), .A2(n_424), .B1(n_361), .B2(n_431), .Y(n_843) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_758), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_809), .B(n_361), .Y(n_845) );
BUFx2_ASAP7_75t_L g846 ( .A(n_816), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_769), .Y(n_847) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_765), .A2(n_424), .B1(n_439), .B2(n_437), .Y(n_848) );
INVx1_ASAP7_75t_SL g849 ( .A(n_792), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_818), .B(n_424), .Y(n_850) );
A2O1A1Ixp33_ASAP7_75t_L g851 ( .A1(n_774), .A2(n_472), .B(n_473), .C(n_470), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_777), .B(n_407), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_716), .B(n_482), .Y(n_853) );
A2O1A1Ixp33_ASAP7_75t_L g854 ( .A1(n_785), .A2(n_488), .B(n_494), .C(n_486), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_716), .B(n_496), .Y(n_855) );
OAI21xp5_ASAP7_75t_L g856 ( .A1(n_723), .A2(n_501), .B(n_500), .Y(n_856) );
AO31x2_ASAP7_75t_L g857 ( .A1(n_811), .A2(n_508), .A3(n_515), .B(n_504), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_787), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_799), .Y(n_859) );
AO31x2_ASAP7_75t_L g860 ( .A1(n_811), .A2(n_520), .A3(n_522), .B(n_518), .Y(n_860) );
NOR2xp33_ASAP7_75t_L g861 ( .A(n_772), .B(n_461), .Y(n_861) );
AND2x4_ASAP7_75t_L g862 ( .A(n_739), .B(n_525), .Y(n_862) );
OAI21xp5_ASAP7_75t_L g863 ( .A1(n_719), .A2(n_527), .B(n_526), .Y(n_863) );
BUFx2_ASAP7_75t_L g864 ( .A(n_795), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_705), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_751), .B(n_533), .Y(n_866) );
AO32x2_ASAP7_75t_L g867 ( .A1(n_821), .A2(n_586), .A3(n_571), .B1(n_551), .B2(n_548), .Y(n_867) );
O2A1O1Ixp33_ASAP7_75t_SL g868 ( .A1(n_761), .A2(n_536), .B(n_537), .C(n_535), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_709), .A2(n_542), .B(n_540), .Y(n_869) );
A2O1A1Ixp33_ASAP7_75t_L g870 ( .A1(n_783), .A2(n_390), .B(n_413), .C(n_378), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_744), .B(n_9), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_764), .B(n_10), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_814), .Y(n_873) );
OAI222xp33_ASAP7_75t_L g874 ( .A1(n_765), .A2(n_413), .B1(n_511), .B2(n_514), .C1(n_13), .C2(n_16), .Y(n_874) );
AO31x2_ASAP7_75t_L g875 ( .A1(n_821), .A2(n_586), .A3(n_551), .B(n_571), .Y(n_875) );
A2O1A1Ixp33_ASAP7_75t_L g876 ( .A1(n_748), .A2(n_756), .B(n_770), .C(n_788), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_790), .Y(n_877) );
AO31x2_ASAP7_75t_L g878 ( .A1(n_778), .A2(n_586), .A3(n_551), .B(n_571), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_780), .A2(n_586), .B(n_551), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_729), .Y(n_880) );
INVx1_ASAP7_75t_L g881 ( .A(n_802), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_801), .A2(n_586), .B1(n_551), .B2(n_571), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_784), .B(n_10), .Y(n_883) );
INVx1_ASAP7_75t_SL g884 ( .A(n_758), .Y(n_884) );
NAND2x1p5_ASAP7_75t_L g885 ( .A(n_768), .B(n_558), .Y(n_885) );
AO31x2_ASAP7_75t_L g886 ( .A1(n_778), .A2(n_551), .A3(n_571), .B(n_548), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_808), .Y(n_887) );
OAI22xp33_ASAP7_75t_L g888 ( .A1(n_765), .A2(n_558), .B1(n_13), .B2(n_11), .Y(n_888) );
NOR2xp67_ASAP7_75t_L g889 ( .A(n_767), .B(n_11), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_746), .B(n_12), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_708), .B(n_17), .Y(n_891) );
NOR2xp33_ASAP7_75t_SL g892 ( .A(n_749), .B(n_558), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_812), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_819), .Y(n_894) );
AOI221xp5_ASAP7_75t_SL g895 ( .A1(n_734), .A2(n_571), .B1(n_20), .B2(n_18), .C(n_19), .Y(n_895) );
OAI21x1_ASAP7_75t_L g896 ( .A1(n_780), .A2(n_160), .B(n_159), .Y(n_896) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_727), .A2(n_558), .B1(n_22), .B2(n_18), .Y(n_897) );
AO31x2_ASAP7_75t_L g898 ( .A1(n_776), .A2(n_24), .A3(n_20), .B(n_23), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_820), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_746), .B(n_24), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_817), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_745), .B(n_26), .Y(n_902) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_715), .A2(n_30), .B1(n_28), .B2(n_29), .C(n_31), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_789), .B(n_30), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_726), .Y(n_905) );
AO32x2_ASAP7_75t_L g906 ( .A1(n_742), .A2(n_33), .A3(n_31), .B1(n_32), .B2(n_34), .Y(n_906) );
OAI21xp5_ASAP7_75t_L g907 ( .A1(n_711), .A2(n_162), .B(n_161), .Y(n_907) );
A2O1A1Ixp33_ASAP7_75t_L g908 ( .A1(n_735), .A2(n_36), .B(n_32), .C(n_33), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_721), .B(n_36), .Y(n_909) );
A2O1A1Ixp33_ASAP7_75t_L g910 ( .A1(n_737), .A2(n_40), .B(n_38), .C(n_39), .Y(n_910) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_742), .A2(n_40), .B1(n_38), .B2(n_39), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_730), .Y(n_912) );
OAI21xp5_ASAP7_75t_L g913 ( .A1(n_711), .A2(n_164), .B(n_163), .Y(n_913) );
OAI21x1_ASAP7_75t_L g914 ( .A1(n_713), .A2(n_166), .B(n_165), .Y(n_914) );
BUFx10_ASAP7_75t_L g915 ( .A(n_752), .Y(n_915) );
OR2x6_ASAP7_75t_L g916 ( .A(n_747), .B(n_41), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g917 ( .A1(n_720), .A2(n_44), .B1(n_41), .B2(n_42), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_717), .B(n_44), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_804), .A2(n_48), .B1(n_45), .B2(n_47), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_796), .B(n_47), .Y(n_920) );
OR2x2_ASAP7_75t_L g921 ( .A(n_750), .B(n_49), .Y(n_921) );
NOR2xp33_ASAP7_75t_SL g922 ( .A(n_752), .B(n_51), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_740), .Y(n_923) );
AND2x4_ASAP7_75t_L g924 ( .A(n_752), .B(n_52), .Y(n_924) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_743), .A2(n_55), .B1(n_52), .B2(n_54), .Y(n_925) );
NAND2x1p5_ASAP7_75t_L g926 ( .A(n_768), .B(n_54), .Y(n_926) );
BUFx3_ASAP7_75t_L g927 ( .A(n_747), .Y(n_927) );
OAI21xp5_ASAP7_75t_L g928 ( .A1(n_712), .A2(n_172), .B(n_170), .Y(n_928) );
AOI221x1_ASAP7_75t_L g929 ( .A1(n_766), .A2(n_56), .B1(n_57), .B2(n_59), .C(n_61), .Y(n_929) );
AO31x2_ASAP7_75t_L g930 ( .A1(n_775), .A2(n_62), .A3(n_56), .B(n_57), .Y(n_930) );
OR2x2_ASAP7_75t_L g931 ( .A(n_750), .B(n_62), .Y(n_931) );
AO31x2_ASAP7_75t_L g932 ( .A1(n_775), .A2(n_66), .A3(n_64), .B(n_65), .Y(n_932) );
A2O1A1Ixp33_ASAP7_75t_L g933 ( .A1(n_763), .A2(n_66), .B(n_64), .C(n_65), .Y(n_933) );
INVx1_ASAP7_75t_L g934 ( .A(n_740), .Y(n_934) );
AOI21xp5_ASAP7_75t_L g935 ( .A1(n_743), .A2(n_182), .B(n_179), .Y(n_935) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_747), .A2(n_69), .B1(n_67), .B2(n_68), .Y(n_936) );
A2O1A1Ixp33_ASAP7_75t_L g937 ( .A1(n_760), .A2(n_72), .B(n_69), .C(n_70), .Y(n_937) );
INVx2_ASAP7_75t_L g938 ( .A(n_762), .Y(n_938) );
OR2x2_ASAP7_75t_L g939 ( .A(n_725), .B(n_70), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_754), .B(n_75), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_803), .Y(n_941) );
INVx3_ASAP7_75t_SL g942 ( .A(n_754), .Y(n_942) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_791), .A2(n_76), .B(n_77), .C(n_78), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_803), .B(n_77), .Y(n_944) );
NOR2xp33_ASAP7_75t_R g945 ( .A(n_782), .B(n_773), .Y(n_945) );
AOI21xp33_ASAP7_75t_L g946 ( .A1(n_806), .A2(n_79), .B(n_80), .Y(n_946) );
INVx3_ASAP7_75t_L g947 ( .A(n_706), .Y(n_947) );
A2O1A1Ixp33_ASAP7_75t_L g948 ( .A1(n_815), .A2(n_80), .B(n_81), .C(n_83), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_731), .B(n_83), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_733), .Y(n_950) );
AO21x2_ASAP7_75t_L g951 ( .A1(n_714), .A2(n_191), .B(n_190), .Y(n_951) );
OAI21xp5_ASAP7_75t_L g952 ( .A1(n_815), .A2(n_194), .B(n_192), .Y(n_952) );
OAI21xp5_ASAP7_75t_L g953 ( .A1(n_771), .A2(n_200), .B(n_197), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_810), .B(n_84), .Y(n_954) );
AO221x2_ASAP7_75t_L g955 ( .A1(n_773), .A2(n_84), .B1(n_85), .B2(n_87), .C(n_88), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_793), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_757), .B(n_85), .Y(n_957) );
AOI21xp5_ASAP7_75t_L g958 ( .A1(n_724), .A2(n_205), .B(n_201), .Y(n_958) );
AOI21xp5_ASAP7_75t_L g959 ( .A1(n_724), .A2(n_212), .B(n_207), .Y(n_959) );
AOI221x1_ASAP7_75t_L g960 ( .A1(n_706), .A2(n_87), .B1(n_88), .B2(n_89), .C(n_90), .Y(n_960) );
BUFx8_ASAP7_75t_L g961 ( .A(n_718), .Y(n_961) );
A2O1A1Ixp33_ASAP7_75t_L g962 ( .A1(n_797), .A2(n_89), .B(n_90), .C(n_91), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_797), .B(n_91), .Y(n_963) );
A2O1A1Ixp33_ASAP7_75t_L g964 ( .A1(n_798), .A2(n_92), .B(n_93), .C(n_94), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_798), .A2(n_214), .B(n_213), .Y(n_965) );
OA21x2_ASAP7_75t_L g966 ( .A1(n_771), .A2(n_219), .B(n_218), .Y(n_966) );
INVx8_ASAP7_75t_L g967 ( .A(n_718), .Y(n_967) );
A2O1A1Ixp33_ASAP7_75t_L g968 ( .A1(n_718), .A2(n_92), .B(n_93), .C(n_95), .Y(n_968) );
AO21x2_ASAP7_75t_L g969 ( .A1(n_771), .A2(n_222), .B(n_220), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_771), .Y(n_970) );
A2O1A1Ixp33_ASAP7_75t_L g971 ( .A1(n_722), .A2(n_95), .B(n_96), .C(n_97), .Y(n_971) );
BUFx12f_ASAP7_75t_L g972 ( .A(n_722), .Y(n_972) );
OAI22x1_ASAP7_75t_L g973 ( .A1(n_781), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_973) );
NOR2xp33_ASAP7_75t_SL g974 ( .A(n_722), .B(n_98), .Y(n_974) );
AO32x2_ASAP7_75t_L g975 ( .A1(n_759), .A2(n_101), .A3(n_102), .B1(n_103), .B2(n_104), .Y(n_975) );
BUFx4f_ASAP7_75t_SL g976 ( .A(n_736), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_707), .B(n_102), .Y(n_977) );
O2A1O1Ixp33_ASAP7_75t_L g978 ( .A1(n_753), .A2(n_103), .B(n_105), .C(n_107), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_772), .A2(n_105), .B1(n_107), .B2(n_108), .Y(n_979) );
AO221x2_ASAP7_75t_L g980 ( .A1(n_742), .A2(n_108), .B1(n_109), .B2(n_110), .C(n_111), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_835), .Y(n_981) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_891), .A2(n_924), .B1(n_955), .B2(n_861), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_825), .Y(n_983) );
INVx2_ASAP7_75t_L g984 ( .A(n_822), .Y(n_984) );
AOI21xp5_ASAP7_75t_L g985 ( .A1(n_856), .A2(n_224), .B(n_223), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_841), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_873), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_905), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_881), .B(n_109), .Y(n_989) );
INVxp33_ASAP7_75t_L g990 ( .A(n_831), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_824), .Y(n_991) );
CKINVDCx11_ASAP7_75t_R g992 ( .A(n_847), .Y(n_992) );
NOR2xp33_ASAP7_75t_SL g993 ( .A(n_922), .B(n_110), .Y(n_993) );
AO31x2_ASAP7_75t_L g994 ( .A1(n_836), .A2(n_111), .A3(n_112), .B(n_113), .Y(n_994) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_942), .B(n_880), .Y(n_995) );
OA21x2_ASAP7_75t_L g996 ( .A1(n_879), .A2(n_270), .B(n_350), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_890), .B(n_114), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_924), .A2(n_114), .B1(n_115), .B2(n_116), .Y(n_998) );
CKINVDCx5p33_ASAP7_75t_R g999 ( .A(n_838), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_949), .Y(n_1000) );
OA21x2_ASAP7_75t_L g1001 ( .A1(n_896), .A2(n_268), .B(n_345), .Y(n_1001) );
INVx2_ASAP7_75t_L g1002 ( .A(n_912), .Y(n_1002) );
OAI221xp5_ASAP7_75t_SL g1003 ( .A1(n_916), .A2(n_115), .B1(n_116), .B2(n_117), .C(n_118), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_955), .A2(n_117), .B1(n_118), .B2(n_119), .Y(n_1004) );
OR2x2_ASAP7_75t_L g1005 ( .A(n_840), .B(n_121), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_923), .B(n_121), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_949), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_934), .B(n_122), .Y(n_1008) );
A2O1A1Ixp33_ASAP7_75t_L g1009 ( .A1(n_842), .A2(n_122), .B(n_124), .C(n_125), .Y(n_1009) );
INVx3_ASAP7_75t_L g1010 ( .A(n_972), .Y(n_1010) );
OA21x2_ASAP7_75t_L g1011 ( .A1(n_928), .A2(n_272), .B(n_340), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_900), .B(n_125), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_926), .Y(n_1013) );
BUFx3_ASAP7_75t_L g1014 ( .A(n_961), .Y(n_1014) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_961), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_941), .B(n_126), .Y(n_1016) );
OR2x2_ASAP7_75t_L g1017 ( .A(n_977), .B(n_127), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_904), .B(n_128), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_846), .B(n_128), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_858), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_845), .Y(n_1021) );
AND2x4_ASAP7_75t_L g1022 ( .A(n_829), .B(n_129), .Y(n_1022) );
AO21x2_ASAP7_75t_L g1023 ( .A1(n_863), .A2(n_273), .B(n_337), .Y(n_1023) );
A2O1A1Ixp33_ASAP7_75t_L g1024 ( .A1(n_876), .A2(n_129), .B(n_130), .C(n_131), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_864), .Y(n_1025) );
BUFx2_ASAP7_75t_L g1026 ( .A(n_916), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_980), .A2(n_130), .B1(n_131), .B2(n_132), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_909), .B(n_132), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_920), .B(n_133), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_829), .Y(n_1030) );
OAI221xp5_ASAP7_75t_L g1031 ( .A1(n_903), .A2(n_134), .B1(n_135), .B2(n_136), .C(n_137), .Y(n_1031) );
OA21x2_ASAP7_75t_L g1032 ( .A1(n_895), .A2(n_278), .B(n_336), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_865), .B(n_877), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_850), .Y(n_1034) );
A2O1A1Ixp33_ASAP7_75t_L g1035 ( .A1(n_978), .A2(n_135), .B(n_136), .C(n_137), .Y(n_1035) );
INVx3_ASAP7_75t_L g1036 ( .A(n_829), .Y(n_1036) );
INVx2_ASAP7_75t_L g1037 ( .A(n_950), .Y(n_1037) );
AO21x2_ASAP7_75t_L g1038 ( .A1(n_907), .A2(n_282), .B(n_334), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_940), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_887), .B(n_138), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_827), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_921), .Y(n_1042) );
OAI221xp5_ASAP7_75t_L g1043 ( .A1(n_832), .A2(n_139), .B1(n_140), .B2(n_142), .C(n_143), .Y(n_1043) );
INVx2_ASAP7_75t_SL g1044 ( .A(n_976), .Y(n_1044) );
INVx2_ASAP7_75t_L g1045 ( .A(n_893), .Y(n_1045) );
BUFx6f_ASAP7_75t_L g1046 ( .A(n_844), .Y(n_1046) );
NOR2x1_ASAP7_75t_SL g1047 ( .A(n_844), .B(n_139), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_894), .Y(n_1048) );
O2A1O1Ixp33_ASAP7_75t_L g1049 ( .A1(n_854), .A2(n_140), .B(n_143), .C(n_145), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_931), .Y(n_1050) );
NAND2xp33_ASAP7_75t_L g1051 ( .A(n_823), .B(n_146), .Y(n_1051) );
NAND2xp5_ASAP7_75t_SL g1052 ( .A(n_844), .B(n_147), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_980), .A2(n_148), .B1(n_150), .B2(n_152), .Y(n_1053) );
BUFx2_ASAP7_75t_L g1054 ( .A(n_859), .Y(n_1054) );
A2O1A1Ixp33_ASAP7_75t_L g1055 ( .A1(n_889), .A2(n_148), .B(n_152), .C(n_153), .Y(n_1055) );
AOI33xp33_ASAP7_75t_L g1056 ( .A1(n_843), .A2(n_153), .A3(n_226), .B1(n_227), .B2(n_229), .B3(n_232), .Y(n_1056) );
AOI21xp5_ASAP7_75t_L g1057 ( .A1(n_869), .A2(n_234), .B(n_235), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_899), .B(n_236), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1059 ( .A(n_823), .Y(n_1059) );
INVx2_ASAP7_75t_SL g1060 ( .A(n_830), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_944), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_852), .A2(n_237), .B1(n_238), .B2(n_239), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_938), .Y(n_1063) );
NAND3xp33_ASAP7_75t_L g1064 ( .A(n_943), .B(n_242), .C(n_244), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_918), .B(n_248), .Y(n_1065) );
INVx4_ASAP7_75t_L g1066 ( .A(n_967), .Y(n_1066) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_849), .B(n_249), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_872), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_871), .Y(n_1069) );
OR2x2_ASAP7_75t_L g1070 ( .A(n_883), .B(n_253), .Y(n_1070) );
INVx1_ASAP7_75t_SL g1071 ( .A(n_884), .Y(n_1071) );
INVx2_ASAP7_75t_L g1072 ( .A(n_878), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_828), .B(n_260), .Y(n_1073) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_823), .A2(n_262), .B1(n_264), .B2(n_265), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_898), .Y(n_1075) );
INVx3_ASAP7_75t_L g1076 ( .A(n_967), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_930), .Y(n_1077) );
AND2x2_ASAP7_75t_L g1078 ( .A(n_902), .B(n_271), .Y(n_1078) );
NOR2x1_ASAP7_75t_L g1079 ( .A(n_927), .B(n_276), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_930), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1081 ( .A1(n_945), .A2(n_285), .B1(n_286), .B2(n_287), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_862), .B(n_289), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_963), .Y(n_1083) );
OA21x2_ASAP7_75t_L g1084 ( .A1(n_914), .A2(n_290), .B(n_291), .Y(n_1084) );
BUFx3_ASAP7_75t_L g1085 ( .A(n_915), .Y(n_1085) );
OAI21x1_ASAP7_75t_L g1086 ( .A1(n_970), .A2(n_292), .B(n_296), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g1087 ( .A1(n_911), .A2(n_299), .B1(n_301), .B2(n_303), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_862), .B(n_305), .Y(n_1088) );
A2O1A1Ixp33_ASAP7_75t_L g1089 ( .A1(n_957), .A2(n_307), .B(n_309), .C(n_310), .Y(n_1089) );
INVx2_ASAP7_75t_L g1090 ( .A(n_886), .Y(n_1090) );
NOR2xp33_ASAP7_75t_L g1091 ( .A(n_939), .B(n_311), .Y(n_1091) );
BUFx4f_ASAP7_75t_SL g1092 ( .A(n_915), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_853), .B(n_312), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1094 ( .A1(n_839), .A2(n_314), .B1(n_315), .B2(n_316), .C(n_317), .Y(n_1094) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_956), .B(n_318), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_954), .A2(n_322), .B1(n_323), .B2(n_324), .Y(n_1096) );
NAND2xp5_ASAP7_75t_L g1097 ( .A(n_851), .B(n_325), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_823), .B(n_327), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_855), .B(n_330), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_885), .Y(n_1100) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_919), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_901), .A2(n_888), .B1(n_946), .B2(n_936), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_833), .B(n_332), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_837), .B(n_866), .Y(n_1104) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_882), .A2(n_979), .B1(n_917), .B2(n_952), .Y(n_1105) );
AOI21xp5_ASAP7_75t_L g1106 ( .A1(n_868), .A2(n_913), .B(n_935), .Y(n_1106) );
OAI211xp5_ASAP7_75t_L g1107 ( .A1(n_897), .A2(n_937), .B(n_929), .C(n_933), .Y(n_1107) );
OR2x6_ASAP7_75t_L g1108 ( .A(n_973), .B(n_953), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_837), .B(n_947), .Y(n_1109) );
AO31x2_ASAP7_75t_L g1110 ( .A1(n_960), .A2(n_870), .A3(n_910), .B(n_908), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g1111 ( .A(n_947), .B(n_892), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_932), .Y(n_1112) );
AO31x2_ASAP7_75t_L g1113 ( .A1(n_962), .A2(n_964), .A3(n_948), .B(n_971), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_857), .B(n_860), .Y(n_1114) );
A2O1A1Ixp33_ASAP7_75t_L g1115 ( .A1(n_968), .A2(n_826), .B(n_834), .C(n_965), .Y(n_1115) );
INVx3_ASAP7_75t_L g1116 ( .A(n_857), .Y(n_1116) );
O2A1O1Ixp33_ASAP7_75t_L g1117 ( .A1(n_874), .A2(n_925), .B(n_848), .C(n_974), .Y(n_1117) );
OAI22xp33_ASAP7_75t_L g1118 ( .A1(n_966), .A2(n_959), .B1(n_958), .B2(n_906), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1119 ( .A(n_857), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_906), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_906), .Y(n_1121) );
OAI21x1_ASAP7_75t_L g1122 ( .A1(n_966), .A2(n_867), .B(n_875), .Y(n_1122) );
OAI21x1_ASAP7_75t_L g1123 ( .A1(n_867), .A2(n_875), .B(n_886), .Y(n_1123) );
INVx11_ASAP7_75t_L g1124 ( .A(n_975), .Y(n_1124) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_837), .B(n_951), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_860), .B(n_875), .Y(n_1126) );
AO31x2_ASAP7_75t_L g1127 ( .A1(n_867), .A2(n_860), .A3(n_975), .B(n_969), .Y(n_1127) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_975), .A2(n_856), .B(n_723), .Y(n_1128) );
A2O1A1Ixp33_ASAP7_75t_L g1129 ( .A1(n_881), .A2(n_842), .B(n_876), .C(n_978), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_835), .Y(n_1130) );
INVx2_ASAP7_75t_L g1131 ( .A(n_825), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_942), .B(n_707), .Y(n_1132) );
A2O1A1Ixp33_ASAP7_75t_L g1133 ( .A1(n_881), .A2(n_842), .B(n_876), .C(n_978), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_835), .Y(n_1134) );
BUFx4f_ASAP7_75t_SL g1135 ( .A(n_847), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_891), .A2(n_765), .B1(n_817), .B2(n_801), .Y(n_1136) );
HB1xp67_ASAP7_75t_L g1137 ( .A(n_840), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_835), .Y(n_1138) );
AND2x4_ASAP7_75t_L g1139 ( .A(n_881), .B(n_825), .Y(n_1139) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_922), .A2(n_661), .B1(n_678), .B2(n_671), .Y(n_1140) );
OAI21xp5_ASAP7_75t_SL g1141 ( .A1(n_924), .A2(n_672), .B(n_671), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g1142 ( .A1(n_881), .A2(n_817), .B1(n_801), .B2(n_949), .Y(n_1142) );
BUFx3_ASAP7_75t_L g1143 ( .A(n_1014), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_991), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1139), .B(n_983), .Y(n_1145) );
INVxp67_ASAP7_75t_L g1146 ( .A(n_1137), .Y(n_1146) );
CKINVDCx5p33_ASAP7_75t_R g1147 ( .A(n_992), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_981), .Y(n_1148) );
AOI21xp5_ASAP7_75t_SL g1149 ( .A1(n_1142), .A2(n_1117), .B(n_1059), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_1139), .B(n_1131), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1151 ( .A1(n_982), .A2(n_1140), .B1(n_1108), .B2(n_1101), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1152 ( .A(n_1141), .B(n_1041), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_984), .B(n_1114), .Y(n_1153) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1019), .B(n_1025), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_988), .B(n_1002), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1156 ( .A(n_1020), .B(n_1045), .Y(n_1156) );
OR2x2_ASAP7_75t_L g1157 ( .A(n_1017), .B(n_1071), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1158 ( .A1(n_1141), .A2(n_1031), .B1(n_1068), .B2(n_1050), .C(n_1042), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1159 ( .A(n_1132), .Y(n_1159) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_1071), .B(n_1005), .Y(n_1160) );
INVx3_ASAP7_75t_L g1161 ( .A(n_1046), .Y(n_1161) );
INVx2_ASAP7_75t_SL g1162 ( .A(n_1015), .Y(n_1162) );
INVx3_ASAP7_75t_SL g1163 ( .A(n_1044), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1048), .B(n_1063), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1033), .B(n_987), .Y(n_1165) );
INVxp67_ASAP7_75t_L g1166 ( .A(n_1026), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_997), .B(n_1012), .Y(n_1167) );
OR2x6_ASAP7_75t_L g1168 ( .A(n_1108), .B(n_1142), .Y(n_1168) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_986), .B(n_1130), .Y(n_1169) );
AO21x2_ASAP7_75t_L g1170 ( .A1(n_1128), .A2(n_1126), .B(n_1118), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1134), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1072), .Y(n_1172) );
INVx4_ASAP7_75t_R g1173 ( .A(n_1060), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1138), .Y(n_1174) );
CKINVDCx20_ASAP7_75t_R g1175 ( .A(n_1135), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1033), .B(n_1037), .Y(n_1176) );
INVx4_ASAP7_75t_L g1177 ( .A(n_1046), .Y(n_1177) );
AOI21xp5_ASAP7_75t_SL g1178 ( .A1(n_1108), .A2(n_1098), .B(n_1055), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_989), .Y(n_1179) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_1010), .Y(n_1180) );
OAI21xp5_ASAP7_75t_SL g1181 ( .A1(n_1136), .A2(n_1004), .B(n_1027), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1061), .B(n_1053), .Y(n_1182) );
AOI21xp5_ASAP7_75t_SL g1183 ( .A1(n_1098), .A2(n_1047), .B(n_1022), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1116), .B(n_989), .Y(n_1184) );
OAI21xp5_ASAP7_75t_L g1185 ( .A1(n_1129), .A2(n_1133), .B(n_1115), .Y(n_1185) );
OR2x6_ASAP7_75t_L g1186 ( .A(n_1022), .B(n_1119), .Y(n_1186) );
INVx3_ASAP7_75t_L g1187 ( .A(n_1036), .Y(n_1187) );
AND2x4_ASAP7_75t_L g1188 ( .A(n_1036), .B(n_1000), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1007), .B(n_1030), .Y(n_1189) );
INVxp67_ASAP7_75t_L g1190 ( .A(n_1054), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1006), .Y(n_1191) );
AOI22xp5_ASAP7_75t_L g1192 ( .A1(n_1051), .A2(n_993), .B1(n_1083), .B2(n_995), .Y(n_1192) );
OR2x2_ASAP7_75t_SL g1193 ( .A(n_1013), .B(n_1067), .Y(n_1193) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_1107), .A2(n_1102), .B(n_1105), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1006), .Y(n_1195) );
NOR2x1p5_ASAP7_75t_L g1196 ( .A(n_999), .B(n_1010), .Y(n_1196) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1116), .B(n_1075), .Y(n_1197) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_1031), .A2(n_1043), .B1(n_1069), .B2(n_1039), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1008), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1008), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1040), .Y(n_1201) );
INVx3_ASAP7_75t_L g1202 ( .A(n_1066), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1120), .B(n_1121), .Y(n_1203) );
INVx2_ASAP7_75t_L g1204 ( .A(n_996), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1077), .B(n_1080), .Y(n_1205) );
OAI211xp5_ASAP7_75t_L g1206 ( .A1(n_1003), .A2(n_998), .B(n_1043), .C(n_1028), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1040), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1016), .Y(n_1208) );
AND2x4_ASAP7_75t_L g1209 ( .A(n_1109), .B(n_1021), .Y(n_1209) );
INVx2_ASAP7_75t_SL g1210 ( .A(n_1066), .Y(n_1210) );
AO21x2_ASAP7_75t_L g1211 ( .A1(n_1112), .A2(n_1106), .B(n_1109), .Y(n_1211) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_1100), .Y(n_1212) );
INVx2_ASAP7_75t_L g1213 ( .A(n_996), .Y(n_1213) );
BUFx3_ASAP7_75t_L g1214 ( .A(n_1076), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1018), .B(n_1078), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1016), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1018), .B(n_994), .Y(n_1217) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_1091), .A2(n_1028), .B1(n_1124), .B2(n_1104), .Y(n_1218) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_1029), .A2(n_1049), .B(n_1024), .C(n_1052), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_990), .B(n_1029), .Y(n_1220) );
INVx2_ASAP7_75t_L g1221 ( .A(n_1001), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_994), .Y(n_1222) );
OAI22xp5_ASAP7_75t_L g1223 ( .A1(n_1105), .A2(n_1097), .B1(n_1088), .B2(n_1082), .Y(n_1223) );
HB1xp67_ASAP7_75t_L g1224 ( .A(n_1076), .Y(n_1224) );
INVx5_ASAP7_75t_L g1225 ( .A(n_1125), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1085), .B(n_1099), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_993), .Y(n_1227) );
AND2x4_ASAP7_75t_SL g1228 ( .A(n_1111), .B(n_1074), .Y(n_1228) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1001), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1127), .B(n_1113), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1079), .Y(n_1231) );
NOR2xp33_ASAP7_75t_L g1232 ( .A(n_1092), .B(n_1099), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1009), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1127), .B(n_1113), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1058), .Y(n_1235) );
INVx2_ASAP7_75t_L g1236 ( .A(n_1084), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1034), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1056), .Y(n_1238) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1084), .Y(n_1239) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1127), .Y(n_1240) );
BUFx3_ASAP7_75t_L g1241 ( .A(n_1093), .Y(n_1241) );
AOI22xp5_ASAP7_75t_L g1242 ( .A1(n_1095), .A2(n_1097), .B1(n_1087), .B2(n_1094), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1035), .Y(n_1243) );
AND2x4_ASAP7_75t_L g1244 ( .A(n_1086), .B(n_1023), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1070), .Y(n_1245) );
AND2x4_ASAP7_75t_L g1246 ( .A(n_1023), .B(n_1113), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1065), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1110), .B(n_1032), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_1094), .A2(n_1064), .B1(n_1073), .B2(n_1103), .Y(n_1249) );
OR2x6_ASAP7_75t_L g1250 ( .A(n_985), .B(n_1057), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g1251 ( .A(n_1103), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1110), .B(n_1038), .Y(n_1252) );
BUFx2_ASAP7_75t_L g1253 ( .A(n_1038), .Y(n_1253) );
INVx1_ASAP7_75t_L g1254 ( .A(n_1089), .Y(n_1254) );
HB1xp67_ASAP7_75t_L g1255 ( .A(n_1011), .Y(n_1255) );
OA21x2_ASAP7_75t_L g1256 ( .A1(n_1096), .A2(n_1062), .B(n_1081), .Y(n_1256) );
OAI221xp5_ASAP7_75t_L g1257 ( .A1(n_1011), .A2(n_982), .B1(n_1141), .B2(n_672), .C(n_695), .Y(n_1257) );
OA21x2_ASAP7_75t_L g1258 ( .A1(n_1122), .A2(n_1123), .B(n_1128), .Y(n_1258) );
INVx2_ASAP7_75t_SL g1259 ( .A(n_1014), .Y(n_1259) );
INVxp67_ASAP7_75t_L g1260 ( .A(n_1137), .Y(n_1260) );
INVxp67_ASAP7_75t_L g1261 ( .A(n_1137), .Y(n_1261) );
AOI21xp5_ASAP7_75t_SL g1262 ( .A1(n_1142), .A2(n_1117), .B(n_949), .Y(n_1262) );
BUFx3_ASAP7_75t_L g1263 ( .A(n_1014), .Y(n_1263) );
OA21x2_ASAP7_75t_L g1264 ( .A1(n_1122), .A2(n_1123), .B(n_1128), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1141), .B(n_772), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1139), .B(n_983), .Y(n_1266) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1090), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1141), .B(n_772), .Y(n_1268) );
OA21x2_ASAP7_75t_L g1269 ( .A1(n_1122), .A2(n_1123), .B(n_1128), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1139), .B(n_983), .Y(n_1270) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1090), .Y(n_1271) );
BUFx3_ASAP7_75t_L g1272 ( .A(n_1014), .Y(n_1272) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1090), .Y(n_1273) );
AO21x2_ASAP7_75t_L g1274 ( .A1(n_1128), .A2(n_1126), .B(n_1118), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1137), .B(n_984), .Y(n_1275) );
INVx2_ASAP7_75t_SL g1276 ( .A(n_1014), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_991), .Y(n_1277) );
BUFx3_ASAP7_75t_L g1278 ( .A(n_1014), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_1159), .Y(n_1279) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_1257), .A2(n_1151), .B1(n_1192), .B2(n_1198), .Y(n_1280) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1205), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1205), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1153), .B(n_1217), .Y(n_1283) );
OAI21xp33_ASAP7_75t_L g1284 ( .A1(n_1151), .A2(n_1194), .B(n_1265), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1203), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1203), .Y(n_1286) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1162), .B(n_1259), .Y(n_1287) );
OR2x6_ASAP7_75t_L g1288 ( .A(n_1168), .B(n_1186), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1153), .B(n_1217), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1290 ( .A(n_1165), .B(n_1152), .Y(n_1290) );
INVx4_ASAP7_75t_L g1291 ( .A(n_1186), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1209), .B(n_1230), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1209), .B(n_1230), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1209), .B(n_1234), .Y(n_1294) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1197), .Y(n_1295) );
NAND2xp5_ASAP7_75t_L g1296 ( .A(n_1165), .B(n_1158), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1234), .B(n_1176), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1298 ( .A(n_1168), .B(n_1268), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1145), .B(n_1150), .Y(n_1299) );
BUFx2_ASAP7_75t_L g1300 ( .A(n_1186), .Y(n_1300) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1145), .B(n_1150), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1197), .Y(n_1302) );
AND2x4_ASAP7_75t_SL g1303 ( .A(n_1186), .B(n_1177), .Y(n_1303) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1176), .B(n_1184), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1172), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1184), .B(n_1168), .Y(n_1306) );
INVx2_ASAP7_75t_SL g1307 ( .A(n_1177), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1266), .B(n_1270), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1309 ( .A(n_1168), .B(n_1266), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_1270), .B(n_1155), .Y(n_1310) );
OAI22xp5_ASAP7_75t_L g1311 ( .A1(n_1198), .A2(n_1193), .B1(n_1241), .B2(n_1218), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1267), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1313 ( .A(n_1267), .B(n_1271), .Y(n_1313) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_1273), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1155), .B(n_1156), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1222), .Y(n_1316) );
BUFx2_ASAP7_75t_L g1317 ( .A(n_1225), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1156), .B(n_1164), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1164), .B(n_1170), .Y(n_1319) );
AND2x4_ASAP7_75t_L g1320 ( .A(n_1225), .B(n_1246), .Y(n_1320) );
INVxp67_ASAP7_75t_SL g1321 ( .A(n_1251), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1170), .B(n_1274), .Y(n_1322) );
INVxp67_ASAP7_75t_SL g1323 ( .A(n_1241), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1144), .B(n_1277), .Y(n_1324) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1148), .B(n_1171), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1274), .B(n_1174), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1185), .B(n_1240), .Y(n_1327) );
OAI211xp5_ASAP7_75t_L g1328 ( .A1(n_1181), .A2(n_1178), .B(n_1206), .C(n_1149), .Y(n_1328) );
OAI211xp5_ASAP7_75t_L g1329 ( .A1(n_1262), .A2(n_1232), .B(n_1166), .C(n_1220), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1237), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1225), .B(n_1215), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1215), .B(n_1252), .Y(n_1332) );
CKINVDCx20_ASAP7_75t_R g1333 ( .A(n_1175), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1252), .B(n_1179), .Y(n_1334) );
OR2x2_ASAP7_75t_L g1335 ( .A(n_1275), .B(n_1157), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1191), .B(n_1195), .Y(n_1336) );
BUFx2_ASAP7_75t_L g1337 ( .A(n_1177), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1169), .B(n_1199), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1200), .B(n_1167), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1211), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1201), .B(n_1207), .Y(n_1341) );
HB1xp67_ASAP7_75t_L g1342 ( .A(n_1146), .Y(n_1342) );
INVx2_ASAP7_75t_SL g1343 ( .A(n_1173), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1247), .B(n_1246), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1246), .B(n_1248), .Y(n_1345) );
NOR2x1_ASAP7_75t_L g1346 ( .A(n_1183), .B(n_1227), .Y(n_1346) );
OR2x2_ASAP7_75t_L g1347 ( .A(n_1160), .B(n_1154), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1208), .B(n_1216), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1258), .B(n_1264), .Y(n_1349) );
NAND2xp5_ASAP7_75t_L g1350 ( .A(n_1182), .B(n_1260), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1269), .B(n_1235), .Y(n_1351) );
OR2x6_ASAP7_75t_L g1352 ( .A(n_1223), .B(n_1250), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1269), .B(n_1189), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1189), .B(n_1238), .Y(n_1354) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1204), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1332), .B(n_1261), .Y(n_1356) );
NOR2xp67_ASAP7_75t_L g1357 ( .A(n_1343), .B(n_1162), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1315), .B(n_1182), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1330), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1330), .Y(n_1360) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_1280), .A2(n_1243), .B1(n_1233), .B2(n_1245), .Y(n_1361) );
OR2x2_ASAP7_75t_L g1362 ( .A(n_1335), .B(n_1190), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1324), .Y(n_1363) );
NAND2x1_ASAP7_75t_SL g1364 ( .A(n_1279), .B(n_1163), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1332), .B(n_1253), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1283), .B(n_1255), .Y(n_1366) );
INVx4_ASAP7_75t_L g1367 ( .A(n_1317), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1325), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1369 ( .A(n_1289), .B(n_1229), .Y(n_1369) );
BUFx3_ASAP7_75t_L g1370 ( .A(n_1337), .Y(n_1370) );
INVx2_ASAP7_75t_SL g1371 ( .A(n_1337), .Y(n_1371) );
INVxp67_ASAP7_75t_SL g1372 ( .A(n_1314), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1285), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1289), .B(n_1221), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1285), .Y(n_1375) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1297), .B(n_1221), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g1377 ( .A(n_1318), .B(n_1212), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1378 ( .A(n_1329), .B(n_1226), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1339), .B(n_1188), .Y(n_1379) );
AND2x4_ASAP7_75t_SL g1380 ( .A(n_1343), .B(n_1202), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1286), .Y(n_1381) );
INVxp67_ASAP7_75t_SL g1382 ( .A(n_1323), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1286), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1348), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1297), .B(n_1236), .Y(n_1385) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1281), .B(n_1180), .Y(n_1386) );
AND2x4_ASAP7_75t_L g1387 ( .A(n_1320), .B(n_1161), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1292), .B(n_1239), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1292), .B(n_1239), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1348), .Y(n_1390) );
INVx3_ASAP7_75t_SL g1391 ( .A(n_1333), .Y(n_1391) );
AND2x4_ASAP7_75t_L g1392 ( .A(n_1320), .B(n_1161), .Y(n_1392) );
OR2x2_ASAP7_75t_L g1393 ( .A(n_1304), .B(n_1276), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1293), .B(n_1294), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1294), .B(n_1213), .Y(n_1395) );
NOR2xp33_ASAP7_75t_L g1396 ( .A(n_1296), .B(n_1232), .Y(n_1396) );
OR2x2_ASAP7_75t_L g1397 ( .A(n_1347), .B(n_1259), .Y(n_1397) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_1347), .B(n_1180), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1336), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1336), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1401 ( .A(n_1339), .B(n_1188), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1341), .B(n_1310), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1334), .B(n_1244), .Y(n_1403) );
AND2x4_ASAP7_75t_L g1404 ( .A(n_1320), .B(n_1161), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1281), .B(n_1244), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1282), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1282), .B(n_1244), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1341), .Y(n_1408) );
AND2x4_ASAP7_75t_SL g1409 ( .A(n_1291), .B(n_1202), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1310), .B(n_1224), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_1295), .B(n_1302), .Y(n_1411) );
NAND2xp5_ASAP7_75t_L g1412 ( .A(n_1290), .B(n_1231), .Y(n_1412) );
AND2x2_ASAP7_75t_SL g1413 ( .A(n_1291), .B(n_1228), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1302), .B(n_1250), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1342), .Y(n_1415) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1299), .B(n_1278), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1417 ( .A(n_1301), .B(n_1278), .Y(n_1417) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1338), .B(n_1228), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1319), .B(n_1250), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1321), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1308), .Y(n_1421) );
NOR2xp67_ASAP7_75t_L g1422 ( .A(n_1328), .B(n_1202), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1423 ( .A(n_1284), .B(n_1210), .Y(n_1423) );
NAND2xp5_ASAP7_75t_L g1424 ( .A(n_1284), .B(n_1210), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1354), .Y(n_1425) );
INVx2_ASAP7_75t_L g1426 ( .A(n_1355), .Y(n_1426) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1326), .Y(n_1427) );
OR2x2_ASAP7_75t_L g1428 ( .A(n_1298), .B(n_1143), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1394), .B(n_1345), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1430 ( .A(n_1402), .B(n_1298), .Y(n_1430) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1394), .B(n_1345), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1420), .Y(n_1432) );
INVx1_ASAP7_75t_SL g1433 ( .A(n_1391), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1425), .B(n_1327), .Y(n_1434) );
INVx1_ASAP7_75t_SL g1435 ( .A(n_1391), .Y(n_1435) );
AOI21xp33_ASAP7_75t_L g1436 ( .A1(n_1378), .A2(n_1311), .B(n_1350), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1399), .B(n_1326), .Y(n_1437) );
OR2x2_ASAP7_75t_L g1438 ( .A(n_1356), .B(n_1313), .Y(n_1438) );
INVx1_ASAP7_75t_SL g1439 ( .A(n_1364), .Y(n_1439) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1359), .Y(n_1440) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1360), .Y(n_1441) );
AND2x4_ASAP7_75t_L g1442 ( .A(n_1419), .B(n_1288), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1443 ( .A(n_1356), .B(n_1313), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1403), .B(n_1319), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1415), .Y(n_1445) );
HB1xp67_ASAP7_75t_L g1446 ( .A(n_1372), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1400), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1408), .B(n_1344), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1403), .B(n_1353), .Y(n_1449) );
NOR2xp33_ASAP7_75t_L g1450 ( .A(n_1396), .B(n_1287), .Y(n_1450) );
AND2x4_ASAP7_75t_L g1451 ( .A(n_1419), .B(n_1288), .Y(n_1451) );
AOI22xp5_ASAP7_75t_L g1452 ( .A1(n_1361), .A2(n_1331), .B1(n_1352), .B2(n_1288), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1369), .B(n_1352), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1369), .B(n_1374), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1384), .B(n_1331), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1390), .Y(n_1456) );
INVx1_ASAP7_75t_L g1457 ( .A(n_1411), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1374), .B(n_1352), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1388), .B(n_1352), .Y(n_1459) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1421), .B(n_1351), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1363), .B(n_1351), .Y(n_1461) );
AND2x4_ASAP7_75t_L g1462 ( .A(n_1414), .B(n_1288), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1368), .B(n_1309), .Y(n_1463) );
AND2x4_ASAP7_75t_L g1464 ( .A(n_1414), .B(n_1288), .Y(n_1464) );
OAI21xp5_ASAP7_75t_L g1465 ( .A1(n_1422), .A2(n_1346), .B(n_1219), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1466 ( .A(n_1393), .B(n_1306), .Y(n_1466) );
OR2x2_ASAP7_75t_L g1467 ( .A(n_1377), .B(n_1306), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1373), .B(n_1309), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1388), .B(n_1352), .Y(n_1469) );
INVx2_ASAP7_75t_L g1470 ( .A(n_1426), .Y(n_1470) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1389), .B(n_1322), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1472 ( .A(n_1389), .B(n_1322), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1473 ( .A(n_1375), .B(n_1316), .Y(n_1473) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_1396), .A2(n_1291), .B1(n_1300), .B2(n_1254), .Y(n_1474) );
OR2x2_ASAP7_75t_L g1475 ( .A(n_1410), .B(n_1305), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1381), .Y(n_1476) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1366), .B(n_1312), .Y(n_1477) );
OR2x2_ASAP7_75t_L g1478 ( .A(n_1366), .B(n_1312), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1395), .B(n_1349), .Y(n_1479) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1383), .Y(n_1480) );
NAND2xp5_ASAP7_75t_SL g1481 ( .A(n_1439), .B(n_1357), .Y(n_1481) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1440), .Y(n_1482) );
NOR2xp33_ASAP7_75t_R g1483 ( .A(n_1433), .B(n_1147), .Y(n_1483) );
INVxp67_ASAP7_75t_L g1484 ( .A(n_1446), .Y(n_1484) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1441), .Y(n_1485) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1432), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1454), .B(n_1365), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1454), .B(n_1365), .Y(n_1488) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1446), .Y(n_1489) );
NAND2xp5_ASAP7_75t_L g1490 ( .A(n_1457), .B(n_1427), .Y(n_1490) );
AND2x4_ASAP7_75t_L g1491 ( .A(n_1442), .B(n_1405), .Y(n_1491) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1476), .Y(n_1492) );
OAI21xp5_ASAP7_75t_SL g1493 ( .A1(n_1465), .A2(n_1380), .B(n_1409), .Y(n_1493) );
BUFx3_ASAP7_75t_L g1494 ( .A(n_1435), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1480), .Y(n_1495) );
INVxp67_ASAP7_75t_SL g1496 ( .A(n_1470), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1477), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1429), .B(n_1376), .Y(n_1498) );
INVxp67_ASAP7_75t_SL g1499 ( .A(n_1478), .Y(n_1499) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1445), .Y(n_1500) );
OAI21xp5_ASAP7_75t_L g1501 ( .A1(n_1436), .A2(n_1378), .B(n_1424), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1429), .B(n_1376), .Y(n_1502) );
INVx2_ASAP7_75t_L g1503 ( .A(n_1447), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1504 ( .A(n_1434), .B(n_1412), .Y(n_1504) );
AOI22xp5_ASAP7_75t_L g1505 ( .A1(n_1450), .A2(n_1361), .B1(n_1413), .B2(n_1418), .Y(n_1505) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1461), .B(n_1406), .Y(n_1506) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1473), .Y(n_1507) );
NAND2xp5_ASAP7_75t_L g1508 ( .A(n_1437), .B(n_1405), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1431), .B(n_1385), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1510 ( .A(n_1460), .B(n_1407), .Y(n_1510) );
AND2x4_ASAP7_75t_L g1511 ( .A(n_1442), .B(n_1407), .Y(n_1511) );
INVx2_ASAP7_75t_L g1512 ( .A(n_1479), .Y(n_1512) );
INVx2_ASAP7_75t_L g1513 ( .A(n_1479), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1431), .B(n_1385), .Y(n_1514) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1438), .Y(n_1515) );
AOI21xp5_ASAP7_75t_L g1516 ( .A1(n_1493), .A2(n_1413), .B(n_1371), .Y(n_1516) );
OAI221xp5_ASAP7_75t_L g1517 ( .A1(n_1493), .A2(n_1474), .B1(n_1452), .B2(n_1450), .C(n_1423), .Y(n_1517) );
AND3x2_ASAP7_75t_L g1518 ( .A(n_1484), .B(n_1317), .C(n_1382), .Y(n_1518) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1503), .Y(n_1519) );
INVxp33_ASAP7_75t_L g1520 ( .A(n_1483), .Y(n_1520) );
INVxp67_ASAP7_75t_L g1521 ( .A(n_1494), .Y(n_1521) );
INVx2_ASAP7_75t_SL g1522 ( .A(n_1494), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1512), .B(n_1449), .Y(n_1523) );
AOI211xp5_ASAP7_75t_L g1524 ( .A1(n_1481), .A2(n_1501), .B(n_1494), .C(n_1505), .Y(n_1524) );
NAND2xp5_ASAP7_75t_SL g1525 ( .A(n_1505), .B(n_1367), .Y(n_1525) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1503), .Y(n_1526) );
AOI21xp5_ASAP7_75t_L g1527 ( .A1(n_1499), .A2(n_1371), .B(n_1367), .Y(n_1527) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1503), .Y(n_1528) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1482), .Y(n_1529) );
AOI222xp33_ASAP7_75t_L g1530 ( .A1(n_1504), .A2(n_1463), .B1(n_1456), .B2(n_1472), .C1(n_1471), .C2(n_1358), .Y(n_1530) );
AOI21xp33_ASAP7_75t_L g1531 ( .A1(n_1489), .A2(n_1428), .B(n_1397), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1482), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1489), .B(n_1471), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1485), .Y(n_1534) );
NAND2xp33_ASAP7_75t_L g1535 ( .A(n_1512), .B(n_1147), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1536 ( .A(n_1507), .B(n_1472), .Y(n_1536) );
NOR2xp33_ASAP7_75t_SL g1537 ( .A(n_1498), .B(n_1143), .Y(n_1537) );
NAND2xp5_ASAP7_75t_SL g1538 ( .A(n_1496), .B(n_1370), .Y(n_1538) );
AOI22xp5_ASAP7_75t_L g1539 ( .A1(n_1515), .A2(n_1453), .B1(n_1458), .B2(n_1459), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1507), .B(n_1444), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g1541 ( .A(n_1487), .B(n_1444), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1485), .Y(n_1542) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1523), .B(n_1512), .Y(n_1543) );
NAND2xp5_ASAP7_75t_L g1544 ( .A(n_1530), .B(n_1487), .Y(n_1544) );
AOI221xp5_ASAP7_75t_L g1545 ( .A1(n_1524), .A2(n_1515), .B1(n_1500), .B2(n_1497), .C(n_1486), .Y(n_1545) );
O2A1O1Ixp33_ASAP7_75t_L g1546 ( .A1(n_1525), .A2(n_1163), .B(n_1272), .C(n_1263), .Y(n_1546) );
O2A1O1Ixp33_ASAP7_75t_L g1547 ( .A1(n_1525), .A2(n_1272), .B(n_1263), .C(n_1500), .Y(n_1547) );
OAI222xp33_ASAP7_75t_L g1548 ( .A1(n_1517), .A2(n_1513), .B1(n_1497), .B2(n_1466), .C1(n_1467), .C2(n_1511), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1549 ( .A(n_1540), .B(n_1488), .Y(n_1549) );
INVxp67_ASAP7_75t_SL g1550 ( .A(n_1538), .Y(n_1550) );
INVxp67_ASAP7_75t_SL g1551 ( .A(n_1538), .Y(n_1551) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1529), .Y(n_1552) );
OAI21xp5_ASAP7_75t_L g1553 ( .A1(n_1520), .A2(n_1488), .B(n_1514), .Y(n_1553) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1519), .Y(n_1554) );
INVx1_ASAP7_75t_L g1555 ( .A(n_1526), .Y(n_1555) );
HB1xp67_ASAP7_75t_L g1556 ( .A(n_1522), .Y(n_1556) );
OAI21xp33_ASAP7_75t_L g1557 ( .A1(n_1537), .A2(n_1490), .B(n_1506), .Y(n_1557) );
AOI22xp33_ASAP7_75t_SL g1558 ( .A1(n_1535), .A2(n_1442), .B1(n_1451), .B2(n_1462), .Y(n_1558) );
NOR2x1_ASAP7_75t_L g1559 ( .A(n_1516), .B(n_1175), .Y(n_1559) );
AOI211xp5_ASAP7_75t_SL g1560 ( .A1(n_1521), .A2(n_1398), .B(n_1451), .C(n_1464), .Y(n_1560) );
NAND4xp25_ASAP7_75t_L g1561 ( .A(n_1559), .B(n_1527), .C(n_1539), .D(n_1531), .Y(n_1561) );
AOI22xp5_ASAP7_75t_L g1562 ( .A1(n_1545), .A2(n_1520), .B1(n_1536), .B2(n_1518), .Y(n_1562) );
AOI211x1_ASAP7_75t_SL g1563 ( .A1(n_1553), .A2(n_1533), .B(n_1541), .C(n_1513), .Y(n_1563) );
OAI21xp33_ASAP7_75t_L g1564 ( .A1(n_1550), .A2(n_1542), .B(n_1534), .Y(n_1564) );
A2O1A1Ixp33_ASAP7_75t_L g1565 ( .A1(n_1560), .A2(n_1409), .B(n_1513), .C(n_1509), .Y(n_1565) );
O2A1O1Ixp33_ASAP7_75t_L g1566 ( .A1(n_1548), .A2(n_1196), .B(n_1362), .C(n_1532), .Y(n_1566) );
OAI211xp5_ASAP7_75t_SL g1567 ( .A1(n_1546), .A2(n_1416), .B(n_1417), .C(n_1486), .Y(n_1567) );
OAI221xp5_ASAP7_75t_L g1568 ( .A1(n_1551), .A2(n_1492), .B1(n_1495), .B2(n_1528), .C(n_1430), .Y(n_1568) );
AOI32xp33_ASAP7_75t_L g1569 ( .A1(n_1558), .A2(n_1509), .A3(n_1498), .B1(n_1514), .B2(n_1502), .Y(n_1569) );
OAI211xp5_ASAP7_75t_L g1570 ( .A1(n_1547), .A2(n_1291), .B(n_1386), .C(n_1379), .Y(n_1570) );
AOI21xp33_ASAP7_75t_L g1571 ( .A1(n_1544), .A2(n_1492), .B(n_1495), .Y(n_1571) );
NAND2xp5_ASAP7_75t_SL g1572 ( .A(n_1557), .B(n_1370), .Y(n_1572) );
OAI211xp5_ASAP7_75t_L g1573 ( .A1(n_1556), .A2(n_1386), .B(n_1401), .C(n_1300), .Y(n_1573) );
OAI222xp33_ASAP7_75t_L g1574 ( .A1(n_1549), .A2(n_1511), .B1(n_1491), .B2(n_1508), .C1(n_1510), .C2(n_1443), .Y(n_1574) );
INVx2_ASAP7_75t_L g1575 ( .A(n_1572), .Y(n_1575) );
NAND3xp33_ASAP7_75t_SL g1576 ( .A(n_1563), .B(n_1518), .C(n_1552), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_1571), .B(n_1543), .Y(n_1577) );
AOI221xp5_ASAP7_75t_L g1578 ( .A1(n_1566), .A2(n_1555), .B1(n_1554), .B2(n_1543), .C(n_1502), .Y(n_1578) );
AOI211x1_ASAP7_75t_L g1579 ( .A1(n_1574), .A2(n_1561), .B(n_1570), .C(n_1564), .Y(n_1579) );
A2O1A1Ixp33_ASAP7_75t_SL g1580 ( .A1(n_1562), .A2(n_1569), .B(n_1568), .C(n_1567), .Y(n_1580) );
NAND3xp33_ASAP7_75t_SL g1581 ( .A(n_1565), .B(n_1242), .C(n_1554), .Y(n_1581) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1573), .B(n_1555), .Y(n_1582) );
NOR2xp33_ASAP7_75t_L g1583 ( .A(n_1572), .B(n_1491), .Y(n_1583) );
NOR2xp67_ASAP7_75t_L g1584 ( .A(n_1562), .B(n_1491), .Y(n_1584) );
AOI221xp5_ASAP7_75t_SL g1585 ( .A1(n_1578), .A2(n_1469), .B1(n_1468), .B2(n_1448), .C(n_1449), .Y(n_1585) );
NOR2xp33_ASAP7_75t_L g1586 ( .A(n_1575), .B(n_1475), .Y(n_1586) );
NOR2xp33_ASAP7_75t_L g1587 ( .A(n_1583), .B(n_1491), .Y(n_1587) );
NOR3xp33_ASAP7_75t_L g1588 ( .A(n_1580), .B(n_1214), .C(n_1187), .Y(n_1588) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1582), .Y(n_1589) );
NOR2x1_ASAP7_75t_L g1590 ( .A(n_1576), .B(n_1214), .Y(n_1590) );
NAND4xp25_ASAP7_75t_L g1591 ( .A(n_1579), .B(n_1249), .C(n_1464), .D(n_1462), .Y(n_1591) );
OAI22xp5_ASAP7_75t_SL g1592 ( .A1(n_1589), .A2(n_1577), .B1(n_1584), .B2(n_1581), .Y(n_1592) );
AO22x1_ASAP7_75t_L g1593 ( .A1(n_1588), .A2(n_1511), .B1(n_1307), .B2(n_1392), .Y(n_1593) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1586), .Y(n_1594) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1590), .Y(n_1595) );
NOR3xp33_ASAP7_75t_SL g1596 ( .A(n_1591), .B(n_1455), .C(n_1340), .Y(n_1596) );
XNOR2x1_ASAP7_75t_L g1597 ( .A(n_1594), .B(n_1585), .Y(n_1597) );
XNOR2xp5_ASAP7_75t_L g1598 ( .A(n_1592), .B(n_1587), .Y(n_1598) );
CKINVDCx20_ASAP7_75t_R g1599 ( .A(n_1595), .Y(n_1599) );
OAI22xp5_ASAP7_75t_SL g1600 ( .A1(n_1596), .A2(n_1256), .B1(n_1250), .B2(n_1404), .Y(n_1600) );
BUFx2_ASAP7_75t_L g1601 ( .A(n_1599), .Y(n_1601) );
INVxp67_ASAP7_75t_SL g1602 ( .A(n_1598), .Y(n_1602) );
AOI21xp5_ASAP7_75t_L g1603 ( .A1(n_1602), .A2(n_1597), .B(n_1600), .Y(n_1603) );
OA21x2_ASAP7_75t_L g1604 ( .A1(n_1601), .A2(n_1596), .B(n_1593), .Y(n_1604) );
OAI21xp33_ASAP7_75t_L g1605 ( .A1(n_1603), .A2(n_1303), .B(n_1404), .Y(n_1605) );
OR2x6_ASAP7_75t_L g1606 ( .A(n_1605), .B(n_1604), .Y(n_1606) );
AOI22xp5_ASAP7_75t_L g1607 ( .A1(n_1606), .A2(n_1387), .B1(n_1404), .B2(n_1392), .Y(n_1607) );
endmodule