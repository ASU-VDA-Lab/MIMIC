module fake_jpeg_27599_n_171 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

OR2x2_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_10),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx12_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_34),
.A2(n_21),
.B1(n_19),
.B2(n_24),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_37),
.B1(n_20),
.B2(n_31),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_17),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_14),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_51),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

NOR2x1_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_14),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_23),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_34),
.B1(n_37),
.B2(n_24),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_54),
.B1(n_60),
.B2(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_53),
.A2(n_57),
.B1(n_42),
.B2(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_70),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_1),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_25),
.C(n_26),
.Y(n_76)
);

BUFx24_ASAP7_75t_SL g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_27),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_14),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_70),
.B(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_80),
.B(n_28),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_63),
.B1(n_42),
.B2(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_48),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_81),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_46),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_44),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_14),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_94),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_67),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_102),
.Y(n_118)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_57),
.C(n_62),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_108),
.C(n_26),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_63),
.B(n_33),
.C(n_32),
.D(n_54),
.Y(n_98)
);

NOR4xp25_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_76),
.C(n_89),
.D(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_106),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_103),
.B(n_107),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_66),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_71),
.B(n_59),
.C(n_47),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_66),
.C(n_42),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_94),
.A2(n_86),
.B1(n_42),
.B2(n_72),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_115),
.B1(n_123),
.B2(n_26),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_105),
.B(n_87),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_28),
.B(n_18),
.C(n_15),
.D(n_23),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_109),
.B(n_90),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_91),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_125),
.C(n_108),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_91),
.B1(n_82),
.B2(n_75),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_115),
.B1(n_92),
.B2(n_119),
.Y(n_126)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_131),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_129),
.C(n_125),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_97),
.C(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

AOI221xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_98),
.B1(n_97),
.B2(n_84),
.C(n_28),
.Y(n_132)
);

AOI321xp33_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_138),
.A3(n_114),
.B1(n_28),
.B2(n_15),
.C(n_121),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_2),
.B(n_3),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_99),
.B1(n_47),
.B2(n_38),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_38),
.B1(n_118),
.B2(n_4),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_139),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_148),
.C(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_3),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_112),
.B(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_147),
.B1(n_137),
.B2(n_130),
.Y(n_150)
);

AOI31xp67_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_138),
.A3(n_127),
.B(n_129),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_13),
.C(n_12),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_144),
.B(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_153),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_152),
.B1(n_147),
.B2(n_146),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_154),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_159),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_155),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_148),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_152),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_11),
.C2(n_6),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_165),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_6),
.C(n_7),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_162),
.Y(n_167)
);

OAI21x1_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_160),
.B(n_9),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_166),
.A2(n_168),
.B(n_8),
.C(n_11),
.Y(n_170)
);


endmodule