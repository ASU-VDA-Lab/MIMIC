module real_aes_442_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_0), .B(n_180), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_1), .A2(n_188), .B(n_210), .Y(n_209) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_2), .A2(n_53), .B1(n_91), .B2(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_3), .B(n_195), .Y(n_258) );
INVx1_ASAP7_75t_L g164 ( .A(n_4), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g132 ( .A1(n_5), .A2(n_38), .B1(n_133), .B2(n_135), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_6), .B(n_195), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g107 ( .A1(n_7), .A2(n_16), .B1(n_108), .B2(n_113), .Y(n_107) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_8), .A2(n_24), .B1(n_91), .B2(n_100), .Y(n_99) );
NAND2xp33_ASAP7_75t_L g196 ( .A(n_9), .B(n_197), .Y(n_196) );
INVx2_ASAP7_75t_L g177 ( .A(n_10), .Y(n_177) );
AOI221x1_ASAP7_75t_L g274 ( .A1(n_11), .A2(n_21), .B1(n_180), .B2(n_188), .C(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_12), .B(n_180), .Y(n_179) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_13), .A2(n_175), .B(n_178), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_14), .B(n_213), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g87 ( .A1(n_15), .A2(n_62), .B1(n_88), .B2(n_104), .Y(n_87) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_17), .B(n_195), .Y(n_222) );
INVx1_ASAP7_75t_L g515 ( .A(n_17), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_18), .A2(n_61), .B1(n_122), .B2(n_123), .Y(n_121) );
AO21x1_ASAP7_75t_L g253 ( .A1(n_19), .A2(n_180), .B(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_20), .A2(n_74), .B1(n_141), .B2(n_142), .Y(n_140) );
NAND2x1_ASAP7_75t_L g244 ( .A(n_22), .B(n_195), .Y(n_244) );
NAND2x1_ASAP7_75t_L g232 ( .A(n_23), .B(n_197), .Y(n_232) );
OAI221xp5_ASAP7_75t_L g156 ( .A1(n_24), .A2(n_53), .B1(n_57), .B2(n_157), .C(n_159), .Y(n_156) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_25), .A2(n_65), .B(n_177), .Y(n_176) );
OR2x2_ASAP7_75t_L g200 ( .A(n_25), .B(n_65), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_26), .A2(n_148), .B1(n_149), .B2(n_150), .Y(n_147) );
INVxp67_ASAP7_75t_L g150 ( .A(n_26), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_27), .B(n_197), .Y(n_212) );
INVx3_ASAP7_75t_L g91 ( .A(n_28), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_29), .B(n_195), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_30), .A2(n_45), .B1(n_138), .B2(n_139), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_31), .B(n_197), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_32), .A2(n_188), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_SL g96 ( .A(n_33), .Y(n_96) );
INVx1_ASAP7_75t_L g166 ( .A(n_34), .Y(n_166) );
AND2x2_ASAP7_75t_L g186 ( .A(n_34), .B(n_164), .Y(n_186) );
AND2x2_ASAP7_75t_L g189 ( .A(n_34), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_35), .B(n_180), .Y(n_267) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_36), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_37), .B(n_197), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_39), .A2(n_188), .B(n_231), .Y(n_230) );
AO22x2_ASAP7_75t_L g90 ( .A1(n_40), .A2(n_57), .B1(n_91), .B2(n_92), .Y(n_90) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_41), .B(n_197), .Y(n_245) );
INVx1_ASAP7_75t_L g183 ( .A(n_42), .Y(n_183) );
INVx1_ASAP7_75t_L g192 ( .A(n_42), .Y(n_192) );
INVx1_ASAP7_75t_L g149 ( .A(n_43), .Y(n_149) );
INVx1_ASAP7_75t_L g97 ( .A(n_44), .Y(n_97) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_46), .B(n_195), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_47), .B(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_48), .A2(n_188), .B(n_243), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_49), .A2(n_64), .B1(n_129), .B2(n_130), .Y(n_128) );
AO21x1_ASAP7_75t_L g255 ( .A1(n_50), .A2(n_188), .B(n_256), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_51), .A2(n_145), .B1(n_146), .B2(n_147), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_51), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_51), .B(n_180), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_52), .B(n_180), .Y(n_234) );
INVxp33_ASAP7_75t_L g161 ( .A(n_53), .Y(n_161) );
AND2x2_ASAP7_75t_L g268 ( .A(n_54), .B(n_214), .Y(n_268) );
INVx1_ASAP7_75t_L g185 ( .A(n_55), .Y(n_185) );
INVx1_ASAP7_75t_L g190 ( .A(n_55), .Y(n_190) );
AND2x2_ASAP7_75t_L g236 ( .A(n_56), .B(n_205), .Y(n_236) );
INVxp67_ASAP7_75t_L g160 ( .A(n_57), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g143 ( .A1(n_58), .A2(n_144), .B1(n_151), .B2(n_152), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_58), .Y(n_151) );
AND2x2_ASAP7_75t_L g204 ( .A(n_59), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_60), .B(n_180), .Y(n_224) );
INVx1_ASAP7_75t_L g497 ( .A(n_60), .Y(n_497) );
AND2x2_ASAP7_75t_L g254 ( .A(n_63), .B(n_199), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_66), .B(n_197), .Y(n_223) );
AND2x2_ASAP7_75t_L g248 ( .A(n_67), .B(n_205), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_68), .B(n_195), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_69), .A2(n_188), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_70), .B(n_197), .Y(n_276) );
INVx1_ASAP7_75t_L g81 ( .A(n_71), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_72), .B(n_195), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_73), .A2(n_82), .B1(n_83), .B2(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_73), .Y(n_505) );
BUFx2_ASAP7_75t_SL g158 ( .A(n_75), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_76), .A2(n_188), .B(n_193), .Y(n_187) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_153), .B1(n_167), .B2(n_489), .C(n_494), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_143), .Y(n_78) );
AOI22xp33_ASAP7_75t_SL g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_82), .A2(n_83), .B1(n_496), .B2(n_497), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
NAND2x1_ASAP7_75t_SL g84 ( .A(n_85), .B(n_126), .Y(n_84) );
NOR2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_116), .Y(n_85) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_107), .Y(n_86) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_98), .Y(n_88) );
AND2x2_ASAP7_75t_L g129 ( .A(n_89), .B(n_109), .Y(n_129) );
AND2x6_ASAP7_75t_L g138 ( .A(n_89), .B(n_119), .Y(n_138) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_93), .Y(n_89) );
AND2x2_ASAP7_75t_L g106 ( .A(n_90), .B(n_94), .Y(n_106) );
INVx2_ASAP7_75t_L g112 ( .A(n_90), .Y(n_112) );
BUFx2_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
INVx1_ASAP7_75t_L g92 ( .A(n_91), .Y(n_92) );
OAI22x1_ASAP7_75t_L g94 ( .A1(n_91), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_91), .Y(n_95) );
INVx2_ASAP7_75t_L g100 ( .A(n_91), .Y(n_100) );
INVx1_ASAP7_75t_L g103 ( .A(n_91), .Y(n_103) );
AND2x4_ASAP7_75t_L g134 ( .A(n_93), .B(n_112), .Y(n_134) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
AND2x2_ASAP7_75t_L g111 ( .A(n_94), .B(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_94), .Y(n_124) );
AND2x4_ASAP7_75t_L g122 ( .A(n_98), .B(n_111), .Y(n_122) );
AND2x2_ASAP7_75t_L g135 ( .A(n_98), .B(n_134), .Y(n_135) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g110 ( .A(n_99), .Y(n_110) );
INVx1_ASAP7_75t_L g120 ( .A(n_99), .Y(n_120) );
AND2x2_ASAP7_75t_L g125 ( .A(n_99), .B(n_102), .Y(n_125) );
INVxp67_ASAP7_75t_L g105 ( .A(n_101), .Y(n_105) );
AND2x4_ASAP7_75t_L g119 ( .A(n_101), .B(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g109 ( .A(n_102), .B(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g113 ( .A(n_106), .B(n_114), .Y(n_113) );
AND2x4_ASAP7_75t_L g118 ( .A(n_106), .B(n_119), .Y(n_118) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x6_ASAP7_75t_L g139 ( .A(n_109), .B(n_134), .Y(n_139) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_110), .Y(n_115) );
AND2x2_ASAP7_75t_L g141 ( .A(n_111), .B(n_119), .Y(n_141) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
AND2x2_ASAP7_75t_L g133 ( .A(n_119), .B(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_SL g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x4_ASAP7_75t_L g130 ( .A(n_125), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g142 ( .A(n_125), .B(n_134), .Y(n_142) );
NOR2x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_136), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_132), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_140), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g152 ( .A(n_144), .Y(n_152) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_154), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_155), .Y(n_154) );
AND3x1_ASAP7_75t_SL g155 ( .A(n_156), .B(n_162), .C(n_165), .Y(n_155) );
INVxp67_ASAP7_75t_L g503 ( .A(n_156), .Y(n_503) );
CKINVDCx8_ASAP7_75t_R g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_162), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_162), .A2(n_511), .B(n_512), .Y(n_510) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_SL g508 ( .A(n_163), .B(n_165), .Y(n_508) );
AND2x2_ASAP7_75t_L g513 ( .A(n_163), .B(n_514), .Y(n_513) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g191 ( .A(n_164), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_165), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2x1p5_ASAP7_75t_L g491 ( .A(n_166), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_410), .Y(n_168) );
NOR3xp33_ASAP7_75t_SL g169 ( .A(n_170), .B(n_322), .C(n_362), .Y(n_169) );
OAI221xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_237), .B1(n_286), .B2(n_301), .C(n_304), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_173), .B(n_201), .Y(n_172) );
INVx2_ASAP7_75t_L g319 ( .A(n_173), .Y(n_319) );
AND2x2_ASAP7_75t_L g349 ( .A(n_173), .B(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g287 ( .A(n_174), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g294 ( .A(n_174), .B(n_227), .Y(n_294) );
INVx2_ASAP7_75t_L g300 ( .A(n_174), .Y(n_300) );
AND2x2_ASAP7_75t_L g309 ( .A(n_174), .B(n_203), .Y(n_309) );
INVx1_ASAP7_75t_L g325 ( .A(n_174), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_174), .B(n_371), .Y(n_370) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx3_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
AND2x4_ASAP7_75t_L g199 ( .A(n_177), .B(n_200), .Y(n_199) );
AND2x2_ASAP7_75t_SL g214 ( .A(n_177), .B(n_200), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_187), .B(n_199), .Y(n_178) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_186), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_182), .B(n_184), .Y(n_181) );
AND2x6_ASAP7_75t_L g197 ( .A(n_182), .B(n_190), .Y(n_197) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x4_ASAP7_75t_L g195 ( .A(n_184), .B(n_192), .Y(n_195) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx5_ASAP7_75t_L g198 ( .A(n_186), .Y(n_198) );
AND2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_191), .Y(n_188) );
INVx2_ASAP7_75t_L g493 ( .A(n_190), .Y(n_493) );
AND2x4_ASAP7_75t_L g490 ( .A(n_191), .B(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g514 ( .A(n_192), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .B(n_198), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_198), .A2(n_211), .B(n_212), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_198), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_232), .B(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_198), .A2(n_244), .B(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_198), .A2(n_257), .B(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_198), .A2(n_265), .B(n_266), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_198), .A2(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_SL g218 ( .A(n_199), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_199), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_202), .B(n_215), .Y(n_201) );
INVx4_ASAP7_75t_L g290 ( .A(n_202), .Y(n_290) );
AND2x2_ASAP7_75t_L g321 ( .A(n_202), .B(n_228), .Y(n_321) );
AND2x2_ASAP7_75t_L g397 ( .A(n_202), .B(n_371), .Y(n_397) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_202), .B(n_227), .Y(n_439) );
INVx5_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_203), .B(n_227), .Y(n_326) );
AND2x2_ASAP7_75t_L g350 ( .A(n_203), .B(n_228), .Y(n_350) );
BUFx2_ASAP7_75t_L g366 ( .A(n_203), .Y(n_366) );
NOR2x1_ASAP7_75t_SL g469 ( .A(n_203), .B(n_371), .Y(n_469) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_207), .Y(n_203) );
INVx3_ASAP7_75t_L g247 ( .A(n_205), .Y(n_247) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_213), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_213), .Y(n_235) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_213), .A2(n_274), .B(n_278), .Y(n_273) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_213), .A2(n_274), .B(n_278), .Y(n_336) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g346 ( .A(n_215), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_215), .A2(n_413), .B1(n_415), .B2(n_417), .C(n_422), .Y(n_412) );
AND2x2_ASAP7_75t_L g432 ( .A(n_215), .B(n_325), .Y(n_432) );
AND2x4_ASAP7_75t_L g215 ( .A(n_216), .B(n_227), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g288 ( .A(n_217), .Y(n_288) );
INVx1_ASAP7_75t_L g341 ( .A(n_217), .Y(n_341) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_218), .B(n_226), .Y(n_225) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_227), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g310 ( .A(n_227), .B(n_298), .Y(n_310) );
INVx2_ASAP7_75t_L g352 ( .A(n_227), .Y(n_352) );
AND2x2_ASAP7_75t_L g485 ( .A(n_227), .B(n_300), .Y(n_485) );
INVx4_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_228), .Y(n_342) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_235), .B(n_236), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_234), .Y(n_229) );
NOR3xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_269), .C(n_284), .Y(n_237) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_249), .Y(n_238) );
INVx2_ASAP7_75t_L g399 ( .A(n_239), .Y(n_399) );
AND2x2_ASAP7_75t_L g444 ( .A(n_239), .B(n_321), .Y(n_444) );
BUFx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g389 ( .A(n_240), .Y(n_389) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_240), .B(n_316), .Y(n_404) );
AO21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_247), .B(n_248), .Y(n_240) );
AO21x2_ASAP7_75t_L g283 ( .A1(n_241), .A2(n_247), .B(n_248), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_246), .Y(n_241) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_247), .A2(n_262), .B(n_268), .Y(n_261) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_247), .A2(n_262), .B(n_268), .Y(n_281) );
INVx2_ASAP7_75t_L g358 ( .A(n_249), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_249), .B(n_388), .Y(n_414) );
AND2x4_ASAP7_75t_L g447 ( .A(n_249), .B(n_394), .Y(n_447) );
AND2x4_ASAP7_75t_L g249 ( .A(n_250), .B(n_261), .Y(n_249) );
AND2x2_ASAP7_75t_L g285 ( .A(n_250), .B(n_280), .Y(n_285) );
OR2x2_ASAP7_75t_L g315 ( .A(n_250), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_250), .B(n_336), .Y(n_384) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
BUFx2_ASAP7_75t_L g329 ( .A(n_251), .Y(n_329) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g303 ( .A(n_252), .Y(n_303) );
OAI21x1_ASAP7_75t_SL g252 ( .A1(n_253), .A2(n_255), .B(n_259), .Y(n_252) );
INVx1_ASAP7_75t_L g260 ( .A(n_254), .Y(n_260) );
INVx2_ASAP7_75t_L g316 ( .A(n_261), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_263), .B(n_267), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_269), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_279), .Y(n_270) );
AND2x2_ASAP7_75t_L g284 ( .A(n_271), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g357 ( .A(n_271), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g442 ( .A(n_271), .Y(n_442) );
BUFx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x4_ASAP7_75t_L g302 ( .A(n_272), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g421 ( .A(n_272), .B(n_281), .Y(n_421) );
AND2x2_ASAP7_75t_L g425 ( .A(n_272), .B(n_291), .Y(n_425) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g394 ( .A(n_273), .Y(n_394) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_273), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_279), .B(n_302), .Y(n_378) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_280), .B(n_303), .Y(n_488) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g292 ( .A(n_281), .B(n_283), .Y(n_292) );
AND2x2_ASAP7_75t_L g374 ( .A(n_281), .B(n_336), .Y(n_374) );
AND2x2_ASAP7_75t_L g393 ( .A(n_281), .B(n_282), .Y(n_393) );
BUFx2_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_282), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx3_ASAP7_75t_L g291 ( .A(n_283), .Y(n_291) );
INVxp67_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
INVx1_ASAP7_75t_L g307 ( .A(n_285), .Y(n_307) );
AND2x2_ASAP7_75t_L g343 ( .A(n_285), .B(n_314), .Y(n_343) );
NAND2xp33_ASAP7_75t_L g424 ( .A(n_285), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g461 ( .A(n_285), .B(n_462), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_289), .B1(n_292), .B2(n_293), .C(n_295), .Y(n_286) );
AND2x2_ASAP7_75t_L g390 ( .A(n_287), .B(n_290), .Y(n_390) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_287), .B(n_350), .Y(n_409) );
AND2x2_ASAP7_75t_L g427 ( .A(n_287), .B(n_352), .Y(n_427) );
AND2x2_ASAP7_75t_L g482 ( .A(n_287), .B(n_321), .Y(n_482) );
INVx1_ASAP7_75t_L g298 ( .A(n_288), .Y(n_298) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_288), .Y(n_354) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_289), .Y(n_434) );
AND2x4_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_290), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_290), .B(n_341), .Y(n_416) );
AND2x2_ASAP7_75t_L g383 ( .A(n_291), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g419 ( .A(n_291), .Y(n_419) );
AND2x2_ASAP7_75t_L g328 ( .A(n_292), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_292), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g470 ( .A(n_292), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_292), .B(n_394), .Y(n_480) );
AND2x4_ASAP7_75t_L g396 ( .A(n_293), .B(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g467 ( .A(n_294), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OR2x2_ASAP7_75t_L g338 ( .A(n_299), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g345 ( .A(n_300), .B(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g376 ( .A(n_300), .B(n_350), .Y(n_376) );
AND2x2_ASAP7_75t_L g450 ( .A(n_300), .B(n_371), .Y(n_450) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g398 ( .A(n_302), .B(n_399), .Y(n_398) );
OAI32xp33_ASAP7_75t_L g463 ( .A1(n_302), .A2(n_464), .A3(n_466), .B1(n_467), .B2(n_470), .Y(n_463) );
AND2x4_ASAP7_75t_L g335 ( .A(n_303), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g433 ( .A(n_303), .B(n_336), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_308), .B1(n_311), .B2(n_317), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_SL g422 ( .A1(n_306), .A2(n_320), .B(n_423), .C(n_424), .Y(n_422) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g406 ( .A(n_307), .B(n_334), .Y(n_406) );
INVx1_ASAP7_75t_SL g477 ( .A(n_308), .Y(n_477) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x4_ASAP7_75t_L g380 ( .A(n_310), .B(n_319), .Y(n_380) );
AOI221xp5_ASAP7_75t_L g458 ( .A1(n_310), .A2(n_459), .B1(n_460), .B2(n_461), .C(n_463), .Y(n_458) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_315), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_318), .A2(n_348), .B1(n_401), .B2(n_402), .Y(n_400) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
OAI211xp5_ASAP7_75t_SL g436 ( .A1(n_319), .A2(n_437), .B(n_445), .C(n_458), .Y(n_436) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g356 ( .A(n_321), .B(n_325), .Y(n_356) );
OAI211xp5_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_327), .B(n_330), .C(n_359), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g353 ( .A(n_325), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g473 ( .A(n_325), .B(n_469), .Y(n_473) );
OAI32xp33_ASAP7_75t_L g430 ( .A1(n_326), .A2(n_431), .A3(n_433), .B1(n_434), .B2(n_435), .Y(n_430) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_SL g420 ( .A(n_329), .B(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_337), .B1(n_343), .B2(n_344), .C(n_347), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_333), .B(n_335), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g487 ( .A(n_334), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_335), .B(n_399), .Y(n_401) );
A2O1A1O1Ixp25_ASAP7_75t_L g472 ( .A1(n_335), .A2(n_404), .B(n_420), .C(n_466), .D(n_473), .Y(n_472) );
AOI31xp33_ASAP7_75t_L g474 ( .A1(n_335), .A2(n_356), .A3(n_466), .B(n_473), .Y(n_474) );
AND2x2_ASAP7_75t_L g388 ( .A(n_336), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_338), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx2_ASAP7_75t_L g465 ( .A(n_340), .Y(n_465) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g460 ( .A(n_341), .B(n_352), .Y(n_460) );
INVx1_ASAP7_75t_L g375 ( .A(n_343), .Y(n_375) );
AND2x2_ASAP7_75t_L g360 ( .A(n_344), .B(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI31xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_351), .A3(n_355), .B(n_357), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_350), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g483 ( .A(n_350), .B(n_429), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x2_ASAP7_75t_L g428 ( .A(n_352), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g454 ( .A(n_352), .Y(n_454) );
INVxp67_ASAP7_75t_L g423 ( .A(n_353), .Y(n_423) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g361 ( .A(n_357), .Y(n_361) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND3xp33_ASAP7_75t_SL g362 ( .A(n_363), .B(n_379), .C(n_395), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_372), .B1(n_376), .B2(n_377), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx2_ASAP7_75t_L g449 ( .A(n_366), .Y(n_449) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_SL g429 ( .A(n_370), .Y(n_429) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_370), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_370), .B(n_439), .Y(n_456) );
NAND2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx1_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_381), .B1(n_390), .B2(n_391), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_382), .B(n_385), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_388), .A2(n_393), .B1(n_427), .B2(n_428), .C(n_430), .Y(n_426) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g466 ( .A(n_393), .Y(n_466) );
AND2x2_ASAP7_75t_L g403 ( .A(n_394), .B(n_404), .Y(n_403) );
O2A1O1Ixp33_ASAP7_75t_SL g451 ( .A1(n_394), .A2(n_452), .B(n_456), .C(n_457), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B(n_400), .C(n_405), .Y(n_395) );
AND2x2_ASAP7_75t_L g446 ( .A(n_399), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g457 ( .A(n_404), .Y(n_457) );
AOI21xp33_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B(n_408), .Y(n_405) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_436), .C(n_471), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g411 ( .A(n_412), .B(n_426), .Y(n_411) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g435 ( .A(n_420), .Y(n_435) );
INVxp67_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_SL g443 ( .A(n_433), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_443), .B2(n_444), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_451), .Y(n_445) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g484 ( .A(n_469), .B(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_474), .B1(n_475), .B2(n_478), .C(n_481), .Y(n_471) );
INVxp67_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI31xp33_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_483), .A3(n_484), .B(n_486), .Y(n_481) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_491), .Y(n_511) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI222xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_498), .B1(n_504), .B2(n_506), .C1(n_509), .C2(n_515), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
endmodule