module real_jpeg_30366_n_13 (n_5, n_4, n_8, n_0, n_12, n_497, n_498, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_497;
input n_498;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_0),
.Y(n_174)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_1),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_1),
.Y(n_466)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_2),
.B(n_183),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_62),
.B1(n_193),
.B2(n_197),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_2),
.A2(n_62),
.B1(n_485),
.B2(n_488),
.Y(n_484)
);

INVx3_ASAP7_75t_R g69 ( 
.A(n_3),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_3),
.A2(n_56),
.B1(n_69),
.B2(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_3),
.A2(n_69),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_3),
.B(n_111),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_99),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_3),
.B(n_393),
.C(n_396),
.Y(n_392)
);

NAND2xp67_ASAP7_75t_L g408 ( 
.A(n_3),
.B(n_409),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_3),
.B(n_26),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_4),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_5),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_6),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_6),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_7),
.B(n_466),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_8),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_9),
.Y(n_114)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_9),
.Y(n_306)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_11),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_11),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_12),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_12),
.A2(n_104),
.B1(n_148),
.B2(n_152),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_12),
.A2(n_104),
.B1(n_233),
.B2(n_237),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g454 ( 
.A1(n_12),
.A2(n_104),
.B1(n_455),
.B2(n_458),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_472),
.B(n_493),
.Y(n_13)
);

OAI32xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_247),
.A3(n_439),
.B1(n_467),
.B2(n_497),
.Y(n_14)
);

OAI321xp33_ASAP7_75t_L g494 ( 
.A1(n_15),
.A2(n_247),
.A3(n_441),
.B1(n_467),
.B2(n_473),
.C(n_498),
.Y(n_494)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp67_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_205),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_18),
.B(n_469),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_185),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_19),
.B(n_185),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_144),
.C(n_157),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_21),
.A2(n_144),
.B1(n_145),
.B2(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_21),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_108),
.B2(n_143),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_66),
.B2(n_67),
.Y(n_23)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_24),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_25),
.B(n_190),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_42),
.B(n_60),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_26),
.A2(n_42),
.B1(n_60),
.B2(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_26),
.B(n_147),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_26),
.A2(n_147),
.B(n_161),
.Y(n_261)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_28),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B1(n_36),
.B2(n_38),
.Y(n_28)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_29),
.Y(n_175)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_29),
.Y(n_238)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_31),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_31),
.Y(n_236)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_35),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_37),
.Y(n_183)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp67_ASAP7_75t_L g161 ( 
.A(n_43),
.B(n_162),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_44),
.A2(n_163),
.B(n_223),
.Y(n_222)
);

OAI22x1_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B1(n_53),
.B2(n_56),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_52),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_52),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_52),
.Y(n_353)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_59),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_62),
.A2(n_177),
.B(n_182),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_67),
.B(n_184),
.C(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_80),
.B1(n_99),
.B2(n_100),
.Y(n_67)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_68),
.A2(n_80),
.B(n_81),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_75),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_69),
.A2(n_136),
.B(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_69),
.B(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_73),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_74),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_75),
.Y(n_368)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_91),
.B1(n_94),
.B2(n_98),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_79),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_80),
.Y(n_200)
);

NOR2x1p5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OAI22x1_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_89),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_84),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_84),
.Y(n_362)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_108),
.B(n_443),
.C(n_445),
.Y(n_442)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

AOI22x1_ASAP7_75t_L g211 ( 
.A1(n_109),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_211)
);

NOR2x1p5_ASAP7_75t_L g242 ( 
.A(n_109),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_109),
.B(n_222),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_110),
.Y(n_215)
);

AO22x2_ASAP7_75t_L g255 ( 
.A1(n_110),
.A2(n_156),
.B1(n_215),
.B2(n_256),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_122),
.B(n_135),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g452 ( 
.A(n_111),
.B(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_111),
.Y(n_460)
);

OAI22x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_115),
.B1(n_118),
.B2(n_120),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_114),
.Y(n_295)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_122),
.Y(n_453)
);

NAND2x1_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_127),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_127),
.Y(n_487)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_133),
.Y(n_302)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_134),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_135),
.Y(n_451)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp33_ASAP7_75t_L g312 ( 
.A(n_139),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_158),
.B1(n_167),
.B2(n_184),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_188),
.B1(n_189),
.B2(n_202),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_143),
.B(n_204),
.C(n_462),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_144),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_155),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_155),
.B(n_222),
.Y(n_333)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_215),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g256 ( 
.A(n_156),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_156),
.B(n_222),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_157),
.B(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2x1_ASAP7_75t_SL g210 ( 
.A(n_159),
.B(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_166),
.B(n_167),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_167),
.A2(n_213),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

NAND2x1_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OR2x6_ASAP7_75t_L g288 ( 
.A(n_169),
.B(n_266),
.Y(n_288)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_174),
.Y(n_409)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_176),
.Y(n_241)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_184),
.B(n_333),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_203),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_187),
.Y(n_444)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_190),
.Y(n_462)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_200),
.B2(n_201),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g448 ( 
.A1(n_191),
.A2(n_192),
.B(n_200),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_196),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_203),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_206),
.B(n_209),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_216),
.C(n_219),
.Y(n_209)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_210),
.B(n_220),
.Y(n_277)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_216),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_217),
.B(n_287),
.C(n_337),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_217),
.A2(n_343),
.B(n_345),
.C(n_369),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_217),
.B(n_377),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_242),
.B(n_244),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_221),
.Y(n_258)
);

NAND2x1p5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_222),
.B(n_265),
.Y(n_264)
);

XOR2x2_ASAP7_75t_SL g284 ( 
.A(n_222),
.B(n_224),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_222),
.A2(n_265),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_222),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_222),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_222),
.A2(n_287),
.B1(n_288),
.B2(n_319),
.Y(n_402)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_222),
.A2(n_319),
.B1(n_387),
.B2(n_388),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B1(n_239),
.B2(n_241),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_225),
.A2(n_232),
.B1(n_266),
.B2(n_271),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_228),
.Y(n_274)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx4f_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_244),
.B(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_242),
.A2(n_246),
.B(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AND3x1_ASAP7_75t_L g322 ( 
.A(n_246),
.B(n_323),
.C(n_324),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_426),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_339),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_313),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_278),
.Y(n_250)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_251),
.Y(n_428)
);

NAND2x1p5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_275),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g438 ( 
.A(n_252),
.B(n_275),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.C(n_262),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_259),
.Y(n_280)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_264),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_255),
.A2(n_257),
.B1(n_286),
.B2(n_317),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_265),
.Y(n_320)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_278),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_279),
.B(n_281),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_283),
.B(n_284),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_285),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_289),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_290),
.Y(n_334)
);

NAND2x1p5_ASAP7_75t_L g373 ( 
.A(n_287),
.B(n_346),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_287),
.A2(n_288),
.B1(n_337),
.B2(n_338),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_287),
.B(n_374),
.C(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_287),
.B(n_416),
.Y(n_415)
);

CKINVDCx11_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_288),
.B(n_346),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_288),
.B(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_288),
.B(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_298),
.B(n_303),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_296),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx4f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_307),
.B(n_312),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx2_ASAP7_75t_SL g308 ( 
.A(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_327),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_314),
.B(n_435),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_325),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_315),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_318),
.C(n_321),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_329),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_321),
.B1(n_322),
.B2(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_319),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_325),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_331),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g435 ( 
.A(n_328),
.B(n_331),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_334),
.C(n_335),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_332),
.B(n_424),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_345),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_336),
.Y(n_424)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21x1_ASAP7_75t_SL g339 ( 
.A1(n_340),
.A2(n_421),
.B(n_425),
.Y(n_339)
);

AOI21x1_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_379),
.B(n_420),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_370),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_344),
.A2(n_372),
.B1(n_373),
.B2(n_374),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_344),
.B(n_373),
.C(n_375),
.Y(n_422)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_350),
.B(n_358),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_363),
.B(n_367),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_366),
.Y(n_391)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_375),
.B1(n_376),
.B2(n_378),
.Y(n_370)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_371),
.Y(n_378)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI21x1_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_384),
.B(n_419),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_381),
.B(n_382),
.Y(n_419)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_383),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_404),
.B(n_417),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_400),
.Y(n_385)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_415),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2x1_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_422),
.B(n_423),
.Y(n_425)
);

AOI21x1_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_430),
.B(n_436),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_428),
.A2(n_437),
.B(n_438),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_463),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_446),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_442),
.B(n_446),
.Y(n_473)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_461),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_452),
.B1(n_454),
.B2(n_460),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

OA22x2_ASAP7_75t_SL g483 ( 
.A1(n_452),
.A2(n_454),
.B1(n_460),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_457),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_459),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_461),
.B(n_480),
.C(n_481),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_463),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_463),
.B(n_476),
.C(n_491),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_L g472 ( 
.A1(n_465),
.A2(n_473),
.B(n_474),
.C(n_475),
.Y(n_472)
);

AND3x1_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_476),
.C(n_491),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_471),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVxp33_ASAP7_75t_SL g476 ( 
.A(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_482),
.Y(n_477)
);

INVxp33_ASAP7_75t_SL g478 ( 
.A(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_479),
.B(n_483),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx4_ASAP7_75t_SL g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);


endmodule