module fake_jpeg_11124_n_202 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx6_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_10),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_31),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_19),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_73),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_90),
.Y(n_109)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_59),
.B(n_0),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_0),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_69),
.B1(n_75),
.B2(n_74),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_72),
.B1(n_61),
.B2(n_63),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_100),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_65),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_105),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_86),
.B1(n_75),
.B2(n_92),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_58),
.B1(n_68),
.B2(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_79),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_76),
.B(n_64),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_117),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_108),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_2),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_97),
.A2(n_84),
.B1(n_71),
.B2(n_80),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_131),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_97),
.A2(n_103),
.B1(n_84),
.B2(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_67),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_125),
.B1(n_126),
.B2(n_131),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_104),
.A2(n_71),
.B1(n_78),
.B2(n_82),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_125)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_63),
.C(n_81),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_148),
.C(n_149),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_2),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_138),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_3),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_4),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_143),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_4),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_5),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_145),
.B(n_153),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_81),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_12),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_81),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_33),
.C(n_55),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_126),
.A2(n_32),
.B1(n_52),
.B2(n_49),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_38),
.B1(n_46),
.B2(n_45),
.Y(n_158)
);

AO22x1_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_56),
.B1(n_28),
.B2(n_29),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_154),
.A2(n_165),
.B(n_16),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_137),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_147),
.B1(n_18),
.B2(n_17),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_140),
.B(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_158),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_47),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_140),
.C(n_147),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_161),
.B(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_139),
.B(n_13),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_164),
.B(n_166),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_14),
.B(n_15),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_14),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_15),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_165),
.B1(n_156),
.B2(n_158),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_175),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_176),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_177),
.A2(n_155),
.B1(n_170),
.B2(n_162),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_34),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_183),
.C(n_43),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_40),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_177),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_181),
.A2(n_154),
.B1(n_160),
.B2(n_17),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_189),
.B1(n_174),
.B2(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_193),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_173),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_178),
.B(n_188),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_187),
.B(n_179),
.C(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_199),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_44),
.Y(n_202)
);


endmodule