module fake_jpeg_25830_n_252 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_1),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_2),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_22),
.B1(n_21),
.B2(n_26),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_61),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_18),
.C(n_32),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_44),
.C(n_24),
.Y(n_98)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_32),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_32),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_22),
.B1(n_21),
.B2(n_26),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_17),
.B1(n_31),
.B2(n_23),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_34),
.B1(n_17),
.B2(n_25),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_73),
.Y(n_95)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_32),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_47),
.B1(n_44),
.B2(n_20),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_98),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_40),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_105),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_40),
.B(n_39),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_47),
.C(n_3),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_82),
.Y(n_120)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_37),
.B1(n_23),
.B2(n_25),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_83),
.A2(n_91),
.B1(n_103),
.B2(n_20),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_94),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_2),
.C(n_3),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_106),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_64),
.A2(n_28),
.B1(n_27),
.B2(n_30),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_72),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_29),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_99),
.Y(n_109)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_3),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_27),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_53),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_53),
.B(n_24),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_60),
.B1(n_70),
.B2(n_63),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_123),
.B1(n_128),
.B2(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_69),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_77),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_77),
.B1(n_87),
.B2(n_83),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_129),
.B1(n_89),
.B2(n_75),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_28),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_75),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_80),
.A2(n_70),
.B1(n_60),
.B2(n_57),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_132),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_52),
.B1(n_44),
.B2(n_28),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_93),
.Y(n_149)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_134),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_124),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_130),
.B(n_100),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_140),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_138),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_110),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_89),
.B1(n_96),
.B2(n_97),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_141),
.A2(n_151),
.B1(n_128),
.B2(n_107),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_146),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_116),
.B(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_127),
.A2(n_82),
.B(n_20),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_154),
.B(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_157),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_20),
.C(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_129),
.A2(n_93),
.B1(n_86),
.B2(n_85),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_117),
.B(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_156),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_115),
.A2(n_76),
.B(n_24),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_4),
.B(n_5),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_122),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_160),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_125),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_137),
.B1(n_144),
.B2(n_149),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_171),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_114),
.C(n_109),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_165),
.B(n_175),
.C(n_177),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_118),
.B1(n_112),
.B2(n_114),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_119),
.B1(n_113),
.B2(n_111),
.Y(n_191)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_178),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_148),
.A2(n_118),
.B(n_126),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_155),
.B(n_154),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_109),
.C(n_113),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_142),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_150),
.Y(n_182)
);

XOR2x1_ASAP7_75t_SL g213 ( 
.A(n_182),
.B(n_190),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_162),
.B1(n_163),
.B2(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_169),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_146),
.B1(n_142),
.B2(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_197),
.B1(n_166),
.B2(n_170),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_159),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_136),
.A3(n_119),
.B1(n_157),
.B2(n_156),
.C1(n_134),
.C2(n_30),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_193),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_176),
.B(n_164),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_135),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_140),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_195),
.B(n_198),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_200),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_107),
.B1(n_111),
.B2(n_8),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_6),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_167),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_210),
.B1(n_183),
.B2(n_185),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_187),
.C(n_165),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_187),
.C(n_177),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_160),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_166),
.Y(n_214)
);

AO21x1_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_203),
.B(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_212),
.C(n_202),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_193),
.B(n_182),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_221),
.B(n_224),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_199),
.B(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_191),
.C(n_167),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_6),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_213),
.B1(n_209),
.B2(n_9),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_198),
.B(n_197),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_174),
.B(n_7),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_174),
.B1(n_210),
.B2(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_226),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_233),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_232),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_6),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_7),
.C(n_9),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_230),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_235),
.B(n_216),
.Y(n_244)
);

AOI31xp33_ASAP7_75t_L g236 ( 
.A1(n_234),
.A2(n_219),
.A3(n_215),
.B(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_238),
.Y(n_241)
);

NAND4xp25_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_7),
.C(n_10),
.D(n_11),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_228),
.B(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_226),
.C(n_12),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_241),
.A2(n_239),
.B(n_235),
.C(n_238),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_245),
.A2(n_13),
.B(n_15),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_10),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_249),
.C(n_247),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_13),
.B(n_15),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_15),
.Y(n_252)
);


endmodule