module fake_netlist_1_9145_n_1170 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1170);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1170;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_1056;
wire n_802;
wire n_985;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1097;
wire n_324;
wire n_1125;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_1169;
wire n_652;
wire n_1042;
wire n_279;
wire n_303;
wire n_975;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_1132;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_844;
wire n_818;
wire n_1160;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1063;
wire n_767;
wire n_828;
wire n_1138;
wire n_293;
wire n_1014;
wire n_506;
wire n_533;
wire n_490;
wire n_393;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_1157;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1017;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_446;
wire n_285;
wire n_423;
wire n_420;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_806;
wire n_881;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_1159;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1069;
wire n_1021;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_912;
wire n_841;
wire n_947;
wire n_924;
wire n_1043;
wire n_378;
wire n_582;
wire n_1141;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_901;
wire n_834;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
wire n_1127;
INVx2_ASAP7_75t_L g272 ( .A(n_204), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_145), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_271), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_111), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_175), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_157), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g278 ( .A(n_134), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_0), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_190), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_267), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_23), .Y(n_282) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_109), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
INVxp33_ASAP7_75t_SL g285 ( .A(n_47), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_243), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_120), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_144), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_104), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_146), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_106), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_184), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_127), .Y(n_293) );
INVx1_ASAP7_75t_SL g294 ( .A(n_235), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_107), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_147), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_149), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_60), .Y(n_298) );
CKINVDCx5p33_ASAP7_75t_R g299 ( .A(n_71), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_211), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_143), .Y(n_301) );
BUFx2_ASAP7_75t_L g302 ( .A(n_165), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_78), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_131), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_229), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_178), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_132), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_135), .Y(n_309) );
BUFx10_ASAP7_75t_L g310 ( .A(n_17), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_96), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_194), .Y(n_312) );
XOR2xp5_ASAP7_75t_L g313 ( .A(n_268), .B(n_92), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_183), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_130), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_121), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_55), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_13), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_155), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_148), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g321 ( .A(n_85), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_193), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_266), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_93), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_32), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_8), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_159), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_138), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_65), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_97), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_13), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_84), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_0), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_93), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_166), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_12), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_168), .Y(n_337) );
BUFx5_ASAP7_75t_L g338 ( .A(n_215), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_79), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_205), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_63), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_66), .Y(n_342) );
INVxp67_ASAP7_75t_L g343 ( .A(n_3), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_117), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_61), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_209), .B(n_181), .Y(n_346) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_217), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_26), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_39), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_108), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_24), .B(n_82), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_244), .Y(n_352) );
BUFx2_ASAP7_75t_SL g353 ( .A(n_50), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_167), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_150), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_208), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_239), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_195), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_265), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_189), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_220), .Y(n_361) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_38), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_27), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_102), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_59), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_27), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_234), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_103), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_79), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_88), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_26), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_185), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_133), .Y(n_373) );
BUFx5_ASAP7_75t_L g374 ( .A(n_52), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_231), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_91), .Y(n_376) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_39), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_4), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_225), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_17), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_73), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_250), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_33), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_214), .Y(n_384) );
CKINVDCx16_ASAP7_75t_R g385 ( .A(n_164), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_67), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_76), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_76), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_52), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_264), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_42), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_170), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_24), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_105), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_113), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_22), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_56), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_212), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_95), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g400 ( .A(n_2), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_128), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_198), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_197), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_256), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_206), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_114), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_173), .Y(n_407) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_385), .B(n_270), .Y(n_408) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_308), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_374), .Y(n_410) );
OA21x2_ASAP7_75t_L g411 ( .A1(n_272), .A2(n_1), .B(n_2), .Y(n_411) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_308), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_374), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_338), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_374), .Y(n_415) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_371), .B(n_1), .Y(n_416) );
AND2x4_ASAP7_75t_L g417 ( .A(n_302), .B(n_3), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_363), .B(n_5), .Y(n_418) );
OA21x2_ASAP7_75t_L g419 ( .A1(n_272), .A2(n_5), .B(n_6), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_338), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_355), .B(n_6), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_324), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_308), .Y(n_424) );
INVxp67_ASAP7_75t_L g425 ( .A(n_360), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_338), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_372), .B(n_7), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_375), .B(n_9), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_338), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_389), .B(n_10), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_389), .B(n_10), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_374), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_283), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_338), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_338), .Y(n_435) );
OA21x2_ASAP7_75t_L g436 ( .A1(n_289), .A2(n_11), .B(n_14), .Y(n_436) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_308), .Y(n_437) );
OA21x2_ASAP7_75t_L g438 ( .A1(n_289), .A2(n_11), .B(n_14), .Y(n_438) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_337), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_374), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_374), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_337), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_371), .B(n_380), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_380), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_337), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_361), .B(n_15), .Y(n_446) );
OAI21x1_ASAP7_75t_L g447 ( .A1(n_361), .A2(n_99), .B(n_98), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_273), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_433), .B(n_365), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_422), .B(n_366), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_425), .B(n_297), .Y(n_452) );
INVx2_ASAP7_75t_SL g453 ( .A(n_417), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_422), .A2(n_388), .B1(n_400), .B2(n_321), .Y(n_455) );
INVx1_ASAP7_75t_SL g456 ( .A(n_418), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_410), .Y(n_457) );
BUFx3_ASAP7_75t_L g458 ( .A(n_443), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_418), .B(n_343), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g460 ( .A(n_408), .B(n_278), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_418), .B(n_310), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_448), .B(n_300), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_410), .Y(n_463) );
INVx8_ASAP7_75t_L g464 ( .A(n_417), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_448), .B(n_311), .Y(n_465) );
OR2x6_ASAP7_75t_L g466 ( .A(n_417), .B(n_353), .Y(n_466) );
INVx1_ASAP7_75t_SL g467 ( .A(n_427), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_443), .B(n_444), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_417), .B(n_281), .Y(n_469) );
NAND2xp33_ASAP7_75t_L g470 ( .A(n_427), .B(n_275), .Y(n_470) );
INVxp67_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_440), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_440), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_443), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_440), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_440), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_443), .B(n_356), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_443), .B(n_310), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_444), .B(n_394), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_413), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_421), .B(n_292), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_414), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_430), .B(n_351), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_428), .B(n_317), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_446), .Y(n_487) );
BUFx2_ASAP7_75t_L g488 ( .A(n_446), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_415), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_415), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_414), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_423), .Y(n_492) );
NAND2xp33_ASAP7_75t_L g493 ( .A(n_464), .B(n_346), .Y(n_493) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_460), .A2(n_408), .B1(n_305), .B2(n_354), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_SL g495 ( .A1(n_480), .A2(n_428), .B(n_432), .C(n_423), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_458), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_458), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_475), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_464), .Y(n_499) );
AND3x1_ASAP7_75t_L g500 ( .A(n_461), .B(n_416), .C(n_313), .Y(n_500) );
OR2x6_ASAP7_75t_L g501 ( .A(n_464), .B(n_430), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_475), .Y(n_502) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_467), .B(n_305), .Y(n_503) );
BUFx12f_ASAP7_75t_L g504 ( .A(n_466), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_479), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_487), .A2(n_431), .B1(n_430), .B2(n_411), .Y(n_506) );
NAND2xp33_ASAP7_75t_L g507 ( .A(n_453), .B(n_292), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_482), .B(n_430), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_453), .B(n_431), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_452), .B(n_431), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_461), .B(n_431), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_459), .B(n_293), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_455), .B(n_279), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_487), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_310), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_468), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_487), .A2(n_411), .B1(n_436), .B2(n_419), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_486), .B(n_282), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_462), .B(n_295), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_488), .A2(n_411), .B1(n_436), .B2(n_419), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_465), .B(n_295), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_466), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_484), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_459), .B(n_404), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_488), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_471), .B(n_404), .Y(n_526) );
AO22x1_ASAP7_75t_L g527 ( .A1(n_451), .A2(n_285), .B1(n_407), .B2(n_405), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_485), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_485), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_449), .B(n_405), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_485), .A2(n_411), .B1(n_436), .B2(n_419), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_485), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_485), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_478), .B(n_274), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_486), .B(n_432), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_469), .B(n_441), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_451), .B(n_441), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_466), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_466), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_472), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_491), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_470), .B(n_299), .Y(n_542) );
OR2x6_ASAP7_75t_L g543 ( .A(n_463), .B(n_447), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_450), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_450), .B(n_286), .Y(n_545) );
AND2x2_ASAP7_75t_SL g546 ( .A(n_454), .B(n_411), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_491), .A2(n_419), .B1(n_436), .B2(n_411), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_454), .B(n_287), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_481), .A2(n_419), .B1(n_438), .B2(n_436), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_457), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_481), .B(n_362), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_483), .B(n_307), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g553 ( .A1(n_489), .A2(n_303), .B(n_318), .C(n_298), .Y(n_553) );
NAND3xp33_ASAP7_75t_SL g554 ( .A(n_489), .B(n_378), .C(n_370), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_473), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_490), .B(n_492), .C(n_474), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_474), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_476), .B(n_276), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_490), .A2(n_354), .B1(n_403), .B2(n_315), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_477), .A2(n_403), .B1(n_315), .B2(n_383), .Y(n_560) );
INVxp67_ASAP7_75t_L g561 ( .A(n_477), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_453), .A2(n_447), .B(n_436), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_464), .Y(n_563) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_464), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_455), .B(n_381), .Y(n_565) );
NAND2xp33_ASAP7_75t_L g566 ( .A(n_464), .B(n_344), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_464), .B(n_350), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_482), .B(n_277), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_458), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_528), .B(n_358), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_562), .A2(n_447), .B(n_420), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_530), .B(n_345), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_505), .B(n_393), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_512), .B(n_349), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_496), .Y(n_576) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_562), .A2(n_420), .B(n_414), .Y(n_577) );
AND2x4_ASAP7_75t_L g578 ( .A(n_499), .B(n_325), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g579 ( .A1(n_528), .A2(n_438), .B1(n_419), .B2(n_369), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_499), .B(n_326), .Y(n_580) );
AO32x2_ASAP7_75t_L g581 ( .A1(n_543), .A2(n_438), .A3(n_409), .B1(n_437), .B2(n_424), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_524), .B(n_349), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_563), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_537), .B(n_396), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_508), .A2(n_509), .B(n_561), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_497), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_503), .A2(n_376), .B1(n_386), .B2(n_369), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_528), .A2(n_386), .B1(n_391), .B2(n_376), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_561), .A2(n_426), .B(n_420), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_553), .A2(n_331), .B(n_332), .C(n_329), .Y(n_590) );
A2O1A1Ixp33_ASAP7_75t_L g591 ( .A1(n_510), .A2(n_568), .B(n_534), .C(n_558), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_551), .B(n_438), .Y(n_592) );
INVx2_ASAP7_75t_SL g593 ( .A(n_504), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_546), .A2(n_434), .B(n_429), .Y(n_594) );
BUFx4f_ASAP7_75t_L g595 ( .A(n_501), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_498), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_563), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_493), .A2(n_438), .B1(n_391), .B2(n_434), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_519), .A2(n_334), .B(n_333), .Y(n_599) );
AOI21xp5_ASAP7_75t_L g600 ( .A1(n_546), .A2(n_434), .B(n_429), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_511), .B(n_336), .Y(n_602) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_564), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_543), .A2(n_435), .B(n_434), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_543), .A2(n_435), .B(n_280), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_544), .A2(n_435), .B(n_284), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_502), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_564), .B(n_339), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_515), .B(n_341), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_521), .B(n_342), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_557), .A2(n_291), .B(n_290), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_525), .B(n_348), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_522), .Y(n_613) );
BUFx8_ASAP7_75t_L g614 ( .A(n_513), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_559), .B(n_387), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_569), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_SL g617 ( .A1(n_495), .A2(n_301), .B(n_304), .C(n_296), .Y(n_617) );
OR2x6_ASAP7_75t_L g618 ( .A(n_501), .B(n_397), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_550), .Y(n_619) );
AOI21xp5_ASAP7_75t_L g620 ( .A1(n_536), .A2(n_309), .B(n_306), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_539), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_506), .A2(n_314), .B(n_312), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_556), .A2(n_319), .B(n_316), .Y(n_623) );
AOI33xp33_ASAP7_75t_L g624 ( .A1(n_553), .A2(n_399), .A3(n_359), .B1(n_320), .B2(n_322), .B3(n_323), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_542), .B(n_288), .Y(n_625) );
NOR2xp33_ASAP7_75t_SL g626 ( .A(n_494), .B(n_367), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_527), .B(n_568), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_516), .B(n_368), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_565), .A2(n_330), .B(n_335), .C(n_328), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_539), .B(n_384), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_526), .B(n_401), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_529), .B(n_294), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_532), .B(n_327), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_533), .B(n_340), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_494), .A2(n_377), .B1(n_352), .B2(n_357), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_555), .Y(n_636) );
INVx3_ASAP7_75t_L g637 ( .A(n_522), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_560), .B(n_15), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_538), .Y(n_639) );
INVx2_ASAP7_75t_SL g640 ( .A(n_552), .Y(n_640) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_531), .A2(n_395), .B1(n_398), .B2(n_392), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_500), .B(n_16), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_540), .B(n_364), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_523), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_531), .A2(n_382), .B(n_390), .C(n_373), .Y(n_645) );
INVxp33_ASAP7_75t_SL g646 ( .A(n_567), .Y(n_646) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_545), .B(n_382), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_520), .A2(n_402), .B1(n_406), .B2(n_390), .Y(n_648) );
INVx3_ASAP7_75t_L g649 ( .A(n_541), .Y(n_649) );
INVxp33_ASAP7_75t_SL g650 ( .A(n_548), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_554), .A2(n_347), .B1(n_379), .B2(n_337), .Y(n_651) );
NAND2xp33_ASAP7_75t_L g652 ( .A(n_517), .B(n_347), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_507), .B(n_18), .Y(n_653) );
AO22x1_ASAP7_75t_L g654 ( .A1(n_566), .A2(n_379), .B1(n_549), .B2(n_547), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g655 ( .A(n_547), .B(n_445), .Y(n_655) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_562), .A2(n_412), .B(n_409), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_562), .A2(n_412), .B(n_409), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_562), .A2(n_412), .B(n_409), .Y(n_658) );
INVx4_ASAP7_75t_L g659 ( .A(n_499), .Y(n_659) );
NOR2xp33_ASAP7_75t_SL g660 ( .A(n_494), .B(n_412), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_505), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_514), .Y(n_662) );
INVx2_ASAP7_75t_SL g663 ( .A(n_504), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_493), .A2(n_437), .B1(n_439), .B2(n_424), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_514), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_518), .B(n_19), .Y(n_666) );
AO21x1_ASAP7_75t_L g667 ( .A1(n_562), .A2(n_437), .B(n_424), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_535), .B(n_19), .Y(n_668) );
AOI21x1_ASAP7_75t_L g669 ( .A1(n_562), .A2(n_437), .B(n_424), .Y(n_669) );
AOI21x1_ASAP7_75t_L g670 ( .A1(n_562), .A2(n_437), .B(n_424), .Y(n_670) );
OAI21xp5_ASAP7_75t_L g671 ( .A1(n_562), .A2(n_442), .B(n_439), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_535), .B(n_20), .Y(n_672) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_528), .A2(n_442), .B1(n_445), .B2(n_439), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_535), .B(n_20), .Y(n_674) );
BUFx6f_ASAP7_75t_L g675 ( .A(n_563), .Y(n_675) );
INVx2_ASAP7_75t_L g676 ( .A(n_514), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_499), .Y(n_677) );
BUFx2_ASAP7_75t_R g678 ( .A(n_627), .Y(n_678) );
INVx3_ASAP7_75t_L g679 ( .A(n_659), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_661), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g681 ( .A1(n_645), .A2(n_442), .B(n_439), .Y(n_681) );
BUFx8_ASAP7_75t_L g682 ( .A(n_593), .Y(n_682) );
NOR2xp33_ASAP7_75t_SL g683 ( .A(n_595), .B(n_21), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_585), .A2(n_445), .B(n_100), .Y(n_684) );
AOI221x1_ASAP7_75t_L g685 ( .A1(n_656), .A2(n_445), .B1(n_28), .B2(n_29), .C(n_30), .Y(n_685) );
OAI21x1_ASAP7_75t_L g686 ( .A1(n_669), .A2(n_445), .B(n_101), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_588), .B(n_25), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_650), .B(n_615), .Y(n_688) );
BUFx10_ASAP7_75t_L g689 ( .A(n_618), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_609), .B(n_30), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_629), .A2(n_445), .B1(n_32), .B2(n_33), .C(n_34), .Y(n_691) );
OAI21x1_ASAP7_75t_L g692 ( .A1(n_657), .A2(n_112), .B(n_110), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_594), .A2(n_116), .B(n_115), .Y(n_693) );
AO32x2_ASAP7_75t_L g694 ( .A1(n_648), .A2(n_31), .A3(n_34), .B1(n_35), .B2(n_36), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_618), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_618), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_592), .A2(n_119), .B(n_118), .Y(n_697) );
NOR2xp67_ASAP7_75t_L g698 ( .A(n_663), .B(n_37), .Y(n_698) );
OAI21x1_ASAP7_75t_L g699 ( .A1(n_658), .A2(n_123), .B(n_122), .Y(n_699) );
BUFx3_ASAP7_75t_L g700 ( .A(n_614), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_598), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_701) );
AO22x2_ASAP7_75t_L g702 ( .A1(n_635), .A2(n_40), .B1(n_41), .B2(n_43), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_600), .A2(n_125), .B(n_124), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_622), .A2(n_44), .B(n_45), .C(n_46), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_614), .Y(n_705) );
OAI21xp5_ASAP7_75t_L g706 ( .A1(n_605), .A2(n_129), .B(n_126), .Y(n_706) );
INVx3_ASAP7_75t_L g707 ( .A(n_659), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_608), .Y(n_708) );
OAI21x1_ASAP7_75t_L g709 ( .A1(n_571), .A2(n_137), .B(n_136), .Y(n_709) );
OAI21x1_ASAP7_75t_L g710 ( .A1(n_577), .A2(n_140), .B(n_139), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_598), .A2(n_44), .B(n_45), .C(n_46), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g712 ( .A1(n_604), .A2(n_142), .B(n_141), .Y(n_712) );
BUFx3_ASAP7_75t_L g713 ( .A(n_601), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_575), .B(n_47), .Y(n_714) );
AO31x2_ASAP7_75t_L g715 ( .A1(n_641), .A2(n_48), .A3(n_49), .B(n_50), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g716 ( .A1(n_666), .A2(n_48), .B(n_49), .C(n_51), .Y(n_716) );
INVx4_ASAP7_75t_L g717 ( .A(n_595), .Y(n_717) );
INVx3_ASAP7_75t_SL g718 ( .A(n_578), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_624), .B(n_53), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_601), .B(n_53), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_677), .B(n_54), .Y(n_721) );
BUFx3_ASAP7_75t_L g722 ( .A(n_603), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_587), .A2(n_54), .B1(n_55), .B2(n_56), .C(n_57), .Y(n_723) );
NOR4xp25_ASAP7_75t_L g724 ( .A(n_590), .B(n_57), .C(n_58), .D(n_59), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_589), .A2(n_152), .B(n_151), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_608), .Y(n_726) );
BUFx10_ASAP7_75t_L g727 ( .A(n_578), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_639), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g729 ( .A1(n_579), .A2(n_154), .B(n_153), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_582), .B(n_62), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_573), .B(n_63), .Y(n_731) );
OR2x2_ASAP7_75t_L g732 ( .A(n_638), .B(n_64), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_668), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_733) );
BUFx2_ASAP7_75t_L g734 ( .A(n_621), .Y(n_734) );
BUFx10_ASAP7_75t_L g735 ( .A(n_580), .Y(n_735) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_603), .Y(n_736) );
AO31x2_ASAP7_75t_L g737 ( .A1(n_672), .A2(n_68), .A3(n_69), .B(n_70), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_606), .A2(n_201), .B(n_263), .Y(n_738) );
OAI21xp5_ASAP7_75t_L g739 ( .A1(n_611), .A2(n_200), .B(n_262), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_646), .Y(n_740) );
AOI21xp5_ASAP7_75t_SL g741 ( .A1(n_664), .A2(n_269), .B(n_199), .Y(n_741) );
OAI21x1_ASAP7_75t_L g742 ( .A1(n_664), .A2(n_196), .B(n_260), .Y(n_742) );
NAND2xp33_ASAP7_75t_L g743 ( .A(n_603), .B(n_156), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_643), .A2(n_202), .B(n_259), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_642), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_576), .Y(n_746) );
BUFx3_ASAP7_75t_L g747 ( .A(n_675), .Y(n_747) );
AO31x2_ASAP7_75t_L g748 ( .A1(n_674), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_748) );
OAI21x1_ASAP7_75t_L g749 ( .A1(n_673), .A2(n_203), .B(n_258), .Y(n_749) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_675), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_586), .Y(n_751) );
AO31x2_ASAP7_75t_L g752 ( .A1(n_623), .A2(n_74), .A3(n_75), .B(n_77), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_647), .A2(n_631), .B(n_628), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_572), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g755 ( .A1(n_610), .A2(n_191), .B(n_255), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_649), .A2(n_188), .B(n_254), .Y(n_756) );
OR2x6_ASAP7_75t_L g757 ( .A(n_640), .B(n_77), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g758 ( .A1(n_620), .A2(n_192), .B(n_253), .Y(n_758) );
OA21x2_ASAP7_75t_L g759 ( .A1(n_651), .A2(n_187), .B(n_252), .Y(n_759) );
OAI21x1_ASAP7_75t_L g760 ( .A1(n_649), .A2(n_186), .B(n_251), .Y(n_760) );
AO31x2_ASAP7_75t_L g761 ( .A1(n_653), .A2(n_78), .A3(n_80), .B(n_81), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_596), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_619), .Y(n_763) );
OAI21x1_ASAP7_75t_L g764 ( .A1(n_636), .A2(n_207), .B(n_249), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_675), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_617), .A2(n_182), .B(n_248), .Y(n_766) );
CKINVDCx6p67_ASAP7_75t_R g767 ( .A(n_570), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_644), .A2(n_180), .B(n_247), .Y(n_768) );
INVx2_ASAP7_75t_L g769 ( .A(n_662), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_602), .A2(n_179), .B(n_246), .Y(n_770) );
AND2x2_ASAP7_75t_L g771 ( .A(n_584), .B(n_80), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_625), .B(n_83), .Y(n_772) );
OAI21x1_ASAP7_75t_L g773 ( .A1(n_665), .A2(n_213), .B(n_245), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_L g774 ( .A1(n_599), .A2(n_84), .B(n_85), .C(n_86), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_676), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_612), .B(n_86), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g777 ( .A1(n_574), .A2(n_216), .B(n_242), .Y(n_777) );
OAI21x1_ASAP7_75t_L g778 ( .A1(n_613), .A2(n_177), .B(n_241), .Y(n_778) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_660), .B(n_87), .C(n_88), .Y(n_779) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_677), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_633), .B(n_89), .Y(n_781) );
AOI21xp5_ASAP7_75t_L g782 ( .A1(n_632), .A2(n_218), .B(n_240), .Y(n_782) );
AO31x2_ASAP7_75t_L g783 ( .A1(n_581), .A2(n_89), .A3(n_90), .B(n_91), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_607), .Y(n_784) );
BUFx8_ASAP7_75t_L g785 ( .A(n_581), .Y(n_785) );
A2O1A1Ixp33_ASAP7_75t_L g786 ( .A1(n_634), .A2(n_92), .B(n_94), .C(n_95), .Y(n_786) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_583), .Y(n_787) );
A2O1A1Ixp33_ASAP7_75t_L g788 ( .A1(n_616), .A2(n_94), .B(n_158), .C(n_160), .Y(n_788) );
OAI22x1_ASAP7_75t_L g789 ( .A1(n_630), .A2(n_161), .B1(n_162), .B2(n_163), .Y(n_789) );
BUFx3_ASAP7_75t_L g790 ( .A(n_583), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_637), .Y(n_791) );
AO31x2_ASAP7_75t_L g792 ( .A1(n_581), .A2(n_169), .A3(n_171), .B(n_172), .Y(n_792) );
AND2x4_ASAP7_75t_L g793 ( .A(n_637), .B(n_174), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_597), .Y(n_794) );
AOI221x1_ASAP7_75t_L g795 ( .A1(n_655), .A2(n_176), .B1(n_219), .B2(n_221), .C(n_222), .Y(n_795) );
NOR2xp67_ASAP7_75t_SL g796 ( .A(n_659), .B(n_223), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_619), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_652), .A2(n_224), .B(n_226), .Y(n_798) );
AO31x2_ASAP7_75t_L g799 ( .A1(n_667), .A2(n_227), .A3(n_228), .B(n_230), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_652), .A2(n_232), .B(n_233), .Y(n_800) );
OAI21xp33_ASAP7_75t_L g801 ( .A1(n_626), .A2(n_236), .B(n_237), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_591), .B(n_238), .Y(n_802) );
AOI21x1_ASAP7_75t_L g803 ( .A1(n_654), .A2(n_261), .B(n_670), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_619), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_652), .A2(n_655), .B(n_671), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_591), .B(n_467), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_688), .B(n_696), .Y(n_807) );
AO21x2_ASAP7_75t_L g808 ( .A1(n_803), .A2(n_681), .B(n_684), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_717), .B(n_695), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_682), .Y(n_810) );
OAI21xp5_ASAP7_75t_L g811 ( .A1(n_802), .A2(n_711), .B(n_753), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_797), .Y(n_812) );
INVxp67_ASAP7_75t_SL g813 ( .A(n_785), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_721), .Y(n_814) );
OA21x2_ASAP7_75t_L g815 ( .A1(n_795), .A2(n_686), .B(n_685), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_680), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_705), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_746), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_727), .B(n_735), .Y(n_819) );
OAI21x1_ASAP7_75t_L g820 ( .A1(n_710), .A2(n_709), .B(n_773), .Y(n_820) );
AO21x2_ASAP7_75t_L g821 ( .A1(n_729), .A2(n_766), .B(n_703), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_804), .B(n_751), .Y(n_822) );
OA21x2_ASAP7_75t_L g823 ( .A1(n_692), .A2(n_699), .B(n_693), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_804), .B(n_762), .Y(n_824) );
AND2x2_ASAP7_75t_SL g825 ( .A(n_683), .B(n_721), .Y(n_825) );
O2A1O1Ixp33_ASAP7_75t_L g826 ( .A1(n_786), .A2(n_716), .B(n_701), .C(n_719), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_763), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_728), .B(n_784), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_734), .B(n_732), .Y(n_829) );
OR2x2_ASAP7_75t_L g830 ( .A(n_687), .B(n_740), .Y(n_830) );
NAND2x1p5_ASAP7_75t_L g831 ( .A(n_679), .B(n_707), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_754), .Y(n_832) );
OA21x2_ASAP7_75t_L g833 ( .A1(n_742), .A2(n_764), .B(n_712), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_771), .B(n_769), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_702), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_775), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_756), .A2(n_760), .B(n_778), .Y(n_837) );
INVx3_ASAP7_75t_L g838 ( .A(n_679), .Y(n_838) );
BUFx2_ASAP7_75t_L g839 ( .A(n_780), .Y(n_839) );
OA21x2_ASAP7_75t_L g840 ( .A1(n_706), .A2(n_800), .B(n_798), .Y(n_840) );
INVx2_ASAP7_75t_SL g841 ( .A(n_689), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_776), .B(n_690), .Y(n_842) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_745), .B(n_735), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_702), .Y(n_844) );
INVx3_ASAP7_75t_L g845 ( .A(n_707), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_730), .B(n_700), .Y(n_846) );
INVx1_ASAP7_75t_L g847 ( .A(n_708), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_714), .B(n_726), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_737), .Y(n_849) );
OR2x2_ASAP7_75t_L g850 ( .A(n_772), .B(n_767), .Y(n_850) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_704), .A2(n_697), .B(n_782), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_781), .B(n_791), .Y(n_852) );
BUFx2_ASAP7_75t_R g853 ( .A(n_713), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_724), .B(n_691), .Y(n_854) );
OR2x6_ASAP7_75t_L g855 ( .A(n_793), .B(n_698), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_737), .Y(n_856) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_750), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_748), .Y(n_858) );
OAI21xp5_ASAP7_75t_L g859 ( .A1(n_777), .A2(n_755), .B(n_758), .Y(n_859) );
NAND2x1p5_ASAP7_75t_L g860 ( .A(n_722), .B(n_747), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_748), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_748), .Y(n_862) );
AO31x2_ASAP7_75t_L g863 ( .A1(n_789), .A2(n_774), .A3(n_788), .B(n_733), .Y(n_863) );
AO21x2_ASAP7_75t_L g864 ( .A1(n_738), .A2(n_739), .B(n_779), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_689), .B(n_794), .Y(n_865) );
OA21x2_ASAP7_75t_L g866 ( .A1(n_801), .A2(n_749), .B(n_770), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_715), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_723), .B(n_765), .Y(n_868) );
OA21x2_ASAP7_75t_L g869 ( .A1(n_725), .A2(n_768), .B(n_744), .Y(n_869) );
NAND2x1p5_ASAP7_75t_L g870 ( .A(n_790), .B(n_796), .Y(n_870) );
BUFx10_ASAP7_75t_L g871 ( .A(n_787), .Y(n_871) );
NAND2x1p5_ASAP7_75t_L g872 ( .A(n_787), .B(n_720), .Y(n_872) );
BUFx2_ASAP7_75t_L g873 ( .A(n_736), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_678), .B(n_694), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_715), .B(n_752), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_715), .B(n_752), .Y(n_876) );
INVx2_ASAP7_75t_L g877 ( .A(n_783), .Y(n_877) );
OA21x2_ASAP7_75t_L g878 ( .A1(n_792), .A2(n_799), .B(n_759), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_761), .Y(n_879) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_761), .Y(n_880) );
INVx2_ASAP7_75t_L g881 ( .A(n_752), .Y(n_881) );
OA21x2_ASAP7_75t_L g882 ( .A1(n_792), .A2(n_799), .B(n_761), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_799), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_741), .B(n_743), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_680), .Y(n_885) );
NAND2x1p5_ASAP7_75t_L g886 ( .A(n_717), .B(n_595), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_806), .B(n_591), .Y(n_887) );
AND2x4_ASAP7_75t_L g888 ( .A(n_717), .B(n_659), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_680), .Y(n_889) );
BUFx12f_ASAP7_75t_L g890 ( .A(n_682), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_680), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_806), .B(n_591), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_688), .B(n_467), .Y(n_893) );
INVx2_ASAP7_75t_SL g894 ( .A(n_682), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_680), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_806), .B(n_591), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_680), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_680), .Y(n_898) );
INVx2_ASAP7_75t_L g899 ( .A(n_797), .Y(n_899) );
CKINVDCx11_ASAP7_75t_R g900 ( .A(n_705), .Y(n_900) );
INVx1_ASAP7_75t_SL g901 ( .A(n_718), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_680), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_806), .B(n_591), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_680), .Y(n_904) );
AND2x2_ASAP7_75t_L g905 ( .A(n_688), .B(n_467), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_797), .Y(n_906) );
OR2x2_ASAP7_75t_L g907 ( .A(n_688), .B(n_588), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_680), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_685), .A2(n_667), .A3(n_645), .B(n_805), .Y(n_909) );
BUFx6f_ASAP7_75t_L g910 ( .A(n_750), .Y(n_910) );
BUFx4f_ASAP7_75t_L g911 ( .A(n_757), .Y(n_911) );
CKINVDCx11_ASAP7_75t_R g912 ( .A(n_705), .Y(n_912) );
A2O1A1Ixp33_ASAP7_75t_L g913 ( .A1(n_753), .A2(n_591), .B(n_806), .C(n_731), .Y(n_913) );
INVx2_ASAP7_75t_L g914 ( .A(n_797), .Y(n_914) );
NAND2x1p5_ASAP7_75t_L g915 ( .A(n_717), .B(n_595), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_835), .B(n_844), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_812), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_899), .B(n_906), .Y(n_918) );
AND2x4_ASAP7_75t_L g919 ( .A(n_914), .B(n_813), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_907), .B(n_830), .Y(n_920) );
INVx2_ASAP7_75t_SL g921 ( .A(n_888), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_828), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_832), .B(n_836), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_816), .Y(n_924) );
INVxp67_ASAP7_75t_SL g925 ( .A(n_814), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_893), .B(n_905), .Y(n_926) );
BUFx2_ASAP7_75t_L g927 ( .A(n_813), .Y(n_927) );
BUFx2_ASAP7_75t_L g928 ( .A(n_857), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_822), .B(n_824), .Y(n_929) );
OA21x2_ASAP7_75t_L g930 ( .A1(n_883), .A2(n_876), .B(n_875), .Y(n_930) );
AO21x1_ASAP7_75t_SL g931 ( .A1(n_875), .A2(n_876), .B(n_880), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_867), .Y(n_932) );
BUFx2_ASAP7_75t_L g933 ( .A(n_825), .Y(n_933) );
OR2x2_ASAP7_75t_L g934 ( .A(n_829), .B(n_887), .Y(n_934) );
INVxp33_ASAP7_75t_L g935 ( .A(n_819), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_807), .B(n_818), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_887), .B(n_892), .Y(n_937) );
AND2x2_ASAP7_75t_L g938 ( .A(n_885), .B(n_889), .Y(n_938) );
INVx2_ASAP7_75t_SL g939 ( .A(n_911), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_891), .Y(n_940) );
AO21x2_ASAP7_75t_L g941 ( .A1(n_849), .A2(n_862), .B(n_856), .Y(n_941) );
OR2x6_ASAP7_75t_L g942 ( .A(n_855), .B(n_870), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_895), .B(n_897), .Y(n_943) );
OR2x6_ASAP7_75t_L g944 ( .A(n_855), .B(n_870), .Y(n_944) );
INVx1_ASAP7_75t_L g945 ( .A(n_881), .Y(n_945) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_890), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_898), .B(n_902), .Y(n_947) );
BUFx3_ASAP7_75t_L g948 ( .A(n_810), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_904), .B(n_908), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g950 ( .A(n_846), .B(n_850), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g951 ( .A1(n_826), .A2(n_842), .B1(n_854), .B2(n_848), .C(n_892), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_877), .Y(n_952) );
OA21x2_ASAP7_75t_L g953 ( .A1(n_858), .A2(n_861), .B(n_879), .Y(n_953) );
AND2x2_ASAP7_75t_L g954 ( .A(n_827), .B(n_896), .Y(n_954) );
INVx5_ASAP7_75t_L g955 ( .A(n_910), .Y(n_955) );
HB1xp67_ASAP7_75t_L g956 ( .A(n_901), .Y(n_956) );
INVx2_ASAP7_75t_SL g957 ( .A(n_886), .Y(n_957) );
INVx2_ASAP7_75t_L g958 ( .A(n_882), .Y(n_958) );
AND2x2_ASAP7_75t_L g959 ( .A(n_896), .B(n_903), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_847), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_903), .B(n_834), .Y(n_961) );
INVx2_ASAP7_75t_L g962 ( .A(n_909), .Y(n_962) );
OR2x2_ASAP7_75t_L g963 ( .A(n_848), .B(n_834), .Y(n_963) );
BUFx2_ASAP7_75t_L g964 ( .A(n_873), .Y(n_964) );
BUFx4f_ASAP7_75t_L g965 ( .A(n_915), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_913), .B(n_874), .Y(n_966) );
BUFx6f_ASAP7_75t_L g967 ( .A(n_871), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_865), .Y(n_968) );
NOR2x1_ASAP7_75t_R g969 ( .A(n_900), .B(n_912), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_842), .B(n_838), .Y(n_970) );
AOI22xp5_ASAP7_75t_SL g971 ( .A1(n_894), .A2(n_817), .B1(n_843), .B2(n_839), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_865), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_909), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_852), .Y(n_974) );
INVx3_ASAP7_75t_L g975 ( .A(n_915), .Y(n_975) );
AO21x2_ASAP7_75t_L g976 ( .A1(n_811), .A2(n_808), .B(n_859), .Y(n_976) );
AND2x4_ASAP7_75t_L g977 ( .A(n_838), .B(n_845), .Y(n_977) );
INVx8_ASAP7_75t_L g978 ( .A(n_809), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_845), .B(n_831), .Y(n_979) );
INVx4_ASAP7_75t_L g980 ( .A(n_942), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_966), .B(n_878), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_932), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_959), .B(n_863), .Y(n_983) );
BUFx2_ASAP7_75t_L g984 ( .A(n_964), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_922), .B(n_868), .Y(n_985) );
AND2x4_ASAP7_75t_L g986 ( .A(n_932), .B(n_884), .Y(n_986) );
HB1xp67_ASAP7_75t_L g987 ( .A(n_964), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_916), .Y(n_988) );
HB1xp67_ASAP7_75t_L g989 ( .A(n_927), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_953), .Y(n_990) );
NOR2xp33_ASAP7_75t_L g991 ( .A(n_926), .B(n_841), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_959), .B(n_815), .Y(n_992) );
AND2x4_ASAP7_75t_L g993 ( .A(n_942), .B(n_837), .Y(n_993) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_927), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_953), .Y(n_995) );
AND2x4_ASAP7_75t_L g996 ( .A(n_942), .B(n_820), .Y(n_996) );
AND2x2_ASAP7_75t_L g997 ( .A(n_954), .B(n_815), .Y(n_997) );
BUFx2_ASAP7_75t_L g998 ( .A(n_928), .Y(n_998) );
BUFx3_ASAP7_75t_L g999 ( .A(n_965), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_945), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_935), .B(n_853), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_961), .B(n_864), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_938), .B(n_860), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1004 ( .A(n_919), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_919), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_938), .Y(n_1006) );
INVx5_ASAP7_75t_L g1007 ( .A(n_942), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_945), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_941), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_934), .B(n_860), .Y(n_1010) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_978), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_941), .Y(n_1012) );
AND2x4_ASAP7_75t_L g1013 ( .A(n_944), .B(n_851), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_943), .B(n_872), .Y(n_1014) );
BUFx3_ASAP7_75t_L g1015 ( .A(n_965), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_961), .B(n_833), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_943), .B(n_872), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1018 ( .A1(n_920), .A2(n_821), .B1(n_833), .B2(n_869), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_947), .B(n_823), .Y(n_1019) );
OR2x6_ASAP7_75t_L g1020 ( .A(n_944), .B(n_823), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_934), .B(n_866), .Y(n_1021) );
AND2x2_ASAP7_75t_L g1022 ( .A(n_947), .B(n_866), .Y(n_1022) );
INVx2_ASAP7_75t_L g1023 ( .A(n_958), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_929), .B(n_840), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_974), .B(n_963), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_918), .B(n_917), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_974), .B(n_963), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_970), .B(n_923), .Y(n_1028) );
NOR2xp33_ASAP7_75t_L g1029 ( .A(n_935), .B(n_950), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_924), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_936), .B(n_951), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1030), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_1006), .B(n_940), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_982), .Y(n_1034) );
AND2x6_ASAP7_75t_SL g1035 ( .A(n_1001), .B(n_969), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_982), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_983), .B(n_931), .Y(n_1037) );
NAND2xp33_ASAP7_75t_L g1038 ( .A(n_1007), .B(n_978), .Y(n_1038) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1023), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g1040 ( .A(n_991), .B(n_948), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_981), .B(n_931), .Y(n_1041) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_988), .B(n_930), .Y(n_1042) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_984), .B(n_930), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1028), .Y(n_1044) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_981), .B(n_930), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1000), .Y(n_1046) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1002), .B(n_952), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_984), .B(n_937), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1000), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1008), .Y(n_1050) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1008), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_999), .Y(n_1052) );
NAND2xp5_ASAP7_75t_SL g1053 ( .A(n_1007), .B(n_933), .Y(n_1053) );
INVx1_ASAP7_75t_L g1054 ( .A(n_987), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_989), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_990), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_994), .Y(n_1057) );
INVx3_ASAP7_75t_L g1058 ( .A(n_993), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1026), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1025), .B(n_960), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1016), .B(n_962), .Y(n_1061) );
OR2x2_ASAP7_75t_L g1062 ( .A(n_998), .B(n_937), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1026), .Y(n_1063) );
INVxp67_ASAP7_75t_L g1064 ( .A(n_1029), .Y(n_1064) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_996), .B(n_962), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1027), .B(n_972), .Y(n_1066) );
AND2x2_ASAP7_75t_L g1067 ( .A(n_1016), .B(n_973), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_995), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_992), .B(n_976), .Y(n_1069) );
AND2x2_ASAP7_75t_L g1070 ( .A(n_997), .B(n_976), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1056), .Y(n_1071) );
AND2x6_ASAP7_75t_SL g1072 ( .A(n_1040), .B(n_944), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1045), .B(n_1022), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1056), .Y(n_1074) );
NOR2xp33_ASAP7_75t_L g1075 ( .A(n_1064), .B(n_971), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_1058), .B(n_996), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1068), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1044), .B(n_1031), .Y(n_1078) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1068), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1034), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1034), .Y(n_1081) );
INVxp67_ASAP7_75t_L g1082 ( .A(n_1054), .Y(n_1082) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1036), .Y(n_1083) );
OR2x2_ASAP7_75t_L g1084 ( .A(n_1048), .B(n_1024), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1069), .B(n_986), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1036), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1087 ( .A(n_1052), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1088 ( .A(n_1070), .B(n_986), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1046), .Y(n_1089) );
NOR2xp67_ASAP7_75t_L g1090 ( .A(n_1058), .B(n_1007), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1070), .B(n_986), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1046), .Y(n_1092) );
INVx1_ASAP7_75t_SL g1093 ( .A(n_1041), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_1048), .B(n_1019), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1062), .B(n_1021), .Y(n_1095) );
INVx3_ASAP7_75t_L g1096 ( .A(n_1058), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1039), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1098 ( .A(n_1061), .B(n_1009), .Y(n_1098) );
HB1xp67_ASAP7_75t_L g1099 ( .A(n_1057), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1067), .B(n_1012), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1067), .B(n_1012), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1049), .Y(n_1102) );
INVxp67_ASAP7_75t_L g1103 ( .A(n_1075), .Y(n_1103) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_1093), .B(n_1059), .Y(n_1104) );
AND2x4_ASAP7_75t_L g1105 ( .A(n_1076), .B(n_1041), .Y(n_1105) );
AND2x4_ASAP7_75t_L g1106 ( .A(n_1076), .B(n_1037), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1107 ( .A(n_1078), .B(n_1055), .Y(n_1107) );
OR2x2_ASAP7_75t_L g1108 ( .A(n_1095), .B(n_1063), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_1076), .B(n_1037), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1080), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1081), .Y(n_1111) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1081), .Y(n_1112) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1084), .B(n_1032), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1084), .B(n_1042), .Y(n_1114) );
O2A1O1Ixp33_ASAP7_75t_SL g1115 ( .A1(n_1087), .A2(n_939), .B(n_1053), .C(n_1011), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1083), .Y(n_1116) );
NOR2xp33_ASAP7_75t_L g1117 ( .A(n_1099), .B(n_1035), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_1073), .B(n_1047), .Y(n_1118) );
NOR2xp33_ASAP7_75t_L g1119 ( .A(n_1082), .B(n_956), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1083), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1097), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1086), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1086), .Y(n_1123) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1097), .Y(n_1124) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1089), .Y(n_1125) );
AOI22xp5_ASAP7_75t_L g1126 ( .A1(n_1117), .A2(n_1091), .B1(n_1085), .B2(n_1088), .Y(n_1126) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_1114), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1113), .Y(n_1128) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_1103), .A2(n_1091), .B1(n_1085), .B2(n_1088), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1121), .Y(n_1130) );
HB1xp67_ASAP7_75t_SL g1131 ( .A(n_1106), .Y(n_1131) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_1114), .B(n_1098), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1107), .B(n_1072), .Y(n_1133) );
AOI222xp33_ASAP7_75t_L g1134 ( .A1(n_1119), .A2(n_1060), .B1(n_1033), .B2(n_1101), .C1(n_1100), .C2(n_1066), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_1118), .B(n_1073), .Y(n_1135) );
OAI21xp5_ASAP7_75t_L g1136 ( .A1(n_1115), .A2(n_1038), .B(n_1090), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g1137 ( .A1(n_1105), .A2(n_980), .B1(n_1076), .B2(n_1096), .Y(n_1137) );
OAI31xp33_ASAP7_75t_L g1138 ( .A1(n_1106), .A2(n_1096), .A3(n_1015), .B(n_1013), .Y(n_1138) );
AOI21xp5_ASAP7_75t_L g1139 ( .A1(n_1109), .A2(n_1090), .B(n_1096), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1127), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_1131), .A2(n_1109), .B1(n_1104), .B2(n_1108), .Y(n_1141) );
OAI322xp33_ASAP7_75t_SL g1142 ( .A1(n_1132), .A2(n_946), .A3(n_985), .B1(n_1123), .B2(n_1122), .C1(n_1120), .C2(n_1116), .Y(n_1142) );
AOI21xp5_ASAP7_75t_L g1143 ( .A1(n_1136), .A2(n_1094), .B(n_1110), .Y(n_1143) );
AOI221xp5_ASAP7_75t_L g1144 ( .A1(n_1133), .A2(n_1125), .B1(n_1112), .B2(n_1111), .C(n_1092), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1135), .B(n_1096), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1134), .B(n_1071), .Y(n_1146) );
AOI21xp33_ASAP7_75t_SL g1147 ( .A1(n_1138), .A2(n_978), .B(n_1043), .Y(n_1147) );
NOR2xp33_ASAP7_75t_L g1148 ( .A(n_1126), .B(n_1071), .Y(n_1148) );
AOI21xp5_ASAP7_75t_L g1149 ( .A1(n_1139), .A2(n_965), .B(n_1124), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1150 ( .A1(n_1137), .A2(n_980), .B1(n_1005), .B2(n_1004), .Y(n_1150) );
AOI221xp5_ASAP7_75t_SL g1151 ( .A1(n_1128), .A2(n_1003), .B1(n_1079), .B2(n_1077), .C(n_1074), .Y(n_1151) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_1129), .A2(n_1013), .B1(n_1065), .B2(n_996), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1153 ( .A1(n_1130), .A2(n_1102), .B1(n_1092), .B2(n_1050), .C(n_1051), .Y(n_1153) );
NOR3xp33_ASAP7_75t_L g1154 ( .A(n_1144), .B(n_1147), .C(n_1141), .Y(n_1154) );
AOI221x1_ASAP7_75t_L g1155 ( .A1(n_1146), .A2(n_1143), .B1(n_1140), .B2(n_1149), .C(n_1150), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_1142), .A2(n_1148), .B1(n_1151), .B2(n_1152), .C(n_1153), .Y(n_1156) );
NOR3xp33_ASAP7_75t_SL g1157 ( .A(n_1017), .B(n_1014), .C(n_949), .Y(n_1157) );
NAND4xp25_ASAP7_75t_L g1158 ( .A(n_1155), .B(n_1145), .C(n_1010), .D(n_975), .Y(n_1158) );
NAND4xp25_ASAP7_75t_L g1159 ( .A(n_1154), .B(n_1145), .C(n_1010), .D(n_975), .Y(n_1159) );
NOR3xp33_ASAP7_75t_SL g1160 ( .A(n_1156), .B(n_968), .C(n_925), .Y(n_1160) );
AND2x2_ASAP7_75t_L g1161 ( .A(n_1160), .B(n_1157), .Y(n_1161) );
XNOR2x1_ASAP7_75t_L g1162 ( .A(n_1159), .B(n_977), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_1158), .Y(n_1163) );
INVx1_ASAP7_75t_SL g1164 ( .A(n_1163), .Y(n_1164) );
OAI22xp5_ASAP7_75t_SL g1165 ( .A1(n_1164), .A2(n_1161), .B1(n_1162), .B2(n_957), .Y(n_1165) );
OA22x2_ASAP7_75t_L g1166 ( .A1(n_1165), .A2(n_921), .B1(n_1018), .B2(n_1020), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1166), .Y(n_1167) );
AOI21xp5_ASAP7_75t_L g1168 ( .A1(n_1167), .A2(n_967), .B(n_955), .Y(n_1168) );
OAI21xp33_ASAP7_75t_L g1169 ( .A1(n_1168), .A2(n_967), .B(n_979), .Y(n_1169) );
AOI21xp33_ASAP7_75t_L g1170 ( .A1(n_1169), .A2(n_967), .B(n_955), .Y(n_1170) );
endmodule