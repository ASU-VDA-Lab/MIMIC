module fake_netlist_1_12528_n_662 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_39, n_662);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_39;
output n_662;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_23), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_31), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_43), .Y(n_99) );
BUFx3_ASAP7_75t_L g100 ( .A(n_28), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_92), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_42), .Y(n_102) );
BUFx2_ASAP7_75t_L g103 ( .A(n_54), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_13), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_8), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_91), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_83), .Y(n_108) );
BUFx5_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_21), .B(n_86), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_1), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_79), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_53), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_41), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_45), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_46), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_55), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_61), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_37), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_38), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_29), .Y(n_122) );
BUFx6f_ASAP7_75t_L g123 ( .A(n_18), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_17), .Y(n_124) );
INVx1_ASAP7_75t_SL g125 ( .A(n_76), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_93), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_8), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_68), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_9), .Y(n_130) );
CKINVDCx14_ASAP7_75t_R g131 ( .A(n_62), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_20), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_81), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_2), .Y(n_134) );
INVx1_ASAP7_75t_SL g135 ( .A(n_78), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_30), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_19), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_0), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_58), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_95), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
OAI22x1_ASAP7_75t_R g143 ( .A1(n_134), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_116), .B(n_3), .Y(n_144) );
OAI22xp5_ASAP7_75t_L g145 ( .A1(n_124), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_98), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_124), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_130), .B(n_6), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_100), .B(n_7), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_109), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_109), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_101), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_109), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_100), .B(n_7), .Y(n_154) );
INVx6_ASAP7_75t_L g155 ( .A(n_109), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_95), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_130), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_128), .B(n_9), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_137), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_159) );
INVx1_ASAP7_75t_SL g160 ( .A(n_157), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_140), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_140), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_150), .Y(n_165) );
BUFx10_ASAP7_75t_L g166 ( .A(n_155), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_142), .B(n_121), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_142), .B(n_105), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_141), .B(n_99), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_141), .B(n_99), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_155), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_154), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g175 ( .A(n_142), .B(n_137), .Y(n_175) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_146), .A2(n_110), .B1(n_127), .B2(n_97), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_154), .A2(n_112), .B1(n_104), .B2(n_123), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_155), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g181 ( .A(n_148), .B(n_138), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_156), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_144), .B(n_131), .Y(n_185) );
AND2x4_ASAP7_75t_SL g186 ( .A(n_144), .B(n_133), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_185), .B(n_146), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_173), .B(n_158), .Y(n_189) );
INVx3_ASAP7_75t_L g190 ( .A(n_173), .Y(n_190) );
AND2x2_ASAP7_75t_SL g191 ( .A(n_186), .B(n_158), .Y(n_191) );
AOI22xp33_ASAP7_75t_SL g192 ( .A1(n_186), .A2(n_139), .B1(n_133), .B2(n_159), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_173), .B(n_158), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_173), .B(n_158), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_167), .B(n_169), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_167), .B(n_152), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_185), .B(n_152), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_185), .B(n_149), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_177), .B(n_149), .Y(n_201) );
NOR2x1_ASAP7_75t_L g202 ( .A(n_175), .B(n_139), .Y(n_202) );
INVxp67_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_167), .B(n_149), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_160), .B(n_138), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_177), .B(n_151), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_175), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_177), .B(n_96), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_184), .B(n_96), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_184), .B(n_102), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_184), .B(n_153), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_171), .Y(n_213) );
OR2x6_ASAP7_75t_L g214 ( .A(n_181), .B(n_145), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g215 ( .A1(n_178), .A2(n_147), .B1(n_106), .B2(n_155), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_181), .B(n_123), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_186), .B(n_102), .Y(n_217) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_184), .B(n_123), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_171), .B(n_107), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_176), .B(n_107), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_172), .B(n_108), .Y(n_221) );
INVx3_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_172), .A2(n_153), .B(n_120), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_176), .B(n_108), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_195), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_197), .Y(n_226) );
INVx2_ASAP7_75t_SL g227 ( .A(n_205), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_190), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_203), .B(n_172), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_189), .A2(n_179), .B(n_165), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_213), .B(n_164), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_189), .A2(n_179), .B(n_165), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_193), .A2(n_179), .B(n_180), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_207), .B(n_113), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_198), .B(n_180), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_196), .B(n_166), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_192), .B(n_129), .C(n_126), .Y(n_237) );
OAI22xp5_ASAP7_75t_L g238 ( .A1(n_188), .A2(n_122), .B1(n_117), .B2(n_115), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_193), .A2(n_120), .B(n_132), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_204), .B(n_166), .Y(n_240) );
O2A1O1Ixp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_118), .B(n_132), .C(n_136), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_194), .A2(n_136), .B(n_118), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_199), .B(n_166), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_194), .A2(n_114), .B(n_183), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_201), .A2(n_114), .B(n_135), .C(n_125), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_201), .A2(n_128), .B(n_111), .C(n_143), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_216), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_206), .A2(n_162), .B(n_183), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_222), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_191), .A2(n_123), .B1(n_95), .B2(n_119), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_217), .B(n_166), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_222), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_206), .A2(n_163), .B(n_183), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_190), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_190), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_212), .A2(n_162), .B(n_182), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_225), .B(n_216), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_249), .Y(n_259) );
AO32x2_ASAP7_75t_L g260 ( .A1(n_250), .A2(n_215), .A3(n_218), .B1(n_191), .B2(n_216), .Y(n_260) );
AOI31xp67_ASAP7_75t_L g261 ( .A1(n_228), .A2(n_163), .A3(n_174), .B(n_182), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_237), .A2(n_214), .B1(n_202), .B2(n_219), .Y(n_262) );
OA21x2_ASAP7_75t_L g263 ( .A1(n_241), .A2(n_223), .B(n_212), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_231), .A2(n_209), .B(n_210), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_227), .A2(n_214), .B1(n_220), .B2(n_224), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_226), .A2(n_214), .B1(n_211), .B2(n_221), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_208), .B(n_218), .Y(n_267) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_239), .A2(n_163), .B(n_182), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_229), .Y(n_269) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_248), .A2(n_208), .B(n_174), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_235), .B(n_214), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_208), .B(n_174), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_249), .Y(n_273) );
NOR2xp67_ASAP7_75t_L g274 ( .A(n_250), .B(n_10), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_229), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_255), .B(n_109), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_238), .B(n_11), .Y(n_277) );
AO32x2_ASAP7_75t_L g278 ( .A1(n_238), .A2(n_143), .A3(n_156), .B1(n_109), .B2(n_95), .Y(n_278) );
INVx1_ASAP7_75t_SL g279 ( .A(n_249), .Y(n_279) );
O2A1O1Ixp5_ASAP7_75t_SL g280 ( .A1(n_256), .A2(n_156), .B(n_109), .C(n_187), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_247), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_252), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_261), .Y(n_283) );
BUFx2_ASAP7_75t_L g284 ( .A(n_259), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_270), .A2(n_257), .B(n_253), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_276), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_258), .B(n_255), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_271), .B(n_243), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_271), .B(n_243), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_259), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_264), .A2(n_236), .B(n_232), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_266), .B(n_252), .Y(n_292) );
AO31x2_ASAP7_75t_L g293 ( .A1(n_267), .A2(n_242), .A3(n_244), .B(n_233), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_270), .A2(n_245), .B(n_254), .Y(n_294) );
AO31x2_ASAP7_75t_L g295 ( .A1(n_277), .A2(n_236), .A3(n_240), .B(n_251), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_276), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_265), .B(n_252), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_272), .A2(n_240), .B(n_234), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_258), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_258), .B(n_234), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_259), .B(n_168), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_259), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_274), .A2(n_246), .B(n_162), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_286), .B(n_260), .Y(n_305) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_283), .A2(n_262), .B(n_280), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
OA21x2_ASAP7_75t_L g308 ( .A1(n_283), .A2(n_280), .B(n_269), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_302), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_302), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_286), .B(n_260), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_296), .B(n_260), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_302), .Y(n_313) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_291), .A2(n_268), .B(n_273), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_284), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_285), .A2(n_273), .B(n_161), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_297), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_295), .B(n_260), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_285), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_295), .B(n_260), .Y(n_321) );
BUFx12f_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_297), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_295), .B(n_278), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_295), .B(n_278), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_284), .B(n_268), .Y(n_326) );
OA21x2_ASAP7_75t_L g327 ( .A1(n_294), .A2(n_161), .B(n_282), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_290), .B(n_268), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
OR2x2_ASAP7_75t_L g330 ( .A(n_288), .B(n_275), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_322), .B(n_298), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_315), .Y(n_334) );
INVx2_ASAP7_75t_SL g335 ( .A(n_315), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_318), .B(n_292), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_316), .B(n_295), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_331), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_315), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_309), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_309), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_316), .B(n_295), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_305), .B(n_304), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_326), .B(n_304), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_305), .B(n_304), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_305), .B(n_304), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_305), .B(n_299), .Y(n_351) );
OR2x6_ASAP7_75t_L g352 ( .A(n_319), .B(n_292), .Y(n_352) );
BUFx3_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_322), .A2(n_300), .B1(n_289), .B2(n_288), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_311), .B(n_299), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_311), .B(n_278), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_318), .B(n_323), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_318), .B(n_289), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_310), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_311), .B(n_278), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_310), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_310), .Y(n_364) );
INVxp67_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_313), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_312), .B(n_300), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_323), .B(n_300), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_313), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
NAND2x1p5_ASAP7_75t_SL g372 ( .A(n_324), .B(n_293), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_312), .B(n_287), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_323), .B(n_324), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_320), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_312), .B(n_287), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_351), .B(n_324), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_374), .B(n_325), .Y(n_378) );
INVx2_ASAP7_75t_SL g379 ( .A(n_334), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_360), .B(n_322), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_349), .B(n_319), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_340), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_349), .B(n_319), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_349), .B(n_321), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_335), .B(n_322), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_373), .B(n_321), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_355), .B(n_325), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_373), .B(n_321), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
CKINVDCx8_ASAP7_75t_R g393 ( .A(n_348), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_358), .B(n_330), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_347), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_340), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_358), .B(n_330), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_376), .B(n_326), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_340), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_347), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_362), .B(n_330), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_343), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_346), .B(n_326), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
NOR2x1_ASAP7_75t_SL g406 ( .A(n_335), .B(n_329), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_374), .B(n_326), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_348), .B(n_326), .Y(n_408) );
INVxp33_ASAP7_75t_L g409 ( .A(n_338), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_334), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_365), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_360), .B(n_329), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_367), .B(n_329), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_369), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_356), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_343), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_334), .Y(n_417) );
AND2x4_ASAP7_75t_L g418 ( .A(n_348), .B(n_328), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_350), .B(n_328), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_372), .B(n_328), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_367), .B(n_332), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_343), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_344), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_336), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_336), .B(n_332), .Y(n_425) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_353), .B(n_332), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_353), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_356), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_335), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_357), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_357), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_366), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_392), .Y(n_434) );
INVx2_ASAP7_75t_SL g435 ( .A(n_410), .Y(n_435) );
INVx1_ASAP7_75t_SL g436 ( .A(n_410), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_392), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_383), .B(n_337), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_383), .B(n_386), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_411), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_398), .B(n_341), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_407), .B(n_352), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_380), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_398), .B(n_341), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_407), .B(n_352), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_378), .B(n_352), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_386), .B(n_345), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_389), .B(n_352), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_389), .B(n_352), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_387), .B(n_345), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_391), .B(n_404), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_379), .B(n_348), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_391), .B(n_352), .Y(n_454) );
AND3x2_ASAP7_75t_L g455 ( .A(n_417), .B(n_333), .C(n_344), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_406), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_381), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_387), .B(n_372), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_384), .Y(n_459) );
INVx3_ASAP7_75t_L g460 ( .A(n_393), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_424), .B(n_372), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_378), .B(n_344), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_413), .B(n_361), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_419), .B(n_328), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_385), .Y(n_465) );
AO22x1_ASAP7_75t_L g466 ( .A1(n_427), .A2(n_361), .B1(n_370), .B2(n_368), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_395), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_421), .B(n_361), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_396), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_377), .B(n_363), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_400), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_402), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_379), .B(n_363), .Y(n_473) );
INVxp67_ASAP7_75t_L g474 ( .A(n_406), .Y(n_474) );
AND2x2_ASAP7_75t_SL g475 ( .A(n_408), .B(n_333), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_405), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_382), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_399), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_390), .B(n_364), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_412), .B(n_364), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_394), .B(n_368), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_409), .B(n_354), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_397), .B(n_368), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_414), .B(n_354), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_409), .B(n_12), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_415), .B(n_375), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_401), .B(n_375), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_429), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_426), .B(n_320), .C(n_308), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_425), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_415), .B(n_314), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_399), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_388), .B(n_327), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_432), .B(n_314), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_432), .B(n_314), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_408), .B(n_314), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_433), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_393), .B(n_320), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_408), .B(n_320), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_403), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_418), .B(n_314), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_418), .B(n_308), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_433), .B(n_308), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_439), .B(n_490), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_444), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_452), .B(n_420), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_438), .B(n_420), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_440), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_461), .B(n_428), .Y(n_509) );
OAI22xp33_ASAP7_75t_SL g510 ( .A1(n_477), .A2(n_430), .B1(n_431), .B2(n_423), .Y(n_510) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_475), .B(n_456), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_461), .B(n_403), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_438), .B(n_416), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_448), .B(n_416), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_448), .B(n_422), .Y(n_516) );
AND2x4_ASAP7_75t_L g517 ( .A(n_456), .B(n_422), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_474), .B(n_423), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_457), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_465), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_436), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_467), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_471), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_451), .B(n_308), .Y(n_524) );
INVxp67_ASAP7_75t_L g525 ( .A(n_435), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_497), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_451), .B(n_306), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_434), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_437), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_474), .A2(n_317), .B1(n_287), .B2(n_327), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g531 ( .A1(n_485), .A2(n_281), .B(n_287), .C(n_308), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_472), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_462), .B(n_306), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_458), .B(n_484), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_473), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_459), .Y(n_537) );
OAI21xp5_ASAP7_75t_SL g538 ( .A1(n_460), .A2(n_301), .B(n_15), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_458), .B(n_482), .Y(n_539) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_460), .A2(n_317), .B1(n_327), .B2(n_306), .Y(n_540) );
NOR2x1_ASAP7_75t_L g541 ( .A(n_493), .B(n_327), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_463), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_468), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_470), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_453), .B(n_293), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_480), .Y(n_547) );
AND2x4_ASAP7_75t_L g548 ( .A(n_453), .B(n_293), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_481), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_483), .Y(n_550) );
INVx2_ASAP7_75t_SL g551 ( .A(n_442), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_459), .Y(n_552) );
OAI33xp33_ASAP7_75t_L g553 ( .A1(n_488), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_486), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_487), .B(n_14), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_445), .B(n_293), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_488), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_464), .B(n_293), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_447), .B(n_16), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g560 ( .A1(n_485), .A2(n_301), .B(n_279), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_469), .Y(n_561) );
AOI31xp33_ASAP7_75t_L g562 ( .A1(n_525), .A2(n_498), .A3(n_443), .B(n_446), .Y(n_562) );
OAI22xp33_ASAP7_75t_SL g563 ( .A1(n_511), .A2(n_498), .B1(n_491), .B2(n_495), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_538), .A2(n_455), .B(n_454), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_538), .A2(n_475), .B(n_489), .Y(n_565) );
AOI211x1_ASAP7_75t_L g566 ( .A1(n_539), .A2(n_466), .B(n_449), .C(n_450), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_506), .B(n_502), .Y(n_568) );
OAI322xp33_ASAP7_75t_L g569 ( .A1(n_555), .A2(n_491), .A3(n_494), .B1(n_495), .B2(n_503), .C1(n_496), .C2(n_501), .Y(n_569) );
OAI21xp33_ASAP7_75t_L g570 ( .A1(n_510), .A2(n_494), .B(n_499), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_521), .B(n_499), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_517), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_521), .Y(n_573) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_510), .A2(n_503), .B(n_500), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_554), .B(n_469), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_536), .B(n_441), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_519), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_524), .B(n_478), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_520), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_522), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_511), .A2(n_492), .B(n_455), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_523), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_504), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_527), .B(n_492), .Y(n_584) );
OAI322xp33_ASAP7_75t_L g585 ( .A1(n_535), .A2(n_161), .A3(n_301), .B1(n_187), .B2(n_168), .C1(n_293), .C2(n_32), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_557), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_536), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_508), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_514), .Y(n_589) );
NAND3xp33_ASAP7_75t_L g590 ( .A(n_531), .B(n_263), .C(n_187), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_517), .Y(n_591) );
NAND4xp25_ASAP7_75t_L g592 ( .A(n_559), .B(n_22), .C(n_24), .D(n_26), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_532), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_546), .B(n_27), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_534), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_526), .Y(n_596) );
O2A1O1Ixp33_ASAP7_75t_L g597 ( .A1(n_553), .A2(n_263), .B(n_35), .C(n_36), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_509), .B(n_263), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_528), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_515), .B(n_187), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_547), .B(n_34), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_529), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_542), .Y(n_603) );
AOI21xp33_ASAP7_75t_L g604 ( .A1(n_597), .A2(n_505), .B(n_560), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_583), .B(n_543), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g606 ( .A1(n_564), .A2(n_518), .B(n_541), .Y(n_606) );
NOR2xp33_ASAP7_75t_R g607 ( .A(n_573), .B(n_551), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_566), .A2(n_544), .B1(n_545), .B2(n_549), .C(n_550), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_565), .A2(n_546), .B1(n_548), .B2(n_556), .Y(n_609) );
OAI31xp33_ASAP7_75t_L g610 ( .A1(n_570), .A2(n_548), .A3(n_558), .B(n_513), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g611 ( .A1(n_562), .A2(n_516), .B(n_512), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_575), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_563), .A2(n_530), .B(n_540), .C(n_533), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g614 ( .A1(n_581), .A2(n_561), .B1(n_552), .B2(n_537), .C(n_168), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_569), .A2(n_168), .B(n_39), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_587), .A2(n_168), .B1(n_40), .B2(n_44), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_575), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_597), .A2(n_47), .B(n_48), .Y(n_618) );
AOI31xp33_ASAP7_75t_L g619 ( .A1(n_574), .A2(n_49), .A3(n_50), .B(n_51), .Y(n_619) );
AOI211xp5_ASAP7_75t_L g620 ( .A1(n_592), .A2(n_52), .B(n_56), .C(n_57), .Y(n_620) );
AOI211xp5_ASAP7_75t_L g621 ( .A1(n_571), .A2(n_59), .B(n_60), .C(n_63), .Y(n_621) );
O2A1O1Ixp33_ASAP7_75t_L g622 ( .A1(n_586), .A2(n_64), .B(n_65), .C(n_66), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_578), .A2(n_67), .B(n_69), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g624 ( .A1(n_603), .A2(n_70), .B1(n_71), .B2(n_73), .C1(n_74), .C2(n_75), .Y(n_624) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_567), .A2(n_77), .B1(n_80), .B2(n_82), .C(n_85), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_601), .A2(n_87), .B(n_89), .C(n_90), .Y(n_626) );
NAND3xp33_ASAP7_75t_SL g627 ( .A(n_590), .B(n_601), .C(n_572), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_589), .B(n_584), .Y(n_628) );
AOI33xp33_ASAP7_75t_L g629 ( .A1(n_577), .A2(n_593), .A3(n_595), .B1(n_579), .B2(n_580), .B3(n_582), .Y(n_629) );
OAI221xp5_ASAP7_75t_SL g630 ( .A1(n_591), .A2(n_584), .B1(n_588), .B2(n_576), .C(n_599), .Y(n_630) );
OAI211xp5_ASAP7_75t_SL g631 ( .A1(n_596), .A2(n_602), .B(n_600), .C(n_598), .Y(n_631) );
AOI322xp5_ASAP7_75t_L g632 ( .A1(n_568), .A2(n_585), .A3(n_594), .B1(n_598), .B2(n_570), .C1(n_539), .C2(n_567), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_594), .B(n_573), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_583), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_566), .A2(n_569), .B1(n_570), .B2(n_562), .C(n_539), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_636), .B(n_604), .C(n_618), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_614), .B(n_604), .C(n_606), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_609), .B(n_607), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_635), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_634), .B(n_630), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g642 ( .A(n_632), .B(n_613), .C(n_615), .Y(n_642) );
NAND4xp75_ASAP7_75t_L g643 ( .A(n_610), .B(n_623), .C(n_633), .D(n_625), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_605), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_637), .B(n_629), .Y(n_645) );
AOI221x1_ASAP7_75t_L g646 ( .A1(n_637), .A2(n_616), .B1(n_631), .B2(n_611), .C(n_627), .Y(n_646) );
NAND3xp33_ASAP7_75t_SL g647 ( .A(n_638), .B(n_620), .C(n_621), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_644), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_640), .B(n_617), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_645), .B(n_639), .Y(n_650) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_648), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_649), .Y(n_652) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_652), .B(n_643), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_650), .A2(n_642), .B(n_646), .Y(n_654) );
BUFx8_ASAP7_75t_L g655 ( .A(n_653), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_654), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_651), .B(n_641), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_655), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_647), .B1(n_612), .B2(n_608), .Y(n_659) );
AO21x2_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_657), .B(n_619), .Y(n_660) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_622), .B(n_624), .Y(n_661) );
AOI21xp33_ASAP7_75t_SL g662 ( .A1(n_661), .A2(n_628), .B(n_626), .Y(n_662) );
endmodule