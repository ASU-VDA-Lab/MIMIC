module real_jpeg_13302_n_18 (n_17, n_8, n_251, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_251;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_68;
wire n_247;
wire n_146;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_188;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_3),
.A2(n_30),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_3),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_4),
.A2(n_66),
.B1(n_67),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_4),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_4),
.A2(n_61),
.B1(n_64),
.B2(n_72),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_4),
.A2(n_45),
.B1(n_47),
.B2(n_72),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_4),
.A2(n_30),
.B1(n_38),
.B2(n_72),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_5),
.A2(n_61),
.B1(n_64),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_5),
.A2(n_66),
.B1(n_67),
.B2(n_81),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_5),
.A2(n_45),
.B1(n_47),
.B2(n_81),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_5),
.A2(n_30),
.B1(n_38),
.B2(n_81),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_7),
.A2(n_66),
.B1(n_67),
.B2(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_7),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_7),
.A2(n_61),
.B1(n_64),
.B2(n_111),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_7),
.A2(n_45),
.B1(n_47),
.B2(n_111),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_7),
.A2(n_30),
.B1(n_38),
.B2(n_111),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_8),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_8),
.A2(n_44),
.B1(n_61),
.B2(n_64),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_8),
.A2(n_30),
.B1(n_38),
.B2(n_44),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_9),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_9),
.A2(n_45),
.B1(n_47),
.B2(n_70),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_9),
.A2(n_30),
.B1(n_38),
.B2(n_70),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_11),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_11),
.A2(n_37),
.B1(n_45),
.B2(n_47),
.Y(n_87)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_13),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_13),
.B(n_114),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_66),
.B(n_167),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_45),
.B1(n_47),
.B2(n_102),
.Y(n_185)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_13),
.A2(n_47),
.B(n_51),
.C(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_13),
.B(n_107),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_13),
.B(n_34),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_13),
.B(n_88),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_13),
.A2(n_64),
.B(n_75),
.C(n_222),
.Y(n_221)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_15),
.A2(n_45),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_15),
.A2(n_30),
.B1(n_38),
.B2(n_55),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_15),
.A2(n_55),
.B1(n_61),
.B2(n_64),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_16),
.A2(n_30),
.B1(n_38),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_16),
.Y(n_92)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_135),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_133),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_115),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_22),
.B(n_115),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_94),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_23),
.A2(n_24),
.B1(n_83),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_56),
.B2(n_57),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_25),
.B(n_58),
.C(n_73),
.Y(n_116)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_41),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_39),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_28),
.A2(n_33),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_29),
.A2(n_34),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_29),
.A2(n_34),
.B1(n_36),
.B2(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_29),
.A2(n_34),
.B(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_29),
.A2(n_34),
.B1(n_98),
.B2(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_29),
.A2(n_34),
.B1(n_149),
.B2(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_29),
.A2(n_34),
.B1(n_161),
.B2(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_29),
.A2(n_34),
.B1(n_102),
.B2(n_207),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_29),
.A2(n_34),
.B1(n_200),
.B2(n_207),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_30),
.B(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_38),
.A2(n_52),
.B(n_102),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_43),
.A2(n_49),
.B1(n_88),
.B2(n_153),
.Y(n_170)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_47),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_45),
.A2(n_64),
.A3(n_77),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_47),
.B(n_78),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_48),
.A2(n_53),
.B1(n_152),
.B2(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_49),
.A2(n_87),
.B1(n_88),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_49),
.A2(n_88),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_49),
.A2(n_88),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_49),
.A2(n_88),
.B1(n_186),
.B2(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_73),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_69),
.B2(n_71),
.Y(n_58)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_59),
.A2(n_60),
.B1(n_71),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_59),
.A2(n_60),
.B1(n_110),
.B2(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_64),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_63),
.A3(n_66),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_61),
.B(n_102),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_64),
.Y(n_100)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_102),
.Y(n_101)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_74),
.A2(n_79),
.B1(n_82),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_74),
.A2(n_79),
.B1(n_105),
.B2(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_75),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_75),
.A2(n_107),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_79),
.A2(n_143),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_83),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_93),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_93),
.Y(n_126)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_94),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_108),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_95),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_101),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_103),
.B(n_108),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_123),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI221xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.C(n_251),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_235),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_178),
.B(n_234),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_162),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_139),
.B(n_162),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_150),
.C(n_154),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_140),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_147),
.C(n_148),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_150),
.A2(n_154),
.B1(n_155),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_156),
.A2(n_157),
.B1(n_160),
.B2(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_158),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_173),
.B2(n_177),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_174),
.C(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_165),
.B(n_169),
.C(n_172),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_228),
.B(n_233),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_216),
.B(n_227),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_196),
.B(n_215),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_182),
.B(n_189),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_183),
.A2(n_184),
.B1(n_187),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_192),
.C(n_194),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_204),
.B(n_214),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_198),
.B(n_202),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_210),
.B(n_213),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_211),
.B(n_212),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_218),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_223),
.C(n_225),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_237),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_240),
.C(n_241),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);


endmodule