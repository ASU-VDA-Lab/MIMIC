module fake_netlist_5_311_n_2114 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_211, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_2114);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2114;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2009;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_433;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1996;
wire n_597;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_54),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_182),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_93),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_77),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_165),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_103),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_67),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_41),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_213),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_140),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_53),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_51),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_151),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_184),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_28),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_97),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_123),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_43),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_51),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_4),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_89),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_10),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_23),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_68),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_61),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_2),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_209),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_52),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_86),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_100),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_124),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_88),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_116),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_118),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_104),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_160),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_2),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_139),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_49),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_126),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_27),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_166),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_25),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_169),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_85),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_107),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_27),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_12),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_94),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_167),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_70),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_47),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_145),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_171),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_152),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_66),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_0),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_115),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_72),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_193),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_204),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_63),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_153),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_125),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_122),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_98),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_155),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_109),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_159),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_0),
.Y(n_298)
);

CKINVDCx12_ASAP7_75t_R g299 ( 
.A(n_83),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_76),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_37),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_15),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_135),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_25),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_60),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_23),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_69),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_121),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_57),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_44),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_67),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_15),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_111),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_91),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_28),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_120),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_37),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_40),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_79),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_129),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_77),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_92),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_73),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_205),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_82),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_59),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_199),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_196),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_210),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_154),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_142),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_58),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_18),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_8),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_62),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_81),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_79),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_90),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_26),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_10),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_22),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_110),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_80),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_84),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_179),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_87),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_176),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_170),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_21),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_141),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_128),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_52),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_18),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_66),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_45),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_201),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_33),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_83),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_127),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_192),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_55),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_173),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_99),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_102),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_80),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_168),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_95),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_31),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_50),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_13),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_36),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_14),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_34),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_50),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_117),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_58),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_187),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_113),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_130),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_39),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_183),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_114),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_131),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_61),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_191),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_190),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_69),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_11),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_73),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_206),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_22),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_63),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_34),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_62),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_137),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_14),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_208),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_40),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_30),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_39),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_8),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_4),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_148),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_132),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_157),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_175),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_20),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_38),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_144),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_186),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_200),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_1),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_178),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_96),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_3),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_57),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_162),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_119),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_53),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_20),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_246),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_227),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_246),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_274),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g427 ( 
.A(n_328),
.B(n_1),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_222),
.B(n_3),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_286),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_303),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_286),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_286),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_344),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_225),
.B(n_5),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_286),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_286),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_361),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_235),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_286),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_384),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_416),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_274),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_286),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_355),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_357),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_286),
.Y(n_446)
);

BUFx6f_ASAP7_75t_SL g447 ( 
.A(n_330),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_286),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_230),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_230),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_230),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_230),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_230),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_357),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_224),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_224),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_412),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_228),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_412),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_228),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_231),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_235),
.Y(n_462)
);

INVxp33_ASAP7_75t_SL g463 ( 
.A(n_355),
.Y(n_463)
);

INVxp67_ASAP7_75t_SL g464 ( 
.A(n_269),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_214),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_218),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_296),
.B(n_6),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_299),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_273),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g470 ( 
.A(n_273),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_253),
.B(n_6),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_231),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_223),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_216),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_233),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_233),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_229),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_329),
.B(n_7),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_241),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_289),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_243),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_217),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_219),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_296),
.B(n_7),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_239),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_220),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_230),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_247),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_250),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_221),
.Y(n_490)
);

BUFx2_ASAP7_75t_SL g491 ( 
.A(n_330),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_226),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_239),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_248),
.B(n_9),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_248),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_252),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_236),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_238),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_269),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_299),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_261),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_314),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_262),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_264),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_242),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_R g506 ( 
.A(n_249),
.B(n_101),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_252),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_251),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_254),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_255),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_256),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_279),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_283),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_225),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_255),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_258),
.B(n_9),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_222),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_258),
.B(n_13),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_284),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_263),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_263),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_257),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_268),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_293),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_260),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_298),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_265),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_418),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_418),
.B(n_16),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_302),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_305),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_L g532 ( 
.A(n_466),
.B(n_310),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_449),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_446),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_449),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_466),
.B(n_312),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_450),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_423),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_451),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

AND3x2_ASAP7_75t_L g542 ( 
.A(n_471),
.B(n_275),
.C(n_270),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_455),
.B(n_314),
.Y(n_543)
);

OA21x2_ASAP7_75t_L g544 ( 
.A1(n_452),
.A2(n_282),
.B(n_268),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_469),
.B(n_330),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_452),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_491),
.B(n_273),
.Y(n_547)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_447),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_453),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_453),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_487),
.Y(n_551)
);

AND2x4_ASAP7_75t_SL g552 ( 
.A(n_465),
.B(n_330),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_528),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_528),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_446),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_464),
.B(n_267),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_481),
.B(n_352),
.Y(n_559)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_429),
.A2(n_287),
.B(n_282),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_448),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_432),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_435),
.Y(n_564)
);

INVx5_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_436),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_499),
.B(n_502),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_439),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_514),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_456),
.B(n_399),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_480),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_514),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_458),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_460),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_461),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_472),
.B(n_276),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_476),
.B(n_277),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_491),
.B(n_273),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_485),
.Y(n_581)
);

CKINVDCx8_ASAP7_75t_R g582 ( 
.A(n_470),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_493),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_496),
.B(n_280),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_438),
.B(n_289),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_507),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_510),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_515),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_520),
.B(n_399),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_521),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_523),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_428),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_434),
.B(n_270),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_494),
.B(n_285),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_467),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_484),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_462),
.B(n_311),
.Y(n_598)
);

OA21x2_ASAP7_75t_L g599 ( 
.A1(n_516),
.A2(n_294),
.B(n_287),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_468),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_500),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_517),
.B(n_311),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_529),
.B(n_275),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_428),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_424),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_427),
.B(n_290),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_518),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_478),
.B(n_288),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_506),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_503),
.B(n_318),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_447),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_L g612 ( 
.A(n_473),
.B(n_319),
.Y(n_612)
);

AND3x2_ASAP7_75t_L g613 ( 
.A(n_444),
.B(n_290),
.C(n_281),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_423),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_447),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_477),
.B(n_291),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_477),
.B(n_292),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_565),
.B(n_479),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_556),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_565),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_566),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_596),
.B(n_597),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_556),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_566),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_560),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_566),
.Y(n_628)
);

BUFx8_ASAP7_75t_SL g629 ( 
.A(n_605),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_565),
.B(n_479),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_557),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_533),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_561),
.Y(n_635)
);

INVx6_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_561),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_597),
.B(n_488),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_543),
.B(n_294),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_534),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_596),
.B(n_488),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_534),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_565),
.B(n_489),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_534),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_533),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_596),
.B(n_489),
.Y(n_647)
);

AO21x2_ASAP7_75t_L g648 ( 
.A1(n_608),
.A2(n_322),
.B(n_317),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_596),
.B(n_364),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_563),
.Y(n_650)
);

NAND3xp33_ASAP7_75t_L g651 ( 
.A(n_607),
.B(n_322),
.C(n_317),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_563),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_539),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_533),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_565),
.B(n_501),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_564),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_609),
.B(n_463),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_566),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_607),
.B(n_501),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_566),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_535),
.Y(n_661)
);

NAND2xp33_ASAP7_75t_L g662 ( 
.A(n_607),
.B(n_504),
.Y(n_662)
);

INVx3_ASAP7_75t_L g663 ( 
.A(n_566),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_535),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_565),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_566),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_568),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_564),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_568),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_564),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_569),
.Y(n_671)
);

AND2x6_ASAP7_75t_L g672 ( 
.A(n_596),
.B(n_364),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_535),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_593),
.B(n_504),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_569),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_546),
.Y(n_676)
);

AND2x6_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_364),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_558),
.B(n_512),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_569),
.Y(n_679)
);

INVx1_ASAP7_75t_SL g680 ( 
.A(n_539),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_565),
.B(n_512),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_567),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_569),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_586),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_536),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_559),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_547),
.B(n_513),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_593),
.A2(n_482),
.B1(n_483),
.B2(n_474),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_546),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_572),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_546),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_536),
.Y(n_692)
);

INVx1_ASAP7_75t_SL g693 ( 
.A(n_614),
.Y(n_693)
);

OAI21xp33_ASAP7_75t_SL g694 ( 
.A1(n_593),
.A2(n_245),
.B(n_240),
.Y(n_694)
);

NAND2xp33_ASAP7_75t_SL g695 ( 
.A(n_545),
.B(n_457),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_558),
.B(n_513),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_609),
.B(n_486),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_547),
.B(n_519),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_553),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_553),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_572),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_553),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_L g703 ( 
.A(n_595),
.B(n_519),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_538),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_538),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_540),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_617),
.B(n_490),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_540),
.Y(n_708)
);

INVx4_ASAP7_75t_L g709 ( 
.A(n_568),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_617),
.B(n_492),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_541),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_580),
.A2(n_232),
.B1(n_237),
.B2(n_234),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_541),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_549),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_580),
.B(n_524),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_586),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_568),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_567),
.B(n_524),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_618),
.B(n_595),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_549),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_560),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_550),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_614),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_608),
.B(n_526),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_550),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_551),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_551),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_602),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_577),
.B(n_526),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_548),
.B(n_530),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_574),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_576),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_581),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_577),
.B(n_530),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_574),
.Y(n_735)
);

XOR2xp5_ASAP7_75t_L g736 ( 
.A(n_548),
.B(n_430),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_568),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_598),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_579),
.B(n_531),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_579),
.B(n_531),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_575),
.Y(n_741)
);

BUFx6f_ASAP7_75t_L g742 ( 
.A(n_581),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_618),
.B(n_616),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_552),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_575),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_616),
.B(n_497),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_581),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_599),
.A2(n_339),
.B1(n_351),
.B2(n_320),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_578),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_585),
.B(n_295),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_599),
.A2(n_396),
.B1(n_320),
.B2(n_351),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_585),
.B(n_297),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_604),
.B(n_425),
.Y(n_753)
);

AND2x6_ASAP7_75t_L g754 ( 
.A(n_615),
.B(n_364),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_578),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_606),
.B(n_309),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_606),
.B(n_315),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_616),
.B(n_425),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_598),
.B(n_426),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_324),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_576),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_571),
.B(n_339),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_583),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_576),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_583),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_588),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_552),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_606),
.B(n_542),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_604),
.B(n_426),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_571),
.B(n_396),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_588),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_624),
.A2(n_590),
.B(n_543),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_719),
.B(n_568),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_771),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_771),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_648),
.A2(n_599),
.B1(n_560),
.B2(n_544),
.Y(n_776)
);

AND2x6_ASAP7_75t_L g777 ( 
.A(n_721),
.B(n_627),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_L g778 ( 
.A(n_662),
.B(n_537),
.C(n_532),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_684),
.A2(n_600),
.B1(n_601),
.B2(n_582),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_682),
.B(n_599),
.Y(n_780)
);

NOR2x1_ASAP7_75t_R g781 ( 
.A(n_723),
.B(n_442),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_743),
.B(n_568),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_718),
.B(n_600),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_684),
.B(n_716),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_642),
.B(n_599),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_716),
.B(n_552),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_647),
.B(n_581),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_621),
.B(n_581),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_731),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_731),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_621),
.B(n_581),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_633),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_625),
.B(n_581),
.Y(n_794)
);

NOR2xp67_ASAP7_75t_L g795 ( 
.A(n_697),
.B(n_611),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_601),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_646),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_762),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_738),
.B(n_602),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_625),
.B(n_542),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_738),
.B(n_364),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_678),
.B(n_364),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_632),
.B(n_560),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_696),
.B(n_610),
.Y(n_804)
);

AO22x1_ASAP7_75t_L g805 ( 
.A1(n_659),
.A2(n_445),
.B1(n_454),
.B2(n_442),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_632),
.B(n_560),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_646),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_721),
.B(n_615),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_634),
.B(n_594),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_634),
.B(n_594),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_659),
.B(n_582),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_721),
.A2(n_590),
.B(n_543),
.C(n_612),
.Y(n_812)
);

AND2x6_ASAP7_75t_L g813 ( 
.A(n_627),
.B(n_615),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_654),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_729),
.B(n_498),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_734),
.B(n_349),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_629),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_638),
.B(n_602),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_739),
.B(n_349),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_740),
.B(n_349),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_654),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_635),
.B(n_594),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_735),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_638),
.B(n_349),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_620),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_650),
.B(n_349),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_635),
.B(n_594),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_620),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_735),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_650),
.B(n_397),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_661),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_741),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_688),
.B(n_698),
.C(n_687),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_661),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_652),
.B(n_397),
.Y(n_835)
);

AO221x1_ASAP7_75t_L g836 ( 
.A1(n_690),
.A2(n_397),
.B1(n_245),
.B2(n_259),
.C(n_266),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_741),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_723),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_637),
.B(n_620),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_649),
.B(n_611),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_745),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_637),
.B(n_603),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_657),
.B(n_505),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_674),
.B(n_707),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_630),
.B(n_603),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_630),
.B(n_603),
.Y(n_846)
);

OR2x2_ASAP7_75t_L g847 ( 
.A(n_753),
.B(n_445),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_745),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_674),
.B(n_508),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_703),
.A2(n_509),
.B1(n_527),
.B2(n_525),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_630),
.B(n_603),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_652),
.B(n_543),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_728),
.B(n_511),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_750),
.B(n_590),
.Y(n_854)
);

AOI22x1_ASAP7_75t_L g855 ( 
.A1(n_640),
.A2(n_454),
.B1(n_590),
.B2(n_571),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_752),
.B(n_397),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_749),
.B(n_584),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_768),
.B(n_397),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_640),
.B(n_582),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_749),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_641),
.B(n_522),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_664),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_759),
.B(n_753),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_755),
.B(n_584),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_755),
.B(n_584),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_641),
.B(n_587),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_690),
.B(n_215),
.Y(n_867)
);

NOR2xp67_ASAP7_75t_L g868 ( 
.A(n_710),
.B(n_589),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_763),
.B(n_587),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_636),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_769),
.B(n_244),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_763),
.B(n_587),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_643),
.B(n_592),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_765),
.B(n_592),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_765),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_643),
.B(n_592),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_636),
.A2(n_748),
.B1(n_751),
.B2(n_701),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_766),
.B(n_544),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_686),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_715),
.B(n_459),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_SL g881 ( 
.A(n_653),
.B(n_433),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_766),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_645),
.B(n_326),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_685),
.B(n_544),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_685),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_639),
.A2(n_651),
.B(n_645),
.C(n_671),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_R g887 ( 
.A(n_695),
.B(n_437),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_692),
.B(n_544),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_636),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_746),
.B(n_613),
.C(n_591),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_636),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_680),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_733),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_692),
.Y(n_894)
);

NOR2x1p5_ASAP7_75t_L g895 ( 
.A(n_770),
.B(n_321),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_705),
.B(n_544),
.Y(n_896)
);

INVx5_ASAP7_75t_L g897 ( 
.A(n_649),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_686),
.B(n_440),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_671),
.B(n_332),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_639),
.B(n_331),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_705),
.B(n_589),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_706),
.B(n_591),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_706),
.Y(n_903)
);

AOI221xp5_ASAP7_75t_L g904 ( 
.A1(n_712),
.A2(n_300),
.B1(n_417),
.B2(n_271),
.C(n_375),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_708),
.B(n_331),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_639),
.A2(n_347),
.B(n_388),
.C(n_413),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_664),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_708),
.B(n_340),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_651),
.B(n_756),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_673),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_673),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_711),
.B(n_340),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_676),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_733),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_758),
.A2(n_441),
.B1(n_348),
.B2(n_353),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_736),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_770),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_711),
.B(n_347),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_720),
.B(n_350),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_712),
.B(n_613),
.C(n_325),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_757),
.A2(n_388),
.B1(n_385),
.B2(n_380),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_686),
.B(n_323),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_676),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_720),
.B(n_350),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_722),
.B(n_366),
.Y(n_925)
);

BUFx6f_ASAP7_75t_L g926 ( 
.A(n_733),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_689),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_722),
.B(n_366),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_675),
.B(n_333),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_726),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_726),
.B(n_639),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_704),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_732),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_689),
.Y(n_934)
);

INVxp33_ASAP7_75t_L g935 ( 
.A(n_736),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_SL g936 ( 
.A(n_693),
.B(n_382),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_730),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_675),
.B(n_679),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_679),
.B(n_380),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_683),
.B(n_385),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_760),
.A2(n_368),
.B1(n_387),
.B2(n_383),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_788),
.A2(n_666),
.B(n_623),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_784),
.B(n_648),
.Y(n_943)
);

OAI321xp33_ASAP7_75t_L g944 ( 
.A1(n_904),
.A2(n_395),
.A3(n_338),
.B1(n_337),
.B2(n_336),
.C(n_335),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_780),
.A2(n_666),
.B(n_623),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_804),
.A2(n_619),
.B1(n_631),
.B2(n_644),
.Y(n_946)
);

AO21x1_ASAP7_75t_L g947 ( 
.A1(n_773),
.A2(n_802),
.B(n_816),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_804),
.B(n_686),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_772),
.A2(n_666),
.B(n_623),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_773),
.A2(n_666),
.B(n_623),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_783),
.A2(n_709),
.B(n_665),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_798),
.B(n_767),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_783),
.A2(n_709),
.B(n_665),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_786),
.A2(n_709),
.B(n_622),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_SL g955 ( 
.A(n_892),
.B(n_744),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_932),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_838),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_817),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_845),
.A2(n_709),
.B(n_622),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_844),
.A2(n_694),
.B(n_681),
.C(n_655),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_L g961 ( 
.A(n_784),
.B(n_694),
.C(n_341),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_867),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_909),
.B(n_683),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_885),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_818),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_825),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_846),
.A2(n_742),
.B(n_733),
.Y(n_967)
);

NOR2xp67_ASAP7_75t_SL g968 ( 
.A(n_897),
.B(n_413),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_863),
.A2(n_345),
.B(n_240),
.C(n_259),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_868),
.B(n_648),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_933),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_894),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_796),
.B(n_799),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_796),
.B(n_704),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_815),
.B(n_713),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_886),
.A2(n_668),
.B(n_656),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_774),
.B(n_713),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_877),
.A2(n_714),
.B1(n_725),
.B2(n_727),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_903),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_825),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_775),
.B(n_714),
.Y(n_981)
);

AO21x1_ASAP7_75t_L g982 ( 
.A1(n_802),
.A2(n_819),
.B(n_816),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_817),
.Y(n_983)
);

NOR3xp33_ASAP7_75t_L g984 ( 
.A(n_843),
.B(n_420),
.C(n_415),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_851),
.A2(n_854),
.B(n_812),
.Y(n_985)
);

INVx5_ASAP7_75t_L g986 ( 
.A(n_777),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_930),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_881),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_825),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_808),
.A2(n_668),
.B(n_656),
.Y(n_990)
);

NOR3xp33_ASAP7_75t_L g991 ( 
.A(n_843),
.B(n_420),
.C(n_415),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_790),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_782),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_791),
.B(n_725),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_823),
.B(n_727),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_931),
.A2(n_778),
.B1(n_863),
.B2(n_839),
.Y(n_996)
);

OR2x2_ASAP7_75t_L g997 ( 
.A(n_847),
.B(n_570),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_936),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_829),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_793),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_832),
.B(n_761),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_833),
.A2(n_337),
.B(n_421),
.C(n_398),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_897),
.B(n_658),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_887),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_837),
.B(n_764),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_L g1006 ( 
.A1(n_819),
.A2(n_764),
.B(n_761),
.C(n_737),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_841),
.B(n_670),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_809),
.A2(n_742),
.B(n_733),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_820),
.A2(n_670),
.B(n_272),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_848),
.B(n_658),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_797),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_860),
.B(n_658),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_875),
.B(n_660),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_882),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_897),
.B(n_660),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_810),
.A2(n_747),
.B(n_742),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_822),
.B(n_660),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_849),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_827),
.A2(n_747),
.B(n_742),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_842),
.B(n_663),
.Y(n_1020)
);

OAI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_884),
.A2(n_667),
.B(n_663),
.Y(n_1021)
);

O2A1O1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_785),
.A2(n_691),
.B(n_699),
.C(n_702),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_849),
.B(n_342),
.C(n_327),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_938),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_785),
.B(n_663),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_808),
.A2(n_699),
.B(n_691),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_893),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_777),
.B(n_667),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_893),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_777),
.B(n_667),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_887),
.Y(n_1031)
);

O2A1O1Ixp5_ASAP7_75t_L g1032 ( 
.A1(n_820),
.A2(n_737),
.B(n_669),
.C(n_702),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_888),
.A2(n_737),
.B(n_669),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_896),
.A2(n_700),
.B(n_555),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_852),
.A2(n_747),
.B(n_742),
.Y(n_1035)
);

AND2x2_ASAP7_75t_SL g1036 ( 
.A(n_815),
.B(n_266),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_803),
.A2(n_747),
.B(n_669),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_917),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_850),
.B(n_570),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_806),
.A2(n_700),
.B(n_573),
.Y(n_1040)
);

INVx4_ASAP7_75t_L g1041 ( 
.A(n_825),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_824),
.A2(n_306),
.B(n_272),
.C(n_278),
.Y(n_1042)
);

AO21x1_ASAP7_75t_L g1043 ( 
.A1(n_856),
.A2(n_801),
.B(n_858),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_897),
.B(n_747),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_777),
.B(n_649),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_828),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_777),
.B(n_649),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_922),
.A2(n_880),
.B(n_878),
.C(n_901),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_853),
.B(n_343),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_857),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_893),
.A2(n_628),
.B(n_626),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_828),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_893),
.A2(n_628),
.B(n_626),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_807),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_914),
.A2(n_628),
.B(n_626),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_864),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_824),
.B(n_649),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_828),
.B(n_626),
.Y(n_1058)
);

OAI21xp33_ASAP7_75t_L g1059 ( 
.A1(n_922),
.A2(n_356),
.B(n_346),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_853),
.B(n_573),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_902),
.B(n_828),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_776),
.A2(n_672),
.B(n_649),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_879),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_776),
.A2(n_672),
.B(n_649),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_779),
.B(n_626),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_871),
.B(n_359),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_914),
.A2(n_628),
.B(n_626),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_895),
.B(n_278),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_865),
.B(n_672),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_880),
.B(n_370),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_869),
.B(n_672),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_795),
.B(n_628),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_859),
.B(n_301),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_914),
.A2(n_628),
.B(n_717),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_872),
.B(n_672),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_914),
.A2(n_717),
.B(n_672),
.Y(n_1076)
);

NAND2xp33_ASAP7_75t_SL g1077 ( 
.A(n_787),
.B(n_358),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_874),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_926),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_800),
.B(n_672),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_937),
.A2(n_811),
.B1(n_787),
.B2(n_891),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_801),
.A2(n_386),
.B(n_304),
.C(n_306),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_805),
.B(n_371),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_866),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_905),
.B(n_677),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_926),
.B(n_717),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_908),
.B(n_677),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_912),
.B(n_677),
.Y(n_1088)
);

OAI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_789),
.A2(n_677),
.B(n_754),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_891),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_883),
.A2(n_677),
.B1(n_754),
.B2(n_362),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_889),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_866),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_814),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_926),
.A2(n_717),
.B(n_677),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_918),
.A2(n_307),
.B(n_421),
.C(n_386),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_926),
.B(n_717),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_873),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_792),
.A2(n_717),
.B(n_677),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_794),
.A2(n_369),
.B(n_392),
.Y(n_1100)
);

NAND2x1p5_ASAP7_75t_L g1101 ( 
.A(n_889),
.B(n_554),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_856),
.A2(n_365),
.B(n_406),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_919),
.B(n_754),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_924),
.B(n_754),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_899),
.A2(n_377),
.B(n_408),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_925),
.B(n_754),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_889),
.B(n_379),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_858),
.A2(n_554),
.B(n_555),
.C(n_301),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_928),
.B(n_754),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_859),
.A2(n_381),
.B1(n_405),
.B2(n_419),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_883),
.B(n_754),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_899),
.A2(n_407),
.B(n_411),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_873),
.A2(n_304),
.B(n_307),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_821),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_915),
.B(n_422),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_861),
.B(n_372),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_929),
.A2(n_308),
.B(n_313),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_L g1118 ( 
.A(n_813),
.B(n_373),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_929),
.B(n_374),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_876),
.A2(n_308),
.B(n_313),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_890),
.A2(n_316),
.B(n_334),
.C(n_335),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_870),
.A2(n_316),
.B(n_334),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_870),
.A2(n_876),
.B(n_862),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_861),
.B(n_376),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_906),
.A2(n_336),
.B(n_338),
.C(n_345),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_831),
.A2(n_354),
.B(n_360),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_813),
.A2(n_414),
.B1(n_410),
.B2(n_409),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_855),
.A2(n_404),
.B1(n_403),
.B2(n_402),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_834),
.B(n_378),
.Y(n_1129)
);

AO21x1_ASAP7_75t_L g1130 ( 
.A1(n_939),
.A2(n_354),
.B(n_360),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_907),
.A2(n_393),
.B(n_367),
.Y(n_1131)
);

INVx4_ASAP7_75t_L g1132 ( 
.A(n_986),
.Y(n_1132)
);

AOI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1034),
.A2(n_963),
.B(n_970),
.Y(n_1133)
);

AND2x6_ASAP7_75t_L g1134 ( 
.A(n_1045),
.B(n_889),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1024),
.B(n_813),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_973),
.B(n_813),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_964),
.Y(n_1137)
);

NOR2xp67_ASAP7_75t_SL g1138 ( 
.A(n_986),
.B(n_920),
.Y(n_1138)
);

OAI221xp5_ASAP7_75t_L g1139 ( 
.A1(n_1049),
.A2(n_898),
.B1(n_921),
.B2(n_941),
.C(n_935),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_965),
.B(n_813),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1036),
.B(n_940),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_1018),
.B(n_781),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_974),
.B(n_910),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_975),
.A2(n_840),
.B(n_927),
.C(n_923),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1036),
.A2(n_900),
.B1(n_916),
.B2(n_836),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_975),
.B(n_948),
.Y(n_1146)
);

OAI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_1049),
.A2(n_389),
.B(n_390),
.Y(n_1147)
);

INVxp67_ASAP7_75t_L g1148 ( 
.A(n_962),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_1041),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1048),
.A2(n_1116),
.B(n_1124),
.C(n_974),
.Y(n_1150)
);

HB1xp67_ASAP7_75t_L g1151 ( 
.A(n_957),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1041),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_972),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_948),
.B(n_911),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1070),
.B(n_913),
.Y(n_1155)
);

XNOR2xp5_ASAP7_75t_L g1156 ( 
.A(n_983),
.B(n_826),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1060),
.B(n_934),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1050),
.B(n_900),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1066),
.B(n_394),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1056),
.B(n_900),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_943),
.A2(n_398),
.B1(n_367),
.B2(n_391),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1116),
.B(n_400),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1124),
.B(n_401),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_971),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1059),
.B(n_900),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_985),
.A2(n_835),
.B(n_830),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_986),
.A2(n_395),
.B1(n_391),
.B2(n_393),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_979),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_986),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_957),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1078),
.B(n_900),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1081),
.B(n_826),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_952),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_945),
.A2(n_363),
.B(n_212),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_949),
.A2(n_1061),
.B(n_954),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_987),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1038),
.B(n_363),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1048),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_942),
.A2(n_202),
.B(n_198),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_984),
.A2(n_197),
.B1(n_195),
.B2(n_194),
.Y(n_1180)
);

INVx3_ASAP7_75t_SL g1181 ( 
.A(n_958),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_R g1182 ( 
.A(n_1063),
.B(n_188),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1062),
.A2(n_185),
.B(n_181),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_952),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1038),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_992),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_999),
.B(n_146),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1046),
.B(n_177),
.Y(n_1188)
);

NOR2xp67_ASAP7_75t_SL g1189 ( 
.A(n_944),
.B(n_19),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_955),
.B(n_164),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1014),
.B(n_138),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1073),
.B(n_21),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_988),
.B(n_24),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1073),
.B(n_24),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1023),
.B(n_29),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1026),
.A2(n_163),
.B(n_161),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_998),
.B(n_29),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1002),
.B(n_30),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1001),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_1004),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_991),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1115),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_R g1203 ( 
.A(n_1031),
.B(n_158),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1005),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_961),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1027),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1068),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_997),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_977),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1039),
.B(n_150),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1064),
.A2(n_149),
.B(n_147),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_1068),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1046),
.B(n_134),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_966),
.B(n_143),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1017),
.A2(n_133),
.B(n_112),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1027),
.Y(n_1216)
);

OAI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1002),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_946),
.B(n_996),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1020),
.A2(n_108),
.B(n_106),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_960),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1027),
.B(n_105),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1119),
.A2(n_1093),
.B(n_1084),
.C(n_1098),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_981),
.B(n_46),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_994),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_995),
.B(n_47),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1083),
.B(n_48),
.C(n_54),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1121),
.B(n_48),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_SL g1228 ( 
.A1(n_1107),
.A2(n_55),
.B(n_56),
.C(n_59),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_1129),
.Y(n_1229)
);

INVx1_ASAP7_75t_SL g1230 ( 
.A(n_1025),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1047),
.A2(n_56),
.B(n_60),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1021),
.A2(n_64),
.B(n_68),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_956),
.B(n_64),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1007),
.B(n_70),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1027),
.B(n_71),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_1121),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1077),
.A2(n_84),
.B1(n_72),
.B2(n_74),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_969),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1128),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1029),
.B(n_75),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1080),
.A2(n_76),
.B(n_78),
.C(n_81),
.Y(n_1241)
);

BUFx2_ASAP7_75t_R g1242 ( 
.A(n_1065),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_993),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1033),
.A2(n_78),
.B(n_82),
.Y(n_1244)
);

O2A1O1Ixp5_ASAP7_75t_SL g1245 ( 
.A1(n_1107),
.A2(n_963),
.B(n_1065),
.C(n_978),
.Y(n_1245)
);

BUFx8_ASAP7_75t_L g1246 ( 
.A(n_1029),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1110),
.B(n_1127),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1092),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_993),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1000),
.B(n_1011),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1029),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_969),
.B(n_1029),
.Y(n_1252)
);

OR2x6_ASAP7_75t_L g1253 ( 
.A(n_1079),
.B(n_966),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1028),
.A2(n_1030),
.B(n_959),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1000),
.Y(n_1255)
);

XOR2xp5_ASAP7_75t_L g1256 ( 
.A(n_1101),
.B(n_1091),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_950),
.A2(n_967),
.B(n_1008),
.Y(n_1257)
);

HB1xp67_ASAP7_75t_L g1258 ( 
.A(n_1092),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1105),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1011),
.B(n_1054),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_976),
.A2(n_1111),
.B(n_1022),
.C(n_1088),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1016),
.A2(n_1019),
.B(n_1037),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_947),
.A2(n_982),
.B(n_1043),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1096),
.B(n_1120),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1054),
.B(n_1114),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1126),
.A2(n_1096),
.B1(n_1052),
.B2(n_980),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_1094),
.B(n_1114),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1118),
.A2(n_1112),
.B1(n_1090),
.B2(n_1052),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1079),
.B(n_989),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1094),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1035),
.A2(n_951),
.B(n_953),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_980),
.A2(n_989),
.B1(n_1057),
.B2(n_1113),
.Y(n_1272)
);

AND2x2_ASAP7_75t_SL g1273 ( 
.A(n_1079),
.B(n_1013),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1130),
.A2(n_1009),
.A3(n_1040),
.B1(n_1125),
.B2(n_1032),
.Y(n_1274)
);

OR2x6_ASAP7_75t_SL g1275 ( 
.A(n_1010),
.B(n_1012),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1117),
.B(n_1090),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1079),
.B(n_1069),
.Y(n_1277)
);

O2A1O1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1042),
.A2(n_1082),
.B(n_1125),
.C(n_1122),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1102),
.B(n_1100),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_990),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1071),
.A2(n_1075),
.B1(n_1085),
.B2(n_1087),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1101),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1103),
.A2(n_1104),
.B1(n_1109),
.B2(n_1106),
.Y(n_1283)
);

NAND2x1_ASAP7_75t_L g1284 ( 
.A(n_1123),
.B(n_1076),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_SL g1285 ( 
.A1(n_1058),
.A2(n_1003),
.B(n_1015),
.C(n_1097),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1006),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1058),
.B(n_1044),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1131),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1170),
.Y(n_1289)
);

O2A1O1Ixp33_ASAP7_75t_SL g1290 ( 
.A1(n_1150),
.A2(n_1072),
.B(n_1044),
.C(n_1097),
.Y(n_1290)
);

AOI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1133),
.A2(n_1072),
.B(n_1099),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1200),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1218),
.A2(n_1089),
.B(n_1086),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1250),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1151),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1267),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_R g1297 ( 
.A(n_1259),
.B(n_1108),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1185),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1254),
.A2(n_1095),
.B(n_1051),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_SL g1300 ( 
.A1(n_1220),
.A2(n_1086),
.B(n_1053),
.C(n_1055),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_1182),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1181),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1239),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1255),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1261),
.A2(n_1067),
.A3(n_1074),
.B(n_968),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1209),
.B(n_1224),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1140),
.B(n_1184),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1175),
.A2(n_1257),
.B(n_1271),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1281),
.A2(n_1262),
.A3(n_1283),
.B(n_1161),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1216),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1148),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1284),
.A2(n_1196),
.B(n_1166),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1245),
.A2(n_1283),
.B(n_1281),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1199),
.B(n_1204),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1208),
.B(n_1159),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1146),
.A2(n_1172),
.B(n_1263),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1277),
.A2(n_1174),
.B(n_1280),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1279),
.A2(n_1143),
.B(n_1165),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1183),
.A2(n_1211),
.B(n_1222),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1230),
.B(n_1143),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1243),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1212),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1155),
.A2(n_1141),
.B(n_1160),
.Y(n_1323)
);

INVx6_ASAP7_75t_SL g1324 ( 
.A(n_1240),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1242),
.B(n_1189),
.Y(n_1325)
);

NOR2x1_ASAP7_75t_L g1326 ( 
.A(n_1206),
.B(n_1251),
.Y(n_1326)
);

AOI221xp5_ASAP7_75t_L g1327 ( 
.A1(n_1162),
.A2(n_1163),
.B1(n_1139),
.B2(n_1147),
.C(n_1161),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1230),
.B(n_1229),
.Y(n_1328)
);

CKINVDCx6p67_ASAP7_75t_R g1329 ( 
.A(n_1240),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1249),
.Y(n_1330)
);

O2A1O1Ixp33_ASAP7_75t_SL g1331 ( 
.A1(n_1178),
.A2(n_1158),
.B(n_1171),
.C(n_1135),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1137),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1246),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1153),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1232),
.A2(n_1244),
.B(n_1247),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1266),
.A2(n_1154),
.A3(n_1272),
.B(n_1286),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1140),
.B(n_1173),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1272),
.A2(n_1266),
.B(n_1136),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_SL g1339 ( 
.A1(n_1158),
.A2(n_1171),
.B(n_1136),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1144),
.A2(n_1132),
.B(n_1169),
.Y(n_1340)
);

AOI31xp67_ASAP7_75t_L g1341 ( 
.A1(n_1268),
.A2(n_1145),
.A3(n_1225),
.B(n_1223),
.Y(n_1341)
);

AOI221x1_ASAP7_75t_L g1342 ( 
.A1(n_1217),
.A2(n_1238),
.B1(n_1231),
.B2(n_1195),
.C(n_1241),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1288),
.A2(n_1234),
.A3(n_1225),
.B(n_1223),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1135),
.A2(n_1228),
.B(n_1264),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1132),
.A2(n_1169),
.B(n_1285),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1236),
.B(n_1260),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1179),
.A2(n_1278),
.B(n_1276),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1238),
.A2(n_1217),
.A3(n_1167),
.B(n_1287),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1216),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1157),
.A2(n_1287),
.B(n_1219),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1216),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1210),
.A2(n_1188),
.B(n_1213),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1168),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1270),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1260),
.B(n_1265),
.Y(n_1355)
);

AOI221xp5_ASAP7_75t_L g1356 ( 
.A1(n_1202),
.A2(n_1177),
.B1(n_1226),
.B2(n_1205),
.C(n_1197),
.Y(n_1356)
);

AOI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1237),
.A2(n_1192),
.B1(n_1194),
.B2(n_1227),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1176),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1269),
.A2(n_1263),
.B(n_1265),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1269),
.A2(n_1273),
.B(n_1252),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1167),
.A2(n_1233),
.A3(n_1201),
.B(n_1198),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1207),
.B(n_1213),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1240),
.A2(n_1186),
.B1(n_1187),
.B2(n_1191),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1193),
.A2(n_1235),
.B(n_1233),
.C(n_1142),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1252),
.A2(n_1256),
.B(n_1215),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1187),
.A2(n_1191),
.B1(n_1210),
.B2(n_1188),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1188),
.A2(n_1275),
.B1(n_1180),
.B2(n_1214),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1203),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1190),
.A2(n_1152),
.B(n_1149),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1164),
.A2(n_1282),
.B(n_1221),
.Y(n_1370)
);

AO31x2_ASAP7_75t_L g1371 ( 
.A1(n_1274),
.A2(n_1251),
.A3(n_1206),
.B(n_1248),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1134),
.A2(n_1138),
.B(n_1214),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1246),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1258),
.B(n_1149),
.Y(n_1374)
);

AOI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1152),
.A2(n_1253),
.B(n_1221),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1156),
.A2(n_1134),
.B1(n_1253),
.B2(n_1274),
.Y(n_1376)
);

AO31x2_ASAP7_75t_L g1377 ( 
.A1(n_1274),
.A2(n_1150),
.A3(n_947),
.B(n_982),
.Y(n_1377)
);

BUFx3_ASAP7_75t_L g1378 ( 
.A(n_1253),
.Y(n_1378)
);

AOI221x1_ASAP7_75t_L g1379 ( 
.A1(n_1134),
.A2(n_1150),
.B1(n_1244),
.B2(n_1232),
.C(n_984),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1134),
.B(n_1036),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1208),
.B(n_867),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1209),
.B(n_1224),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1162),
.B(n_1018),
.Y(n_1383)
);

O2A1O1Ixp33_ASAP7_75t_SL g1384 ( 
.A1(n_1150),
.A2(n_1218),
.B(n_1220),
.C(n_1178),
.Y(n_1384)
);

AOI211x1_ASAP7_75t_L g1385 ( 
.A1(n_1189),
.A2(n_1217),
.B(n_1238),
.C(n_1139),
.Y(n_1385)
);

O2A1O1Ixp5_ASAP7_75t_L g1386 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1218),
.C(n_1150),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1388)
);

A2O1A1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1150),
.C(n_804),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1208),
.B(n_867),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1208),
.B(n_1018),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1393)
);

INVx5_ASAP7_75t_L g1394 ( 
.A(n_1216),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1137),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1232),
.A2(n_1244),
.B(n_1171),
.Y(n_1397)
);

BUFx4_ASAP7_75t_SL g1398 ( 
.A(n_1170),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1150),
.A2(n_947),
.A3(n_982),
.B(n_1261),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1400)
);

AO31x2_ASAP7_75t_L g1401 ( 
.A1(n_1150),
.A2(n_947),
.A3(n_982),
.B(n_1261),
.Y(n_1401)
);

AO32x2_ASAP7_75t_L g1402 ( 
.A1(n_1161),
.A2(n_1238),
.A3(n_1217),
.B1(n_1266),
.B2(n_1281),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1162),
.A2(n_1036),
.B1(n_1163),
.B2(n_991),
.Y(n_1403)
);

BUFx8_ASAP7_75t_L g1404 ( 
.A(n_1212),
.Y(n_1404)
);

INVx5_ASAP7_75t_L g1405 ( 
.A(n_1216),
.Y(n_1405)
);

BUFx12f_ASAP7_75t_L g1406 ( 
.A(n_1200),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1407)
);

BUFx12f_ASAP7_75t_L g1408 ( 
.A(n_1200),
.Y(n_1408)
);

AOI221x1_ASAP7_75t_L g1409 ( 
.A1(n_1150),
.A2(n_1244),
.B1(n_1232),
.B2(n_984),
.C(n_991),
.Y(n_1409)
);

INVx3_ASAP7_75t_L g1410 ( 
.A(n_1132),
.Y(n_1410)
);

AOI221x1_ASAP7_75t_L g1411 ( 
.A1(n_1150),
.A2(n_1244),
.B1(n_1232),
.B2(n_984),
.C(n_991),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1208),
.B(n_1036),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_SL g1413 ( 
.A(n_1242),
.B(n_1036),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1209),
.B(n_1224),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1415)
);

CKINVDCx11_ASAP7_75t_R g1416 ( 
.A(n_1181),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1162),
.A2(n_1036),
.B1(n_1163),
.B2(n_1195),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1250),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1209),
.B(n_1224),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1423)
);

NOR2xp67_ASAP7_75t_L g1424 ( 
.A(n_1200),
.B(n_892),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1150),
.A2(n_1218),
.B(n_1245),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1150),
.A2(n_1218),
.B(n_1245),
.Y(n_1426)
);

AO31x2_ASAP7_75t_L g1427 ( 
.A1(n_1150),
.A2(n_947),
.A3(n_982),
.B(n_1261),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1185),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1162),
.B(n_1018),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1162),
.A2(n_1163),
.B(n_1150),
.C(n_804),
.Y(n_1431)
);

NAND3x1_ASAP7_75t_L g1432 ( 
.A(n_1162),
.B(n_712),
.C(n_904),
.Y(n_1432)
);

AO221x2_ASAP7_75t_L g1433 ( 
.A1(n_1217),
.A2(n_1238),
.B1(n_1226),
.B2(n_1161),
.C(n_1198),
.Y(n_1433)
);

XOR2xp5_ASAP7_75t_L g1434 ( 
.A(n_1200),
.B(n_605),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1170),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1150),
.A2(n_1036),
.B1(n_1242),
.B2(n_973),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1162),
.A2(n_904),
.B1(n_1163),
.B2(n_843),
.C(n_944),
.Y(n_1437)
);

NAND3x1_ASAP7_75t_L g1438 ( 
.A(n_1162),
.B(n_712),
.C(n_904),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1209),
.B(n_1224),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_SL g1440 ( 
.A1(n_1150),
.A2(n_1218),
.B(n_1220),
.C(n_1178),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1218),
.A2(n_1261),
.B(n_1175),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1216),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1218),
.A2(n_1261),
.B(n_1175),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1218),
.A2(n_985),
.B(n_986),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1137),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1150),
.A2(n_1036),
.B1(n_1242),
.B2(n_973),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1448)
);

AOI221x1_ASAP7_75t_L g1449 ( 
.A1(n_1150),
.A2(n_1244),
.B1(n_1232),
.B2(n_984),
.C(n_991),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1208),
.B(n_1036),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1254),
.A2(n_1040),
.B(n_1175),
.Y(n_1451)
);

BUFx8_ASAP7_75t_L g1452 ( 
.A(n_1212),
.Y(n_1452)
);

OA21x2_ASAP7_75t_L g1453 ( 
.A1(n_1218),
.A2(n_1261),
.B(n_1175),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1200),
.B(n_892),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1162),
.B(n_1018),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1437),
.A2(n_1418),
.B1(n_1403),
.B2(n_1433),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1418),
.A2(n_1433),
.B1(n_1327),
.B2(n_1356),
.Y(n_1457)
);

BUFx4f_ASAP7_75t_L g1458 ( 
.A(n_1292),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1436),
.A2(n_1446),
.B1(n_1413),
.B2(n_1455),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1389),
.A2(n_1431),
.B1(n_1366),
.B2(n_1432),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1438),
.A2(n_1429),
.B1(n_1383),
.B2(n_1363),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1332),
.Y(n_1462)
);

BUFx12f_ASAP7_75t_L g1463 ( 
.A(n_1416),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1328),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1334),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1410),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1353),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1311),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1301),
.Y(n_1469)
);

OAI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1413),
.A2(n_1325),
.B1(n_1446),
.B2(n_1436),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1358),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1435),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1371),
.Y(n_1473)
);

OAI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1325),
.A2(n_1357),
.B1(n_1342),
.B2(n_1439),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1335),
.A2(n_1357),
.B1(n_1365),
.B2(n_1367),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1306),
.B(n_1314),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1395),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1410),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1310),
.B(n_1394),
.Y(n_1479)
);

INVx1_ASAP7_75t_SL g1480 ( 
.A(n_1315),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1306),
.A2(n_1439),
.B1(n_1414),
.B2(n_1422),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1367),
.A2(n_1335),
.B1(n_1363),
.B2(n_1380),
.Y(n_1482)
);

NAND2x1p5_ASAP7_75t_L g1483 ( 
.A(n_1394),
.B(n_1405),
.Y(n_1483)
);

BUFx12f_ASAP7_75t_L g1484 ( 
.A(n_1322),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1425),
.A2(n_1426),
.B1(n_1412),
.B2(n_1450),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1428),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1294),
.B(n_1296),
.Y(n_1487)
);

NAND2x1p5_ASAP7_75t_L g1488 ( 
.A(n_1405),
.B(n_1378),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1352),
.A2(n_1422),
.B1(n_1382),
.B2(n_1314),
.Y(n_1489)
);

INVx6_ASAP7_75t_L g1490 ( 
.A(n_1404),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1406),
.Y(n_1491)
);

OAI22x1_ASAP7_75t_L g1492 ( 
.A1(n_1376),
.A2(n_1320),
.B1(n_1391),
.B2(n_1382),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1424),
.A2(n_1454),
.B1(n_1362),
.B2(n_1434),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1445),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1408),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1330),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1404),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1414),
.A2(n_1329),
.B1(n_1320),
.B2(n_1324),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1354),
.Y(n_1499)
);

BUFx10_ASAP7_75t_L g1500 ( 
.A(n_1368),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1295),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1304),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1452),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1297),
.A2(n_1303),
.B1(n_1319),
.B2(n_1360),
.Y(n_1504)
);

CKINVDCx16_ASAP7_75t_R g1505 ( 
.A(n_1302),
.Y(n_1505)
);

BUFx4_ASAP7_75t_R g1506 ( 
.A(n_1333),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1326),
.B(n_1375),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1452),
.Y(n_1508)
);

INVx4_ASAP7_75t_L g1509 ( 
.A(n_1349),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1425),
.A2(n_1426),
.B1(n_1420),
.B2(n_1324),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_SL g1511 ( 
.A1(n_1319),
.A2(n_1372),
.B1(n_1386),
.B2(n_1373),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1313),
.A2(n_1453),
.B1(n_1443),
.B2(n_1441),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1313),
.A2(n_1453),
.B1(n_1443),
.B2(n_1441),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1362),
.A2(n_1337),
.B1(n_1307),
.B2(n_1390),
.Y(n_1514)
);

BUFx8_ASAP7_75t_SL g1515 ( 
.A(n_1307),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1347),
.A2(n_1346),
.B1(n_1385),
.B2(n_1323),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1337),
.B(n_1381),
.Y(n_1517)
);

AOI22xp5_ASAP7_75t_L g1518 ( 
.A1(n_1372),
.A2(n_1298),
.B1(n_1384),
.B2(n_1440),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1349),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1398),
.Y(n_1520)
);

INVx6_ASAP7_75t_L g1521 ( 
.A(n_1351),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1351),
.Y(n_1522)
);

CKINVDCx20_ASAP7_75t_R g1523 ( 
.A(n_1442),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1347),
.A2(n_1346),
.B1(n_1397),
.B2(n_1344),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1374),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1350),
.A2(n_1339),
.B1(n_1364),
.B2(n_1411),
.Y(n_1526)
);

CKINVDCx11_ASAP7_75t_R g1527 ( 
.A(n_1442),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1344),
.A2(n_1350),
.B1(n_1316),
.B2(n_1293),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1370),
.Y(n_1529)
);

BUFx12f_ASAP7_75t_L g1530 ( 
.A(n_1442),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1374),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1316),
.A2(n_1387),
.B1(n_1393),
.B2(n_1444),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1392),
.A2(n_1396),
.B1(n_1400),
.B2(n_1421),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1355),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1355),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_SL g1536 ( 
.A1(n_1409),
.A2(n_1449),
.B1(n_1402),
.B2(n_1419),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1379),
.A2(n_1402),
.B1(n_1415),
.B2(n_1430),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1338),
.A2(n_1402),
.B1(n_1318),
.B2(n_1359),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1369),
.A2(n_1345),
.B1(n_1340),
.B2(n_1308),
.Y(n_1539)
);

CKINVDCx11_ASAP7_75t_R g1540 ( 
.A(n_1341),
.Y(n_1540)
);

INVx11_ASAP7_75t_L g1541 ( 
.A(n_1371),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1317),
.A2(n_1348),
.B1(n_1361),
.B2(n_1417),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1371),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_SL g1544 ( 
.A1(n_1348),
.A2(n_1361),
.B1(n_1312),
.B2(n_1299),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1343),
.B(n_1361),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1343),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1348),
.A2(n_1388),
.B1(n_1448),
.B2(n_1447),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_SL g1548 ( 
.A1(n_1407),
.A2(n_1451),
.B1(n_1423),
.B2(n_1309),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1343),
.Y(n_1549)
);

BUFx12f_ASAP7_75t_L g1550 ( 
.A(n_1331),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1291),
.A2(n_1290),
.B1(n_1300),
.B2(n_1336),
.Y(n_1551)
);

OAI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1399),
.A2(n_1401),
.B1(n_1427),
.B2(n_1309),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1336),
.B(n_1305),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1309),
.A2(n_1399),
.B1(n_1401),
.B2(n_1427),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1399),
.A2(n_1401),
.B1(n_1427),
.B2(n_1377),
.Y(n_1555)
);

BUFx10_ASAP7_75t_L g1556 ( 
.A(n_1305),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1377),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1305),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1437),
.A2(n_1036),
.B1(n_1418),
.B2(n_1403),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1332),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1321),
.Y(n_1561)
);

INVx5_ASAP7_75t_L g1562 ( 
.A(n_1310),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1437),
.A2(n_1036),
.B1(n_1418),
.B2(n_1403),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1310),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1321),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_SL g1566 ( 
.A(n_1404),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1437),
.B2(n_1431),
.Y(n_1567)
);

BUFx4f_ASAP7_75t_SL g1568 ( 
.A(n_1292),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1311),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1321),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1437),
.A2(n_1036),
.B1(n_1418),
.B2(n_1403),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1383),
.B(n_1429),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1418),
.A2(n_1413),
.B1(n_1437),
.B2(n_1325),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1416),
.Y(n_1574)
);

INVx6_ASAP7_75t_L g1575 ( 
.A(n_1404),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1413),
.A2(n_1036),
.B1(n_1163),
.B2(n_1162),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1404),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1412),
.B(n_1450),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1321),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1371),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1437),
.A2(n_1036),
.B1(n_1418),
.B2(n_1403),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1321),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1437),
.A2(n_1036),
.B1(n_1418),
.B2(n_1403),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1383),
.B(n_1429),
.Y(n_1584)
);

BUFx12f_ASAP7_75t_L g1585 ( 
.A(n_1416),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1428),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_R g1587 ( 
.A1(n_1383),
.A2(n_244),
.B1(n_300),
.B2(n_215),
.Y(n_1587)
);

BUFx2_ASAP7_75t_SL g1588 ( 
.A(n_1424),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_SL g1589 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1036),
.B2(n_1383),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1437),
.B2(n_1431),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1437),
.B2(n_1431),
.Y(n_1591)
);

CKINVDCx11_ASAP7_75t_R g1592 ( 
.A(n_1416),
.Y(n_1592)
);

BUFx12f_ASAP7_75t_L g1593 ( 
.A(n_1416),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_SL g1594 ( 
.A1(n_1413),
.A2(n_1036),
.B1(n_1163),
.B2(n_1162),
.Y(n_1594)
);

AOI22xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1413),
.A2(n_1036),
.B1(n_1163),
.B2(n_1162),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_SL g1596 ( 
.A(n_1404),
.Y(n_1596)
);

CKINVDCx11_ASAP7_75t_R g1597 ( 
.A(n_1416),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1289),
.Y(n_1598)
);

CKINVDCx16_ASAP7_75t_R g1599 ( 
.A(n_1292),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1310),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1413),
.A2(n_1036),
.B1(n_1163),
.B2(n_1162),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1389),
.A2(n_1431),
.B(n_1335),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1332),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1413),
.A2(n_1036),
.B1(n_1163),
.B2(n_1162),
.Y(n_1604)
);

OAI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1418),
.A2(n_1413),
.B1(n_1437),
.B2(n_1325),
.Y(n_1605)
);

BUFx8_ASAP7_75t_SL g1606 ( 
.A(n_1292),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1437),
.B2(n_1431),
.Y(n_1607)
);

BUFx2_ASAP7_75t_L g1608 ( 
.A(n_1311),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1332),
.Y(n_1609)
);

CKINVDCx11_ASAP7_75t_R g1610 ( 
.A(n_1416),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1332),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1437),
.B2(n_1431),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1546),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1539),
.A2(n_1547),
.B(n_1533),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1549),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1485),
.B(n_1475),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1462),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1520),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1547),
.A2(n_1533),
.B(n_1532),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1589),
.A2(n_1612),
.B1(n_1607),
.B2(n_1567),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1532),
.A2(n_1551),
.B(n_1542),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1471),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1542),
.A2(n_1553),
.B(n_1529),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1545),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1559),
.A2(n_1583),
.B1(n_1563),
.B2(n_1581),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1512),
.A2(n_1513),
.B(n_1602),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1557),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1559),
.A2(n_1583),
.B1(n_1563),
.B2(n_1571),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1473),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1576),
.A2(n_1595),
.B1(n_1594),
.B2(n_1601),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1512),
.A2(n_1513),
.B(n_1538),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1473),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1477),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1538),
.A2(n_1524),
.B(n_1528),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1543),
.Y(n_1636)
);

CKINVDCx14_ASAP7_75t_R g1637 ( 
.A(n_1592),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1485),
.B(n_1475),
.Y(n_1638)
);

OA21x2_ASAP7_75t_L g1639 ( 
.A1(n_1524),
.A2(n_1528),
.B(n_1554),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1580),
.Y(n_1640)
);

AOI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1590),
.A2(n_1591),
.B(n_1460),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1580),
.Y(n_1642)
);

INVx3_ASAP7_75t_SL g1643 ( 
.A(n_1562),
.Y(n_1643)
);

AOI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1481),
.A2(n_1476),
.B(n_1537),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1494),
.B(n_1560),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1525),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1554),
.B(n_1555),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1558),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1562),
.Y(n_1649)
);

OA21x2_ASAP7_75t_L g1650 ( 
.A1(n_1555),
.A2(n_1516),
.B(n_1510),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1541),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1537),
.A2(n_1552),
.B(n_1481),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1468),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1597),
.Y(n_1654)
);

INVx3_ASAP7_75t_L g1655 ( 
.A(n_1556),
.Y(n_1655)
);

BUFx2_ASAP7_75t_R g1656 ( 
.A(n_1606),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1464),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1553),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1486),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1603),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_L g1661 ( 
.A1(n_1571),
.A2(n_1581),
.B1(n_1604),
.B2(n_1456),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1507),
.A2(n_1516),
.B(n_1518),
.Y(n_1662)
);

NAND2x1p5_ASAP7_75t_L g1663 ( 
.A(n_1562),
.B(n_1534),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1609),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1492),
.Y(n_1665)
);

BUFx2_ASAP7_75t_L g1666 ( 
.A(n_1550),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1578),
.B(n_1482),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1611),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1507),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_SL g1670 ( 
.A1(n_1461),
.A2(n_1535),
.B1(n_1573),
.B2(n_1605),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1544),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1496),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1510),
.A2(n_1457),
.B(n_1456),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1499),
.Y(n_1674)
);

OAI21x1_ASAP7_75t_L g1675 ( 
.A1(n_1489),
.A2(n_1570),
.B(n_1561),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1531),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1565),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1487),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1579),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1457),
.B(n_1536),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1582),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1608),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1466),
.A2(n_1478),
.B(n_1502),
.Y(n_1683)
);

OAI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1466),
.A2(n_1478),
.B(n_1488),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1526),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1488),
.A2(n_1548),
.B(n_1479),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1540),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1474),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1572),
.B(n_1584),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1515),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1474),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1498),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1498),
.Y(n_1693)
);

CKINVDCx20_ASAP7_75t_R g1694 ( 
.A(n_1610),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1511),
.Y(n_1695)
);

OAI21x1_ASAP7_75t_L g1696 ( 
.A1(n_1479),
.A2(n_1483),
.B(n_1514),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1573),
.A2(n_1605),
.B(n_1504),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_SL g1698 ( 
.A1(n_1587),
.A2(n_1470),
.B1(n_1490),
.B2(n_1575),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1483),
.Y(n_1699)
);

OR2x6_ASAP7_75t_L g1700 ( 
.A(n_1490),
.B(n_1575),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1519),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1459),
.A2(n_1470),
.B(n_1493),
.Y(n_1702)
);

BUFx3_ASAP7_75t_L g1703 ( 
.A(n_1523),
.Y(n_1703)
);

NAND2x1p5_ASAP7_75t_L g1704 ( 
.A(n_1564),
.B(n_1600),
.Y(n_1704)
);

CKINVDCx20_ASAP7_75t_R g1705 ( 
.A(n_1469),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1459),
.A2(n_1586),
.B(n_1569),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1501),
.B(n_1472),
.Y(n_1708)
);

OAI21x1_ASAP7_75t_L g1709 ( 
.A1(n_1564),
.A2(n_1600),
.B(n_1521),
.Y(n_1709)
);

INVx2_ASAP7_75t_SL g1710 ( 
.A(n_1598),
.Y(n_1710)
);

CKINVDCx20_ASAP7_75t_R g1711 ( 
.A(n_1568),
.Y(n_1711)
);

INVx4_ASAP7_75t_SL g1712 ( 
.A(n_1490),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1598),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1509),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1509),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1530),
.Y(n_1716)
);

OAI21x1_ASAP7_75t_SL g1717 ( 
.A1(n_1522),
.A2(n_1506),
.B(n_1596),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1588),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_1527),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1577),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1500),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1566),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1505),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1577),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1508),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1497),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1620),
.A2(n_1631),
.B1(n_1697),
.B2(n_1661),
.Y(n_1727)
);

CKINVDCx5p33_ASAP7_75t_R g1728 ( 
.A(n_1618),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1651),
.B(n_1497),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_SL g1730 ( 
.A(n_1652),
.B(n_1463),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1706),
.B(n_1503),
.Y(n_1731)
);

AO22x1_ASAP7_75t_SL g1732 ( 
.A1(n_1687),
.A2(n_1593),
.B1(n_1585),
.B2(n_1484),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1623),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1700),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1706),
.B(n_1503),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1657),
.B(n_1599),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1630),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1651),
.B(n_1491),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1678),
.B(n_1458),
.Y(n_1739)
);

BUFx3_ASAP7_75t_L g1740 ( 
.A(n_1717),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1622),
.A2(n_1495),
.B(n_1574),
.Y(n_1741)
);

AO32x1_ASAP7_75t_L g1742 ( 
.A1(n_1680),
.A2(n_1458),
.A3(n_1500),
.B1(n_1568),
.B2(n_1688),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1662),
.B(n_1644),
.Y(n_1743)
);

O2A1O1Ixp33_ASAP7_75t_L g1744 ( 
.A1(n_1702),
.A2(n_1685),
.B(n_1695),
.C(n_1626),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1652),
.A2(n_1614),
.B(n_1635),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1653),
.Y(n_1746)
);

AO32x2_ASAP7_75t_L g1747 ( 
.A1(n_1710),
.A2(n_1649),
.A3(n_1636),
.B1(n_1652),
.B2(n_1640),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1641),
.B(n_1695),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1719),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1621),
.B(n_1645),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1662),
.B(n_1663),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1619),
.A2(n_1622),
.B(n_1614),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1634),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1629),
.A2(n_1670),
.B1(n_1698),
.B2(n_1673),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1673),
.A2(n_1689),
.B1(n_1685),
.B2(n_1641),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1700),
.A2(n_1673),
.B(n_1663),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1667),
.B(n_1665),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1646),
.B(n_1676),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1616),
.A2(n_1638),
.B1(n_1691),
.B2(n_1688),
.C(n_1680),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1713),
.B(n_1687),
.Y(n_1760)
);

OAI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1616),
.A2(n_1638),
.B(n_1692),
.Y(n_1761)
);

AOI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1707),
.A2(n_1693),
.B1(n_1671),
.B2(n_1659),
.C(n_1682),
.Y(n_1762)
);

O2A1O1Ixp33_ASAP7_75t_SL g1763 ( 
.A1(n_1718),
.A2(n_1720),
.B(n_1721),
.C(n_1710),
.Y(n_1763)
);

BUFx4f_ASAP7_75t_SL g1764 ( 
.A(n_1694),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1621),
.B(n_1645),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1618),
.Y(n_1766)
);

NOR2x1p5_ASAP7_75t_L g1767 ( 
.A(n_1690),
.B(n_1719),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1675),
.A2(n_1619),
.B(n_1673),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1675),
.A2(n_1718),
.B(n_1696),
.Y(n_1769)
);

NAND3xp33_ASAP7_75t_L g1770 ( 
.A(n_1708),
.B(n_1676),
.C(n_1679),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1686),
.A2(n_1624),
.B(n_1683),
.Y(n_1771)
);

AO32x2_ASAP7_75t_L g1772 ( 
.A1(n_1649),
.A2(n_1636),
.A3(n_1630),
.B1(n_1633),
.B2(n_1640),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1669),
.B(n_1660),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1635),
.A2(n_1627),
.B(n_1639),
.Y(n_1774)
);

INVx2_ASAP7_75t_SL g1775 ( 
.A(n_1719),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1682),
.B(n_1708),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1696),
.A2(n_1663),
.B(n_1684),
.Y(n_1777)
);

AO32x2_ASAP7_75t_L g1778 ( 
.A1(n_1633),
.A2(n_1642),
.A3(n_1647),
.B1(n_1625),
.B2(n_1639),
.Y(n_1778)
);

AND2x6_ASAP7_75t_L g1779 ( 
.A(n_1669),
.B(n_1658),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_SL g1780 ( 
.A1(n_1719),
.A2(n_1690),
.B(n_1720),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1677),
.B(n_1679),
.C(n_1681),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_L g1782 ( 
.A1(n_1723),
.A2(n_1726),
.B1(n_1725),
.B2(n_1724),
.C(n_1666),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_SL g1783 ( 
.A(n_1628),
.B(n_1648),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1719),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1726),
.A2(n_1716),
.B1(n_1722),
.B2(n_1703),
.Y(n_1785)
);

O2A1O1Ixp33_ASAP7_75t_L g1786 ( 
.A1(n_1717),
.A2(n_1669),
.B(n_1674),
.C(n_1672),
.Y(n_1786)
);

INVx4_ASAP7_75t_L g1787 ( 
.A(n_1712),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1650),
.A2(n_1635),
.B1(n_1639),
.B2(n_1637),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1617),
.Y(n_1789)
);

NOR2x1_ASAP7_75t_L g1790 ( 
.A(n_1714),
.B(n_1715),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1664),
.B(n_1668),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1716),
.A2(n_1701),
.B1(n_1703),
.B2(n_1650),
.Y(n_1792)
);

OAI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1684),
.A2(n_1709),
.B(n_1699),
.Y(n_1793)
);

OA21x2_ASAP7_75t_L g1794 ( 
.A1(n_1624),
.A2(n_1613),
.B(n_1615),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1747),
.Y(n_1795)
);

NOR2x1_ASAP7_75t_L g1796 ( 
.A(n_1790),
.B(n_1655),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1737),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1794),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1752),
.B(n_1632),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1747),
.B(n_1632),
.Y(n_1800)
);

INVx1_ASAP7_75t_SL g1801 ( 
.A(n_1736),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1794),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1747),
.B(n_1768),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1747),
.B(n_1632),
.Y(n_1804)
);

INVxp67_ASAP7_75t_SL g1805 ( 
.A(n_1781),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1778),
.B(n_1627),
.Y(n_1806)
);

HB1xp67_ASAP7_75t_L g1807 ( 
.A(n_1733),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1753),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1778),
.B(n_1627),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1778),
.B(n_1635),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1743),
.B(n_1639),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1771),
.B(n_1773),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1751),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1774),
.B(n_1615),
.Y(n_1814)
);

BUFx5_ASAP7_75t_L g1815 ( 
.A(n_1779),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1774),
.B(n_1650),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1745),
.B(n_1650),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1789),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1751),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1772),
.Y(n_1821)
);

INVx5_ASAP7_75t_L g1822 ( 
.A(n_1751),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1808),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1805),
.B(n_1791),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1825)
);

NAND4xp25_ASAP7_75t_L g1826 ( 
.A(n_1817),
.B(n_1727),
.C(n_1744),
.D(n_1754),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1802),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1802),
.Y(n_1828)
);

OAI221xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1805),
.A2(n_1744),
.B1(n_1759),
.B2(n_1762),
.C(n_1788),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1812),
.B(n_1777),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1800),
.B(n_1741),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1804),
.B(n_1788),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1802),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1820),
.B(n_1748),
.Y(n_1835)
);

AOI221xp5_ASAP7_75t_L g1836 ( 
.A1(n_1817),
.A2(n_1755),
.B1(n_1759),
.B2(n_1748),
.C(n_1762),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1814),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1814),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1814),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1820),
.B(n_1770),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1798),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1798),
.Y(n_1842)
);

INVx3_ASAP7_75t_L g1843 ( 
.A(n_1812),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1804),
.B(n_1772),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1812),
.B(n_1793),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1812),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1801),
.A2(n_1761),
.B1(n_1792),
.B2(n_1776),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1821),
.B(n_1783),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1806),
.B(n_1772),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_SL g1850 ( 
.A(n_1822),
.B(n_1787),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1801),
.A2(n_1776),
.B1(n_1757),
.B2(n_1746),
.Y(n_1851)
);

NOR2x1_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_1756),
.Y(n_1852)
);

AOI211xp5_ASAP7_75t_L g1853 ( 
.A1(n_1817),
.A2(n_1780),
.B(n_1782),
.C(n_1786),
.Y(n_1853)
);

AOI221xp5_ASAP7_75t_L g1854 ( 
.A1(n_1803),
.A2(n_1758),
.B1(n_1786),
.B2(n_1785),
.C(n_1769),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1813),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1816),
.A2(n_1742),
.B(n_1730),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1796),
.B(n_1734),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1806),
.B(n_1750),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1813),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1807),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1807),
.Y(n_1861)
);

INVx4_ASAP7_75t_L g1862 ( 
.A(n_1815),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1812),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1809),
.B(n_1765),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1827),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1823),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1837),
.B(n_1803),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1849),
.B(n_1803),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1849),
.B(n_1844),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1837),
.B(n_1795),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1851),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1837),
.B(n_1795),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1835),
.B(n_1797),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1827),
.Y(n_1874)
);

BUFx3_ASAP7_75t_L g1875 ( 
.A(n_1855),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1862),
.B(n_1822),
.Y(n_1876)
);

BUFx2_ASAP7_75t_L g1877 ( 
.A(n_1852),
.Y(n_1877)
);

NOR2x1_ASAP7_75t_L g1878 ( 
.A(n_1852),
.B(n_1767),
.Y(n_1878)
);

INVxp67_ASAP7_75t_SL g1879 ( 
.A(n_1841),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1849),
.B(n_1811),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1837),
.B(n_1797),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1827),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1827),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1860),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1849),
.B(n_1811),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1844),
.B(n_1811),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1844),
.B(n_1810),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1838),
.B(n_1809),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1838),
.B(n_1839),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1860),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1835),
.B(n_1810),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1857),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1828),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1828),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1839),
.B(n_1816),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1839),
.B(n_1816),
.Y(n_1897)
);

OAI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1826),
.A2(n_1763),
.B(n_1799),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1857),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1861),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1828),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1834),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1835),
.B(n_1818),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1861),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1884),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1873),
.B(n_1840),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1873),
.B(n_1840),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1903),
.B(n_1840),
.Y(n_1908)
);

HB1xp67_ASAP7_75t_L g1909 ( 
.A(n_1875),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1903),
.B(n_1824),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1871),
.B(n_1824),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1884),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1891),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1890),
.Y(n_1914)
);

AND2x4_ASAP7_75t_L g1915 ( 
.A(n_1878),
.B(n_1852),
.Y(n_1915)
);

BUFx3_ASAP7_75t_L g1916 ( 
.A(n_1875),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1891),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1869),
.B(n_1855),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1890),
.Y(n_1919)
);

INVx1_ASAP7_75t_SL g1920 ( 
.A(n_1878),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1871),
.A2(n_1826),
.B1(n_1836),
.B2(n_1854),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1869),
.B(n_1855),
.Y(n_1922)
);

AOI211xp5_ASAP7_75t_L g1923 ( 
.A1(n_1898),
.A2(n_1826),
.B(n_1829),
.C(n_1836),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1875),
.B(n_1862),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1893),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.B(n_1824),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1875),
.B(n_1862),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1900),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_L g1929 ( 
.A(n_1898),
.B(n_1846),
.Y(n_1929)
);

INVxp67_ASAP7_75t_L g1930 ( 
.A(n_1877),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1869),
.B(n_1859),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1868),
.B(n_1859),
.Y(n_1932)
);

OAI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1877),
.A2(n_1854),
.B(n_1853),
.C(n_1847),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1900),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1876),
.B(n_1862),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1904),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1867),
.B(n_1848),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1890),
.Y(n_1938)
);

AOI32xp33_ASAP7_75t_L g1939 ( 
.A1(n_1877),
.A2(n_1833),
.A3(n_1853),
.B1(n_1847),
.B2(n_1825),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1904),
.Y(n_1940)
);

NAND2x1p5_ASAP7_75t_L g1941 ( 
.A(n_1893),
.B(n_1822),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1867),
.B(n_1848),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1899),
.B(n_1851),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1892),
.B(n_1848),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1868),
.B(n_1859),
.Y(n_1945)
);

INVx1_ASAP7_75t_SL g1946 ( 
.A(n_1899),
.Y(n_1946)
);

AOI21xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1876),
.A2(n_1654),
.B(n_1728),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1866),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1866),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1870),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1881),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1911),
.B(n_1892),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1923),
.B(n_1833),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1928),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1928),
.Y(n_1955)
);

OAI31xp33_ASAP7_75t_SL g1956 ( 
.A1(n_1933),
.A2(n_1868),
.A3(n_1833),
.B(n_1876),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1936),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1936),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1915),
.B(n_1876),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1921),
.B(n_1833),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1905),
.Y(n_1961)
);

INVx2_ASAP7_75t_SL g1962 ( 
.A(n_1916),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1920),
.Y(n_1963)
);

INVx1_ASAP7_75t_SL g1964 ( 
.A(n_1925),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1943),
.B(n_1880),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1912),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1913),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1939),
.B(n_1864),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1946),
.B(n_1880),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1918),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1915),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1916),
.Y(n_1972)
);

NOR2xp67_ASAP7_75t_SL g1973 ( 
.A(n_1909),
.B(n_1654),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1910),
.B(n_1880),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1917),
.B(n_1864),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1915),
.B(n_1929),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1918),
.B(n_1885),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1934),
.B(n_1864),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1940),
.B(n_1864),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1922),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1949),
.Y(n_1981)
);

OR2x2_ASAP7_75t_L g1982 ( 
.A(n_1910),
.B(n_1885),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1932),
.B(n_1858),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1947),
.B(n_1764),
.Y(n_1984)
);

NAND2x1p5_ASAP7_75t_L g1985 ( 
.A(n_1935),
.B(n_1784),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1949),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1932),
.B(n_1858),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1926),
.B(n_1885),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1908),
.B(n_1764),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1948),
.Y(n_1990)
);

AOI21xp33_ASAP7_75t_L g1991 ( 
.A1(n_1956),
.A2(n_1930),
.B(n_1927),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1960),
.A2(n_1829),
.B(n_1853),
.Y(n_1992)
);

O2A1O1Ixp33_ASAP7_75t_L g1993 ( 
.A1(n_1953),
.A2(n_1941),
.B(n_1906),
.C(n_1907),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1968),
.A2(n_1964),
.B1(n_1976),
.B2(n_1963),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1989),
.B(n_1656),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1959),
.Y(n_1996)
);

INVxp67_ASAP7_75t_L g1997 ( 
.A(n_1989),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1976),
.A2(n_1941),
.B(n_1766),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1976),
.A2(n_1941),
.B(n_1856),
.Y(n_1999)
);

AND2x2_ASAP7_75t_SL g2000 ( 
.A(n_1984),
.B(n_1784),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1962),
.B(n_1945),
.Y(n_2001)
);

OAI21x1_ASAP7_75t_L g2002 ( 
.A1(n_1985),
.A2(n_1919),
.B(n_1914),
.Y(n_2002)
);

NAND2x1p5_ASAP7_75t_L g2003 ( 
.A(n_1973),
.B(n_1784),
.Y(n_2003)
);

INVxp67_ASAP7_75t_L g2004 ( 
.A(n_1962),
.Y(n_2004)
);

OAI221xp5_ASAP7_75t_SL g2005 ( 
.A1(n_1971),
.A2(n_1856),
.B1(n_1926),
.B2(n_1937),
.C(n_1942),
.Y(n_2005)
);

OAI21xp33_ASAP7_75t_SL g2006 ( 
.A1(n_1972),
.A2(n_1945),
.B(n_1931),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1972),
.B(n_1922),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1965),
.A2(n_1935),
.B1(n_1876),
.B2(n_1931),
.Y(n_2008)
);

OAI21xp33_ASAP7_75t_L g2009 ( 
.A1(n_1952),
.A2(n_1907),
.B(n_1906),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1981),
.Y(n_2010)
);

NAND3xp33_ASAP7_75t_SL g2011 ( 
.A(n_1969),
.B(n_1942),
.C(n_1937),
.Y(n_2011)
);

AOI32xp33_ASAP7_75t_L g2012 ( 
.A1(n_1959),
.A2(n_1825),
.A3(n_1831),
.B1(n_1832),
.B2(n_1935),
.Y(n_2012)
);

OAI32xp33_ASAP7_75t_L g2013 ( 
.A1(n_1970),
.A2(n_1944),
.A3(n_1908),
.B1(n_1870),
.B2(n_1872),
.Y(n_2013)
);

AOI21xp33_ASAP7_75t_SL g2014 ( 
.A1(n_1984),
.A2(n_1766),
.B(n_1728),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1961),
.B(n_1966),
.Y(n_2015)
);

AOI22xp5_ASAP7_75t_L g2016 ( 
.A1(n_1959),
.A2(n_1850),
.B1(n_1830),
.B2(n_1845),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1970),
.A2(n_1850),
.B1(n_1830),
.B2(n_1845),
.Y(n_2017)
);

OAI21xp5_ASAP7_75t_SL g2018 ( 
.A1(n_1985),
.A2(n_1738),
.B(n_1732),
.Y(n_2018)
);

OR2x2_ASAP7_75t_L g2019 ( 
.A(n_1980),
.B(n_1944),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1992),
.A2(n_1967),
.B(n_1955),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_2018),
.A2(n_1980),
.B1(n_1850),
.B2(n_1876),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_2010),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_SL g2023 ( 
.A1(n_2018),
.A2(n_1994),
.B(n_1998),
.Y(n_2023)
);

AOI221xp5_ASAP7_75t_L g2024 ( 
.A1(n_2005),
.A2(n_1954),
.B1(n_1957),
.B2(n_1958),
.C(n_1990),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2015),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1991),
.A2(n_1986),
.B1(n_1977),
.B2(n_1950),
.C(n_1938),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2001),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1996),
.B(n_1977),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_2002),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2007),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1997),
.A2(n_1739),
.B1(n_1749),
.B2(n_1775),
.Y(n_2031)
);

INVxp67_ASAP7_75t_L g2032 ( 
.A(n_2004),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_2011),
.B(n_1988),
.Y(n_2033)
);

OAI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_2006),
.A2(n_1982),
.B1(n_1974),
.B2(n_1979),
.C(n_1978),
.Y(n_2034)
);

INVxp67_ASAP7_75t_SL g2035 ( 
.A(n_2003),
.Y(n_2035)
);

O2A1O1Ixp33_ASAP7_75t_L g2036 ( 
.A1(n_1993),
.A2(n_1879),
.B(n_1975),
.C(n_1924),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2019),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2009),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2000),
.B(n_2003),
.Y(n_2039)
);

CKINVDCx16_ASAP7_75t_R g2040 ( 
.A(n_1995),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2008),
.B(n_1983),
.Y(n_2041)
);

AOI322xp5_ASAP7_75t_L g2042 ( 
.A1(n_2017),
.A2(n_1887),
.A3(n_1888),
.B1(n_1886),
.B2(n_1825),
.C1(n_1832),
.C2(n_1831),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2032),
.B(n_2014),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2037),
.Y(n_2044)
);

OAI22xp33_ASAP7_75t_L g2045 ( 
.A1(n_2023),
.A2(n_1999),
.B1(n_2016),
.B2(n_1987),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_2029),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_2028),
.B(n_1924),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2028),
.Y(n_2048)
);

OAI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_2020),
.A2(n_2013),
.B(n_1927),
.Y(n_2049)
);

OAI21xp33_ASAP7_75t_L g2050 ( 
.A1(n_2038),
.A2(n_2041),
.B(n_2033),
.Y(n_2050)
);

XNOR2x1_ASAP7_75t_L g2051 ( 
.A(n_2025),
.B(n_1701),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2039),
.B(n_1924),
.Y(n_2052)
);

INVx1_ASAP7_75t_SL g2053 ( 
.A(n_2040),
.Y(n_2053)
);

INVxp67_ASAP7_75t_L g2054 ( 
.A(n_2035),
.Y(n_2054)
);

AOI31xp33_ASAP7_75t_L g2055 ( 
.A1(n_2027),
.A2(n_1927),
.A3(n_1729),
.B(n_1738),
.Y(n_2055)
);

OAI21xp33_ASAP7_75t_SL g2056 ( 
.A1(n_2021),
.A2(n_2012),
.B(n_1950),
.Y(n_2056)
);

BUFx2_ASAP7_75t_SL g2057 ( 
.A(n_2029),
.Y(n_2057)
);

NOR3xp33_ASAP7_75t_L g2058 ( 
.A(n_2053),
.B(n_2030),
.C(n_2026),
.Y(n_2058)
);

NOR2x1_ASAP7_75t_L g2059 ( 
.A(n_2057),
.B(n_2048),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_2054),
.B(n_2022),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_2024),
.Y(n_2061)
);

NOR2x1_ASAP7_75t_L g2062 ( 
.A(n_2057),
.B(n_1711),
.Y(n_2062)
);

XNOR2xp5_ASAP7_75t_L g2063 ( 
.A(n_2051),
.B(n_2031),
.Y(n_2063)
);

OAI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_2049),
.A2(n_2043),
.B(n_2046),
.C(n_2036),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2044),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_2045),
.A2(n_2031),
.B1(n_2034),
.B2(n_1846),
.Y(n_2066)
);

AOI221xp5_ASAP7_75t_L g2067 ( 
.A1(n_2056),
.A2(n_1938),
.B1(n_1919),
.B2(n_1914),
.C(n_1879),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2051),
.Y(n_2068)
);

NAND2xp67_ASAP7_75t_SL g2069 ( 
.A(n_2047),
.B(n_1886),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_2047),
.B(n_2042),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2052),
.B(n_1886),
.Y(n_2071)
);

OAI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2055),
.A2(n_2052),
.B1(n_1951),
.B2(n_1740),
.C(n_1862),
.Y(n_2072)
);

OAI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2053),
.A2(n_1846),
.B1(n_1830),
.B2(n_1872),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_2061),
.A2(n_1705),
.B(n_1865),
.Y(n_2074)
);

NAND2xp33_ASAP7_75t_SL g2075 ( 
.A(n_2063),
.B(n_1729),
.Y(n_2075)
);

NAND3xp33_ASAP7_75t_SL g2076 ( 
.A(n_2064),
.B(n_1735),
.C(n_1731),
.Y(n_2076)
);

XNOR2xp5_ASAP7_75t_L g2077 ( 
.A(n_2062),
.B(n_1740),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2059),
.B(n_2058),
.Y(n_2078)
);

AOI221xp5_ASAP7_75t_L g2079 ( 
.A1(n_2066),
.A2(n_1825),
.B1(n_1832),
.B2(n_1831),
.C(n_1841),
.Y(n_2079)
);

AOI221x1_ASAP7_75t_L g2080 ( 
.A1(n_2068),
.A2(n_1842),
.B1(n_1841),
.B2(n_1883),
.C(n_1894),
.Y(n_2080)
);

INVx1_ASAP7_75t_SL g2081 ( 
.A(n_2071),
.Y(n_2081)
);

NAND4xp75_ASAP7_75t_L g2082 ( 
.A(n_2060),
.B(n_1832),
.C(n_1831),
.D(n_1896),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2081),
.Y(n_2083)
);

OAI221xp5_ASAP7_75t_SL g2084 ( 
.A1(n_2078),
.A2(n_2070),
.B1(n_2072),
.B2(n_2067),
.C(n_2065),
.Y(n_2084)
);

OAI322xp33_ASAP7_75t_L g2085 ( 
.A1(n_2074),
.A2(n_2073),
.A3(n_2069),
.B1(n_1870),
.B2(n_1872),
.C1(n_1842),
.C2(n_1841),
.Y(n_2085)
);

AOI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_2076),
.A2(n_1842),
.B1(n_1830),
.B2(n_1845),
.C(n_1763),
.Y(n_2086)
);

NOR3xp33_ASAP7_75t_L g2087 ( 
.A(n_2075),
.B(n_2079),
.C(n_2082),
.Y(n_2087)
);

OAI321xp33_ASAP7_75t_L g2088 ( 
.A1(n_2077),
.A2(n_2080),
.A3(n_1819),
.B1(n_1813),
.B2(n_1704),
.C(n_1846),
.Y(n_2088)
);

NOR4xp75_ASAP7_75t_L g2089 ( 
.A(n_2078),
.B(n_1760),
.C(n_1843),
.D(n_1863),
.Y(n_2089)
);

AOI21xp33_ASAP7_75t_L g2090 ( 
.A1(n_2078),
.A2(n_1842),
.B(n_1865),
.Y(n_2090)
);

NAND4xp75_ASAP7_75t_L g2091 ( 
.A(n_2083),
.B(n_1712),
.C(n_1896),
.D(n_1897),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2089),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2088),
.Y(n_2093)
);

BUFx3_ASAP7_75t_L g2094 ( 
.A(n_2084),
.Y(n_2094)
);

NAND2xp33_ASAP7_75t_L g2095 ( 
.A(n_2087),
.B(n_1881),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2086),
.A2(n_1830),
.B1(n_1845),
.B2(n_1887),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_2095),
.A2(n_2090),
.B1(n_2085),
.B2(n_1712),
.Y(n_2097)
);

OR2x2_ASAP7_75t_L g2098 ( 
.A(n_2092),
.B(n_1889),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2094),
.B(n_1896),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_2093),
.B(n_1712),
.Y(n_2100)
);

OAI221xp5_ASAP7_75t_L g2101 ( 
.A1(n_2097),
.A2(n_2096),
.B1(n_2091),
.B2(n_1862),
.C(n_1843),
.Y(n_2101)
);

INVxp67_ASAP7_75t_L g2102 ( 
.A(n_2099),
.Y(n_2102)
);

AO22x2_ASAP7_75t_L g2103 ( 
.A1(n_2102),
.A2(n_2100),
.B1(n_2098),
.B2(n_2096),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_2103),
.Y(n_2104)
);

CKINVDCx20_ASAP7_75t_R g2105 ( 
.A(n_2103),
.Y(n_2105)
);

OAI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_2105),
.A2(n_2101),
.B(n_1897),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2104),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_2107),
.A2(n_1897),
.B1(n_1863),
.B2(n_1843),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2106),
.B(n_1865),
.Y(n_2109)
);

OAI322xp33_ASAP7_75t_L g2110 ( 
.A1(n_2109),
.A2(n_1902),
.A3(n_1883),
.B1(n_1865),
.B2(n_1874),
.C1(n_1901),
.C2(n_1895),
.Y(n_2110)
);

OAI21xp5_ASAP7_75t_SL g2111 ( 
.A1(n_2110),
.A2(n_2108),
.B(n_1704),
.Y(n_2111)
);

OAI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_2111),
.A2(n_1902),
.B1(n_1874),
.B2(n_1901),
.Y(n_2112)
);

AOI221xp5_ASAP7_75t_L g2113 ( 
.A1(n_2112),
.A2(n_1882),
.B1(n_1883),
.B2(n_1874),
.C(n_1901),
.Y(n_2113)
);

AOI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2113),
.A2(n_1643),
.B(n_1709),
.C(n_1715),
.Y(n_2114)
);


endmodule