module real_aes_17061_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_735;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g111 ( .A(n_0), .B(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_1), .A2(n_4), .B1(n_272), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_2), .A2(n_44), .B1(n_153), .B2(n_245), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_3), .A2(n_22), .B1(n_213), .B2(n_245), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_5), .A2(n_15), .B1(n_185), .B2(n_187), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_6), .A2(n_62), .B1(n_149), .B2(n_215), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_7), .A2(n_16), .B1(n_153), .B2(n_158), .Y(n_504) );
INVx1_ASAP7_75t_L g112 ( .A(n_8), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_9), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_10), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_11), .A2(n_17), .B1(n_148), .B2(n_152), .Y(n_147) );
BUFx2_ASAP7_75t_L g106 ( .A(n_12), .Y(n_106) );
OR2x2_ASAP7_75t_L g126 ( .A(n_12), .B(n_39), .Y(n_126) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_13), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_14), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_18), .A2(n_99), .B1(n_185), .B2(n_272), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g176 ( .A1(n_19), .A2(n_40), .B1(n_177), .B2(n_179), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_20), .B(n_186), .Y(n_234) );
OAI21x1_ASAP7_75t_L g164 ( .A1(n_21), .A2(n_59), .B(n_165), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_23), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g136 ( .A1(n_24), .A2(n_55), .B1(n_137), .B2(n_138), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_24), .Y(n_137) );
INVx4_ASAP7_75t_R g529 ( .A(n_25), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_26), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_27), .B(n_156), .Y(n_566) );
INVx1_ASAP7_75t_L g838 ( .A(n_28), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_29), .A2(n_48), .B1(n_198), .B2(n_201), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_30), .A2(n_54), .B1(n_185), .B2(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_31), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_32), .B(n_177), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_33), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_34), .B(n_245), .Y(n_572) );
INVx1_ASAP7_75t_L g611 ( .A(n_35), .Y(n_611) );
A2O1A1Ixp33_ASAP7_75t_SL g547 ( .A1(n_36), .A2(n_153), .B(n_155), .C(n_548), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_37), .Y(n_127) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_38), .A2(n_56), .B1(n_153), .B2(n_201), .Y(n_556) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_41), .A2(n_87), .B1(n_153), .B2(n_212), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_42), .A2(n_80), .B1(n_820), .B2(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_42), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_43), .A2(n_47), .B1(n_153), .B2(n_158), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_45), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_46), .A2(n_61), .B1(n_185), .B2(n_199), .Y(n_274) );
INVx1_ASAP7_75t_L g569 ( .A(n_49), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_50), .B(n_153), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_51), .Y(n_588) );
INVx2_ASAP7_75t_L g488 ( .A(n_52), .Y(n_488) );
BUFx3_ASAP7_75t_L g115 ( .A(n_53), .Y(n_115) );
INVx1_ASAP7_75t_L g124 ( .A(n_53), .Y(n_124) );
INVx1_ASAP7_75t_L g138 ( .A(n_55), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_57), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_58), .A2(n_88), .B1(n_153), .B2(n_201), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_60), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_63), .A2(n_75), .B1(n_198), .B2(n_199), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_64), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_65), .A2(n_77), .B1(n_153), .B2(n_158), .Y(n_222) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_66), .A2(n_98), .B1(n_152), .B2(n_185), .Y(n_221) );
INVx1_ASAP7_75t_L g165 ( .A(n_67), .Y(n_165) );
AND2x4_ASAP7_75t_L g167 ( .A(n_68), .B(n_168), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_69), .A2(n_90), .B1(n_198), .B2(n_201), .Y(n_607) );
AO22x1_ASAP7_75t_L g516 ( .A1(n_70), .A2(n_76), .B1(n_179), .B2(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g168 ( .A(n_71), .Y(n_168) );
AND2x2_ASAP7_75t_L g550 ( .A(n_72), .B(n_240), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_73), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_74), .B(n_215), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_78), .B(n_245), .Y(n_589) );
INVx2_ASAP7_75t_L g156 ( .A(n_79), .Y(n_156) );
INVx1_ASAP7_75t_L g821 ( .A(n_80), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_81), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_82), .B(n_240), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_83), .A2(n_97), .B1(n_201), .B2(n_215), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_84), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_85), .B(n_163), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_86), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_89), .B(n_240), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_91), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_92), .B(n_240), .Y(n_585) );
INVx1_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_93), .B(n_123), .Y(n_122) );
NAND2xp33_ASAP7_75t_L g237 ( .A(n_94), .B(n_186), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_95), .A2(n_160), .B(n_215), .C(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g531 ( .A(n_96), .B(n_532), .Y(n_531) );
NAND2xp33_ASAP7_75t_L g593 ( .A(n_100), .B(n_178), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_116), .B(n_837), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
BUFx4f_ASAP7_75t_L g839 ( .A(n_104), .Y(n_839) );
AND2x6_ASAP7_75t_L g104 ( .A(n_105), .B(n_109), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
INVxp33_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
NOR3x1_ASAP7_75t_L g109 ( .A(n_110), .B(n_113), .C(n_115), .Y(n_109) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AND3x2_ASAP7_75t_L g133 ( .A(n_113), .B(n_125), .C(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g817 ( .A(n_114), .Y(n_817) );
INVx1_ASAP7_75t_L g828 ( .A(n_115), .Y(n_828) );
NOR2x1_ASAP7_75t_L g836 ( .A(n_115), .B(n_126), .Y(n_836) );
OR2x6_ASAP7_75t_L g116 ( .A(n_117), .B(n_128), .Y(n_116) );
NOR2x1_ASAP7_75t_L g129 ( .A(n_117), .B(n_130), .Y(n_129) );
NOR2x1_ASAP7_75t_SL g117 ( .A(n_118), .B(n_127), .Y(n_117) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx8_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_SL g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g134 ( .A(n_124), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_125), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_484), .B(n_489), .Y(n_128) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_135), .Y(n_130) );
BUFx2_ASAP7_75t_SL g131 ( .A(n_132), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
XNOR2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_139), .Y(n_135) );
NAND4xp25_ASAP7_75t_L g139 ( .A(n_140), .B(n_359), .C(n_413), .D(n_452), .Y(n_139) );
NAND4xp75_ASAP7_75t_L g818 ( .A(n_140), .B(n_359), .C(n_413), .D(n_452), .Y(n_818) );
NOR2x1_ASAP7_75t_L g140 ( .A(n_141), .B(n_317), .Y(n_140) );
NAND3xp33_ASAP7_75t_SL g141 ( .A(n_142), .B(n_260), .C(n_299), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_207), .B1(n_250), .B2(n_255), .Y(n_142) );
INVx1_ASAP7_75t_L g423 ( .A(n_143), .Y(n_423) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_172), .Y(n_143) );
INVx1_ASAP7_75t_L g286 ( .A(n_144), .Y(n_286) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_SL g252 ( .A(n_145), .Y(n_252) );
AND2x2_ASAP7_75t_L g304 ( .A(n_145), .B(n_193), .Y(n_304) );
AND2x2_ASAP7_75t_L g343 ( .A(n_145), .B(n_174), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_145), .B(n_280), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_145), .B(n_479), .Y(n_478) );
AO31x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_161), .A3(n_166), .B(n_169), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_154), .B1(n_157), .B2(n_159), .Y(n_146) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_150), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_151), .Y(n_153) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_151), .Y(n_178) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
INVx1_ASAP7_75t_L g188 ( .A(n_151), .Y(n_188) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_151), .Y(n_201) );
INVx2_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
INVx1_ASAP7_75t_L g215 ( .A(n_151), .Y(n_215) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_151), .Y(n_245) );
INVx1_ASAP7_75t_L g273 ( .A(n_151), .Y(n_273) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g158 ( .A(n_153), .Y(n_158) );
INVx1_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_154), .A2(n_176), .B1(n_181), .B2(n_184), .Y(n_175) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_154), .A2(n_181), .B1(n_197), .B2(n_200), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_154), .A2(n_211), .B1(n_214), .B2(n_216), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_154), .A2(n_159), .B1(n_221), .B2(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_154), .A2(n_236), .B(n_237), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_154), .A2(n_181), .B1(n_244), .B2(n_246), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_154), .A2(n_181), .B1(n_271), .B2(n_274), .Y(n_270) );
OAI22x1_ASAP7_75t_L g503 ( .A1(n_154), .A2(n_216), .B1(n_504), .B2(n_505), .Y(n_503) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_154), .A2(n_512), .B1(n_555), .B2(n_556), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_154), .A2(n_216), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx6_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g232 ( .A1(n_155), .A2(n_158), .B(n_233), .C(n_234), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_155), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_155), .A2(n_593), .B(n_594), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_155), .A2(n_511), .B(n_516), .C(n_519), .Y(n_632) );
BUFx8_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g160 ( .A(n_156), .Y(n_160) );
INVx2_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
INVx1_ASAP7_75t_L g546 ( .A(n_156), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_L g587 ( .A1(n_158), .A2(n_588), .B(n_589), .C(n_590), .Y(n_587) );
INVx1_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
AO31x2_ASAP7_75t_L g219 ( .A1(n_161), .A2(n_220), .A3(n_223), .B(n_225), .Y(n_219) );
AOI21x1_ASAP7_75t_L g538 ( .A1(n_161), .A2(n_539), .B(n_550), .Y(n_538) );
AO31x2_ASAP7_75t_L g605 ( .A1(n_161), .A2(n_202), .A3(n_606), .B(n_610), .Y(n_605) );
BUFx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_162), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g532 ( .A(n_162), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_162), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_162), .B(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g170 ( .A(n_163), .Y(n_170) );
INVx2_ASAP7_75t_L g206 ( .A(n_163), .Y(n_206) );
OAI21xp33_ASAP7_75t_L g519 ( .A1(n_163), .A2(n_514), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
AO31x2_ASAP7_75t_L g174 ( .A1(n_166), .A2(n_175), .A3(n_189), .B(n_191), .Y(n_174) );
INVx2_ASAP7_75t_L g224 ( .A(n_166), .Y(n_224) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_166), .A2(n_243), .A3(n_247), .B(n_248), .Y(n_242) );
AO31x2_ASAP7_75t_L g502 ( .A1(n_166), .A2(n_206), .A3(n_503), .B(n_506), .Y(n_502) );
BUFx10_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g203 ( .A(n_167), .Y(n_203) );
INVx1_ASAP7_75t_L g520 ( .A(n_167), .Y(n_520) );
BUFx10_ASAP7_75t_L g557 ( .A(n_167), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g169 ( .A(n_170), .B(n_171), .Y(n_169) );
INVx2_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_170), .B(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g327 ( .A(n_173), .B(n_302), .Y(n_327) );
OR2x2_ASAP7_75t_L g369 ( .A(n_173), .B(n_349), .Y(n_369) );
OR2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_193), .Y(n_173) );
INVx2_ASAP7_75t_L g254 ( .A(n_174), .Y(n_254) );
INVx1_ASAP7_75t_L g280 ( .A(n_174), .Y(n_280) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_174), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_174), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g434 ( .A(n_174), .Y(n_434) );
AND2x2_ASAP7_75t_L g439 ( .A(n_174), .B(n_268), .Y(n_439) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g198 ( .A(n_178), .Y(n_198) );
OAI22xp33_ASAP7_75t_L g528 ( .A1(n_178), .A2(n_188), .B1(n_529), .B2(n_530), .Y(n_528) );
OAI21xp33_ASAP7_75t_SL g565 ( .A1(n_179), .A2(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g512 ( .A(n_182), .Y(n_512) );
BUFx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g591 ( .A(n_183), .Y(n_591) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_186), .Y(n_517) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AO31x2_ASAP7_75t_L g209 ( .A1(n_189), .A2(n_202), .A3(n_210), .B(n_217), .Y(n_209) );
BUFx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_190), .B(n_192), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_190), .B(n_226), .Y(n_225) );
INVx2_ASAP7_75t_SL g230 ( .A(n_190), .Y(n_230) );
INVx4_ASAP7_75t_L g240 ( .A(n_190), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_190), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g573 ( .A(n_190), .B(n_557), .Y(n_573) );
AND2x4_ASAP7_75t_L g253 ( .A(n_193), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g277 ( .A(n_193), .Y(n_277) );
INVx2_ASAP7_75t_L g326 ( .A(n_193), .Y(n_326) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_193), .Y(n_342) );
INVx1_ASAP7_75t_L g479 ( .A(n_193), .Y(n_479) );
AO31x2_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_196), .A3(n_202), .B(n_204), .Y(n_193) );
AO31x2_ASAP7_75t_L g269 ( .A1(n_194), .A2(n_223), .A3(n_270), .B(n_275), .Y(n_269) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_194), .A2(n_523), .B(n_531), .Y(n_522) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_201), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g609 ( .A(n_201), .Y(n_609) );
INVx2_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_SL g238 ( .A(n_203), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_206), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_227), .Y(n_207) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_208), .Y(n_307) );
AND2x2_ASAP7_75t_L g314 ( .A(n_208), .B(n_310), .Y(n_314) );
AND2x2_ASAP7_75t_L g371 ( .A(n_208), .B(n_358), .Y(n_371) );
AND2x4_ASAP7_75t_SL g480 ( .A(n_208), .B(n_282), .Y(n_480) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
BUFx2_ASAP7_75t_L g261 ( .A(n_209), .Y(n_261) );
OR2x2_ASAP7_75t_L g298 ( .A(n_209), .B(n_284), .Y(n_298) );
AND2x4_ASAP7_75t_L g311 ( .A(n_209), .B(n_259), .Y(n_311) );
INVx2_ASAP7_75t_L g339 ( .A(n_209), .Y(n_339) );
OR2x2_ASAP7_75t_L g365 ( .A(n_209), .B(n_242), .Y(n_365) );
INVx1_ASAP7_75t_L g418 ( .A(n_209), .Y(n_418) );
INVx2_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_213), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_216), .B(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g259 ( .A(n_219), .Y(n_259) );
BUFx2_ASAP7_75t_L g337 ( .A(n_219), .Y(n_337) );
AND2x2_ASAP7_75t_L g425 ( .A(n_219), .B(n_339), .Y(n_425) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_224), .A2(n_524), .B(n_527), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_227), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
AND2x4_ASAP7_75t_L g338 ( .A(n_228), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g412 ( .A(n_228), .B(n_259), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_228), .B(n_261), .Y(n_430) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
BUFx2_ASAP7_75t_L g363 ( .A(n_229), .Y(n_363) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_229) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_230), .A2(n_231), .B(n_239), .Y(n_265) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_235), .B(n_238), .Y(n_231) );
INVx2_ASAP7_75t_L g247 ( .A(n_240), .Y(n_247) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_240), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_241), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g283 ( .A(n_241), .Y(n_283) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
INVx1_ASAP7_75t_L g333 ( .A(n_242), .Y(n_333) );
AND2x2_ASAP7_75t_L g358 ( .A(n_242), .B(n_265), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_245), .B(n_542), .Y(n_541) );
AO31x2_ASAP7_75t_L g553 ( .A1(n_247), .A2(n_554), .A3(n_557), .B(n_558), .Y(n_553) );
AND2x2_ASAP7_75t_L g450 ( .A(n_250), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g483 ( .A(n_250), .B(n_348), .Y(n_483) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
INVx1_ASAP7_75t_L g446 ( .A(n_251), .Y(n_446) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g278 ( .A(n_252), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g313 ( .A(n_252), .B(n_268), .Y(n_313) );
INVx1_ASAP7_75t_L g323 ( .A(n_252), .Y(n_323) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_252), .Y(n_330) );
INVx2_ASAP7_75t_L g355 ( .A(n_252), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_252), .B(n_277), .Y(n_368) );
OR2x2_ASAP7_75t_L g377 ( .A(n_252), .B(n_331), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_252), .B(n_325), .Y(n_387) );
AND2x2_ASAP7_75t_L g456 ( .A(n_252), .B(n_434), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_253), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g312 ( .A(n_253), .B(n_313), .Y(n_312) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_253), .Y(n_399) );
NAND2x1p5_ASAP7_75t_L g406 ( .A(n_253), .B(n_289), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_253), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g468 ( .A(n_253), .B(n_354), .Y(n_468) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_256), .A2(n_322), .B1(n_406), .B2(n_407), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_257), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g462 ( .A(n_258), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g482 ( .A(n_258), .B(n_358), .Y(n_482) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g294 ( .A(n_259), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_259), .B(n_283), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_259), .B(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_259), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B1(n_288), .B2(n_292), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_261), .B(n_263), .Y(n_350) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_261), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g465 ( .A(n_261), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B1(n_281), .B2(n_285), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_264), .Y(n_421) );
INVx1_ASAP7_75t_L g463 ( .A(n_264), .Y(n_463) );
INVx1_ASAP7_75t_L g284 ( .A(n_265), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_278), .Y(n_266) );
AOI211xp5_ASAP7_75t_L g351 ( .A1(n_267), .A2(n_352), .B(n_356), .C(n_357), .Y(n_351) );
INVx1_ASAP7_75t_L g389 ( .A(n_267), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_267), .B(n_343), .Y(n_427) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_277), .Y(n_267) );
INVx3_ASAP7_75t_L g349 ( .A(n_268), .Y(n_349) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g287 ( .A(n_269), .B(n_277), .Y(n_287) );
INVx2_ASAP7_75t_L g291 ( .A(n_269), .Y(n_291) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_273), .B(n_544), .Y(n_543) );
NAND2x1_ASAP7_75t_L g370 ( .A(n_278), .B(n_348), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_278), .B(n_341), .Y(n_380) );
INVx1_ASAP7_75t_L g409 ( .A(n_278), .Y(n_409) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_281), .A2(n_467), .B(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g300 ( .A1(n_282), .A2(n_301), .B(n_305), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_282), .B(n_436), .Y(n_472) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx3_ASAP7_75t_L g331 ( .A(n_287), .Y(n_331) );
AND2x4_ASAP7_75t_L g449 ( .A(n_287), .B(n_316), .Y(n_449) );
AND2x2_ASAP7_75t_L g455 ( .A(n_287), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g386 ( .A(n_289), .Y(n_386) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g306 ( .A(n_290), .B(n_297), .Y(n_306) );
AND2x2_ASAP7_75t_L g432 ( .A(n_290), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g303 ( .A(n_291), .Y(n_303) );
OR2x2_ASAP7_75t_L g353 ( .A(n_291), .B(n_326), .Y(n_353) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_295), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NOR2x1p5_ASAP7_75t_L g364 ( .A(n_294), .B(n_365), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_294), .B(n_298), .Y(n_451) );
INVx1_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
NOR2x1_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NOR2xp67_ASAP7_75t_SL g381 ( .A(n_298), .B(n_382), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_307), .B1(n_308), .B2(n_312), .C1(n_314), .C2(n_315), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g344 ( .A1(n_301), .A2(n_345), .B(n_350), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_302), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g469 ( .A(n_302), .Y(n_469) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_303), .Y(n_475) );
AND2x4_ASAP7_75t_L g315 ( .A(n_304), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_304), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g459 ( .A(n_304), .Y(n_459) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
AND2x2_ASAP7_75t_L g400 ( .A(n_309), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g393 ( .A(n_310), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_334), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B1(n_328), .B2(n_332), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp33_ASAP7_75t_L g321 ( .A(n_322), .B(n_327), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g346 ( .A(n_324), .Y(n_346) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
AND2x4_ASAP7_75t_L g383 ( .A(n_333), .B(n_338), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_333), .B(n_436), .Y(n_435) );
AOI211x1_ASAP7_75t_SL g334 ( .A1(n_335), .A2(n_340), .B(n_344), .C(n_351), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_335), .A2(n_449), .B(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_338), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g401 ( .A(n_337), .B(n_338), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_338), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_338), .Y(n_394) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g458 ( .A(n_341), .B(n_439), .Y(n_458) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g356 ( .A(n_343), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_343), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g376 ( .A(n_349), .B(n_368), .Y(n_376) );
OR2x2_ASAP7_75t_L g477 ( .A(n_349), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_353), .Y(n_410) );
INVx2_ASAP7_75t_L g447 ( .A(n_353), .Y(n_447) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND5xp2_ASAP7_75t_L g453 ( .A(n_356), .B(n_406), .C(n_454), .D(n_457), .E(n_459), .Y(n_453) );
AND2x2_ASAP7_75t_L g424 ( .A(n_358), .B(n_425), .Y(n_424) );
NOR2x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_397), .Y(n_359) );
NAND2xp67_ASAP7_75t_SL g360 ( .A(n_361), .B(n_378), .Y(n_360) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B1(n_371), .B2(n_372), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .C(n_370), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g403 ( .A(n_370), .Y(n_403) );
NAND3xp33_ASAP7_75t_SL g372 ( .A(n_373), .B(n_376), .C(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g396 ( .A(n_375), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_SL g408 ( .A1(n_376), .A2(n_409), .B(n_410), .C(n_411), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B1(n_383), .B2(n_384), .C(n_388), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_385), .B(n_474), .Y(n_473) );
OR2x2_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_393), .B2(n_395), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g440 ( .A1(n_389), .A2(n_415), .B(n_441), .C(n_443), .Y(n_440) );
INVx1_ASAP7_75t_L g404 ( .A(n_390), .Y(n_404) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g429 ( .A(n_392), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_402), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g407 ( .A(n_401), .Y(n_407) );
AOI211xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_405), .C(n_408), .Y(n_402) );
AND3x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_440), .C(n_448), .Y(n_413) );
AOI221x1_ASAP7_75t_SL g414 ( .A1(n_415), .A2(n_422), .B1(n_424), .B2(n_426), .C(n_428), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_431), .B1(n_435), .B2(n_438), .Y(n_428) );
INVx1_ASAP7_75t_L g442 ( .A(n_433), .Y(n_442) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
AOI211x1_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_460), .B(n_466), .C(n_481), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_473), .B1(n_476), .B2(n_480), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g826 ( .A(n_488), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_488), .B(n_834), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_824), .B(n_829), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_819), .B1(n_822), .B2(n_823), .Y(n_490) );
INVx2_ASAP7_75t_L g822 ( .A(n_491), .Y(n_822) );
AO22x2_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_814), .B1(n_815), .B2(n_818), .Y(n_491) );
INVx1_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
NOR2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_728), .Y(n_493) );
NAND4xp75_ASAP7_75t_L g494 ( .A(n_495), .B(n_633), .C(n_675), .D(n_699), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_533), .B(n_574), .C(n_612), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g719 ( .A(n_499), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g813 ( .A(n_499), .B(n_750), .Y(n_813) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_508), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g628 ( .A(n_501), .B(n_584), .Y(n_628) );
AND2x2_ASAP7_75t_L g669 ( .A(n_501), .B(n_630), .Y(n_669) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g580 ( .A(n_502), .B(n_522), .Y(n_580) );
OR2x2_ASAP7_75t_L g598 ( .A(n_502), .B(n_522), .Y(n_598) );
INVx2_ASAP7_75t_L g620 ( .A(n_502), .Y(n_620) );
AND2x2_ASAP7_75t_L g650 ( .A(n_502), .B(n_584), .Y(n_650) );
AND2x2_ASAP7_75t_L g679 ( .A(n_502), .B(n_521), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_502), .B(n_631), .Y(n_715) );
AND2x2_ASAP7_75t_L g692 ( .A(n_508), .B(n_621), .Y(n_692) );
INVx2_ASAP7_75t_L g787 ( .A(n_508), .Y(n_787) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
INVx2_ASAP7_75t_L g579 ( .A(n_509), .Y(n_579) );
AND2x4_ASAP7_75t_L g618 ( .A(n_509), .B(n_522), .Y(n_618) );
AOI21x1_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_515), .B(n_518), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI21x1_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_514), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_512), .A2(n_571), .B(n_572), .Y(n_570) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_520), .A2(n_540), .B(n_547), .Y(n_539) );
AND2x2_ASAP7_75t_L g777 ( .A(n_521), .B(n_579), .Y(n_777) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g641 ( .A(n_522), .Y(n_641) );
AND2x2_ASAP7_75t_L g698 ( .A(n_522), .B(n_584), .Y(n_698) );
AND2x2_ASAP7_75t_L g713 ( .A(n_522), .B(n_621), .Y(n_713) );
AND2x2_ASAP7_75t_L g735 ( .A(n_522), .B(n_579), .Y(n_735) );
OAI211xp5_ASAP7_75t_SL g782 ( .A1(n_533), .A2(n_783), .B(n_785), .C(n_792), .Y(n_782) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_560), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g769 ( .A(n_536), .B(n_705), .Y(n_769) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_551), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_537), .B(n_562), .Y(n_668) );
INVxp67_ASAP7_75t_L g682 ( .A(n_537), .Y(n_682) );
AND2x2_ASAP7_75t_L g702 ( .A(n_537), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_537), .B(n_615), .Y(n_709) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g602 ( .A(n_538), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_543), .B(n_545), .Y(n_540) );
BUFx4f_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_546), .B(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g643 ( .A(n_551), .B(n_625), .Y(n_643) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g691 ( .A(n_552), .B(n_602), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_552), .B(n_605), .Y(n_697) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g601 ( .A(n_553), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g666 ( .A(n_553), .B(n_605), .Y(n_666) );
BUFx2_ASAP7_75t_L g673 ( .A(n_553), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_553), .B(n_605), .Y(n_753) );
INVx1_ASAP7_75t_L g596 ( .A(n_557), .Y(n_596) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g683 ( .A(n_561), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g812 ( .A(n_561), .B(n_601), .Y(n_812) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx3_ASAP7_75t_L g615 ( .A(n_562), .Y(n_615) );
AND2x2_ASAP7_75t_L g626 ( .A(n_562), .B(n_605), .Y(n_626) );
AND2x2_ASAP7_75t_L g672 ( .A(n_562), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g705 ( .A(n_562), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_562), .B(n_616), .Y(n_722) );
AND2x2_ASAP7_75t_L g761 ( .A(n_562), .B(n_762), .Y(n_761) );
AND2x4_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_570), .B(n_573), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_581), .B(n_599), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_576), .A2(n_740), .B1(n_741), .B2(n_743), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
AND2x2_ASAP7_75t_L g737 ( .A(n_577), .B(n_628), .Y(n_737) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g652 ( .A(n_578), .Y(n_652) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g801 ( .A(n_579), .B(n_621), .Y(n_801) );
AND2x2_ASAP7_75t_L g765 ( .A(n_580), .B(n_660), .Y(n_765) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_597), .Y(n_581) );
OR2x2_ASAP7_75t_L g662 ( .A(n_582), .B(n_639), .Y(n_662) );
OR2x2_ASAP7_75t_L g774 ( .A(n_582), .B(n_598), .Y(n_774) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g637 ( .A(n_583), .Y(n_637) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g621 ( .A(n_584), .Y(n_621) );
BUFx3_ASAP7_75t_L g703 ( .A(n_584), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_592), .B(n_595), .Y(n_586) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g771 ( .A(n_598), .B(n_630), .Y(n_771) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
AND2x2_ASAP7_75t_L g613 ( .A(n_601), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g654 ( .A(n_601), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g791 ( .A(n_601), .Y(n_791) );
INVx1_ASAP7_75t_L g810 ( .A(n_601), .Y(n_810) );
INVx2_ASAP7_75t_L g625 ( .A(n_602), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_602), .B(n_605), .Y(n_674) );
INVx1_ASAP7_75t_L g738 ( .A(n_603), .Y(n_738) );
BUFx3_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g799 ( .A(n_604), .Y(n_799) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g616 ( .A(n_605), .Y(n_616) );
INVx1_ASAP7_75t_L g706 ( .A(n_605), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_617), .B1(n_622), .B2(n_627), .Y(n_612) );
AND2x4_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx2_ASAP7_75t_L g655 ( .A(n_615), .Y(n_655) );
AND2x2_ASAP7_75t_L g657 ( .A(n_615), .B(n_642), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_615), .B(n_625), .Y(n_717) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx3_ASAP7_75t_L g648 ( .A(n_618), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_618), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g742 ( .A(n_618), .B(n_726), .Y(n_742) );
INVx1_ASAP7_75t_L g646 ( .A(n_619), .Y(n_646) );
AOI222xp33_ASAP7_75t_L g656 ( .A1(n_619), .A2(n_657), .B1(n_658), .B2(n_663), .C1(n_669), .C2(n_670), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_619), .A2(n_687), .B(n_688), .Y(n_686) );
AND2x2_ASAP7_75t_L g710 ( .A(n_619), .B(n_629), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_619), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
OR2x2_ASAP7_75t_L g639 ( .A(n_620), .B(n_631), .Y(n_639) );
INVx1_ASAP7_75t_L g727 ( .A(n_620), .Y(n_727) );
BUFx2_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_624), .B(n_665), .Y(n_694) );
OR2x2_ASAP7_75t_L g806 ( .A(n_624), .B(n_666), .Y(n_806) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x4_ASAP7_75t_L g689 ( .A(n_626), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g804 ( .A(n_626), .Y(n_804) );
OAI31xp33_ASAP7_75t_L g785 ( .A1(n_627), .A2(n_786), .A3(n_788), .B(n_789), .Y(n_785) );
AND2x4_ASAP7_75t_SL g627 ( .A(n_628), .B(n_629), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_628), .B(n_777), .Y(n_776) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_656), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_642), .B(n_644), .Y(n_634) );
NOR2x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x6_ASAP7_75t_L g755 ( .A(n_637), .B(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
INVx1_ASAP7_75t_L g687 ( .A(n_640), .Y(n_687) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g778 ( .A(n_641), .B(n_715), .Y(n_778) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_643), .A2(n_732), .B1(n_734), .B2(n_736), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g792 ( .A1(n_643), .A2(n_704), .B(n_766), .C(n_793), .Y(n_792) );
AOI21xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_649), .B(n_653), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g745 ( .A(n_648), .B(n_746), .C(n_747), .D(n_749), .Y(n_745) );
NAND2x1_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_650), .B(n_652), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_650), .B(n_735), .Y(n_758) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g724 ( .A(n_655), .B(n_684), .Y(n_724) );
NAND2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_662), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_662), .A2(n_806), .B1(n_807), .B2(n_809), .Y(n_805) );
AOI221x1_ASAP7_75t_L g744 ( .A1(n_663), .A2(n_745), .B1(n_751), .B2(n_754), .C(n_757), .Y(n_744) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_667), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g684 ( .A(n_666), .Y(n_684) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g696 ( .A(n_668), .B(n_697), .Y(n_696) );
NAND2x1p5_ASAP7_75t_L g759 ( .A(n_669), .B(n_750), .Y(n_759) );
O2A1O1Ixp5_ASAP7_75t_L g772 ( .A1(n_670), .A2(n_754), .B(n_773), .C(n_775), .Y(n_772) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
INVx2_ASAP7_75t_L g721 ( .A(n_673), .Y(n_721) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_685), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_677), .A2(n_695), .B1(n_765), .B2(n_766), .C(n_768), .Y(n_764) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g701 ( .A(n_679), .B(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_679), .B(n_750), .Y(n_749) );
AND2x2_ASAP7_75t_L g800 ( .A(n_679), .B(n_801), .Y(n_800) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVxp67_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
NAND2x1_ASAP7_75t_L g779 ( .A(n_682), .B(n_780), .Y(n_779) );
OR2x2_ASAP7_75t_L g803 ( .A(n_682), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g743 ( .A(n_683), .Y(n_743) );
AOI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_692), .B2(n_693), .C1(n_695), .C2(n_698), .Y(n_685) );
INVx1_ASAP7_75t_L g770 ( .A(n_689), .Y(n_770) );
INVx1_ASAP7_75t_L g733 ( .A(n_690), .Y(n_733) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g767 ( .A(n_691), .Y(n_767) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g708 ( .A(n_697), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g762 ( .A(n_697), .Y(n_762) );
AND2x2_ASAP7_75t_L g725 ( .A(n_698), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_718), .Y(n_699) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_704), .B1(n_707), .B2(n_710), .C1(n_711), .C2(n_716), .Y(n_700) );
INVx3_ASAP7_75t_L g750 ( .A(n_703), .Y(n_750) );
BUFx2_ASAP7_75t_L g808 ( .A(n_703), .Y(n_808) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g780 ( .A(n_705), .Y(n_780) );
OR2x2_ASAP7_75t_L g790 ( .A(n_705), .B(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx2_ASAP7_75t_SL g748 ( .A(n_713), .Y(n_748) );
AND2x2_ASAP7_75t_L g793 ( .A(n_714), .B(n_750), .Y(n_793) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_715), .Y(n_746) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g752 ( .A(n_717), .B(n_753), .Y(n_752) );
NOR2x1_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
OR2x2_ASAP7_75t_L g809 ( .A(n_722), .B(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g740 ( .A(n_724), .Y(n_740) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g747 ( .A(n_727), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g797 ( .A(n_727), .Y(n_797) );
NAND4xp75_ASAP7_75t_L g728 ( .A(n_729), .B(n_763), .C(n_781), .D(n_794), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_744), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_738), .B(n_739), .Y(n_730) );
INVxp33_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_733), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g756 ( .A(n_735), .Y(n_756) );
AND2x2_ASAP7_75t_L g796 ( .A(n_735), .B(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g766 ( .A(n_738), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g784 ( .A(n_749), .Y(n_784) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI22xp33_ASAP7_75t_SL g775 ( .A1(n_752), .A2(n_776), .B1(n_778), .B2(n_779), .Y(n_775) );
INVx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AOI21xp33_ASAP7_75t_SL g757 ( .A1(n_758), .A2(n_759), .B(n_760), .Y(n_757) );
INVx1_ASAP7_75t_L g788 ( .A(n_759), .Y(n_788) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
AND2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_772), .Y(n_763) );
AOI21xp5_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_770), .B(n_771), .Y(n_768) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx3_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_811), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_798), .B1(n_800), .B2(n_802), .C(n_805), .Y(n_795) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
BUFx12f_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_817), .Y(n_816) );
AND2x2_ASAP7_75t_L g835 ( .A(n_817), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g823 ( .A(n_819), .Y(n_823) );
BUFx12f_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AND2x6_ASAP7_75t_SL g825 ( .A(n_826), .B(n_827), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
INVx5_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
BUFx10_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NOR2xp33_ASAP7_75t_SL g837 ( .A(n_838), .B(n_839), .Y(n_837) );
endmodule