module fake_netlist_5_688_n_1030 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_1030);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1030;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_419;
wire n_380;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_785;
wire n_316;
wire n_855;
wire n_389;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_998;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_612;
wire n_1001;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_947;
wire n_373;
wire n_820;
wire n_936;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_1024;
wire n_556;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_394;
wire n_579;
wire n_250;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_449;
wire n_325;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_647;
wire n_240;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_696;
wire n_255;
wire n_897;
wire n_798;
wire n_350;
wire n_1020;
wire n_662;
wire n_459;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_681;
wire n_584;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_673;
wire n_631;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_680;
wire n_974;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_249;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_693;
wire n_571;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_1028;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_736;
wire n_595;
wire n_502;
wire n_892;
wire n_893;
wire n_1015;
wire n_1000;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_607;
wire n_575;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_710;
wire n_707;
wire n_795;
wire n_832;
wire n_695;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_403;
wire n_453;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_233;
wire n_686;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_895;
wire n_644;
wire n_728;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1025;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_666;
wire n_538;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_100),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_21),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_89),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_221),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_165),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_95),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_15),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_96),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_78),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_182),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

CKINVDCx11_ASAP7_75t_R g240 ( 
.A(n_177),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_181),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_154),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_214),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_19),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_149),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_27),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_29),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_69),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_86),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_72),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_12),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_39),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_53),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_73),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_77),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_156),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_218),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_9),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_205),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_36),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_84),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_193),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_60),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_106),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_158),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_110),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_211),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_21),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_219),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_163),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_27),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_12),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_20),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_208),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_178),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_5),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_85),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_9),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_45),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_81),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_200),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_151),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_117),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_121),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_135),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_137),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_152),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_6),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_146),
.Y(n_302)
);

BUFx5_ASAP7_75t_L g303 ( 
.A(n_35),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_93),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_63),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_161),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_16),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_195),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_171),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_179),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_141),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_170),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_24),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_105),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_189),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_124),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_198),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_122),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_104),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_36),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_150),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_103),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_33),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_0),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g327 ( 
.A(n_237),
.B(n_41),
.Y(n_327)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_247),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_242),
.B(n_0),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_303),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_237),
.B(n_42),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_1),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_291),
.B(n_1),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_2),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_274),
.B(n_43),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_264),
.B(n_2),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_3),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_240),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_3),
.Y(n_342)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_274),
.B(n_4),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

INVx5_ASAP7_75t_L g346 ( 
.A(n_247),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_305),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_303),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_296),
.B(n_4),
.Y(n_349)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_305),
.Y(n_350)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_245),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_44),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_262),
.B(n_306),
.Y(n_353)
);

BUFx8_ASAP7_75t_SL g354 ( 
.A(n_246),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_315),
.B(n_5),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_226),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_244),
.B(n_6),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_262),
.B(n_7),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_245),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_225),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_245),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_232),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_245),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_314),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_249),
.B(n_7),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_243),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_236),
.B(n_8),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_239),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_250),
.B(n_255),
.Y(n_370)
);

BUFx12f_ASAP7_75t_L g371 ( 
.A(n_240),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_257),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_259),
.B(n_8),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_260),
.B(n_46),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_224),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_261),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_270),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_318),
.B(n_10),
.Y(n_378)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_227),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_279),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_251),
.B(n_256),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_354),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_338),
.B1(n_330),
.B2(n_339),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_363),
.B(n_347),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_359),
.A2(n_291),
.B1(n_297),
.B2(n_276),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_228),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_351),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_267),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_335),
.A2(n_268),
.B1(n_324),
.B2(n_266),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_358),
.A2(n_297),
.B1(n_258),
.B2(n_284),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_357),
.B(n_229),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_378),
.A2(n_283),
.B1(n_301),
.B2(n_246),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_351),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_321),
.B1(n_289),
.B2(n_287),
.Y(n_395)
);

BUFx10_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_329),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_360),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_360),
.Y(n_400)
);

NOR2x1p5_ASAP7_75t_L g401 ( 
.A(n_371),
.B(n_282),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_321),
.B1(n_307),
.B2(n_272),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_363),
.A2(n_340),
.B1(n_381),
.B2(n_373),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_364),
.Y(n_404)
);

INVx3_ASAP7_75t_SL g405 ( 
.A(n_365),
.Y(n_405)
);

AO22x2_ASAP7_75t_L g406 ( 
.A1(n_327),
.A2(n_269),
.B1(n_273),
.B2(n_275),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_344),
.A2(n_323),
.B1(n_322),
.B2(n_230),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

AO22x2_ASAP7_75t_L g412 ( 
.A1(n_327),
.A2(n_333),
.B1(n_352),
.B2(n_337),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_L g413 ( 
.A1(n_371),
.A2(n_320),
.B1(n_281),
.B2(n_285),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_344),
.A2(n_295),
.B1(n_302),
.B2(n_316),
.Y(n_414)
);

OAI22xp33_ASAP7_75t_L g415 ( 
.A1(n_326),
.A2(n_304),
.B1(n_309),
.B2(n_311),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_327),
.A2(n_337),
.B1(n_352),
.B2(n_333),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_333),
.A2(n_319),
.B1(n_317),
.B2(n_313),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_337),
.A2(n_277),
.B1(n_310),
.B2(n_308),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_231),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_352),
.A2(n_271),
.B1(n_299),
.B2(n_298),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_L g421 ( 
.A1(n_334),
.A2(n_312),
.B1(n_294),
.B2(n_293),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_365),
.Y(n_422)
);

AO22x2_ASAP7_75t_L g423 ( 
.A1(n_366),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_343),
.A2(n_292),
.B1(n_290),
.B2(n_288),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_374),
.A2(n_252),
.B1(n_280),
.B2(n_278),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_365),
.B(n_233),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_374),
.A2(n_248),
.B1(n_265),
.B2(n_263),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_331),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_356),
.Y(n_429)
);

OA22x2_ASAP7_75t_L g430 ( 
.A1(n_377),
.A2(n_286),
.B1(n_254),
.B2(n_253),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_374),
.A2(n_238),
.B1(n_235),
.B2(n_234),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_365),
.B(n_241),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_343),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_366),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_342),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_R g438 ( 
.A1(n_349),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_384),
.B(n_375),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_382),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_416),
.B(n_365),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_428),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_347),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_392),
.B(n_375),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_385),
.B(n_375),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_370),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_430),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_411),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_393),
.B(n_361),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_407),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_394),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_397),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_391),
.B(n_361),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_408),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_429),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

AND2x2_ASAP7_75t_SL g466 ( 
.A(n_435),
.B(n_355),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_402),
.B(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_418),
.B(n_379),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_440),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_423),
.B(n_367),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_SL g474 ( 
.A(n_433),
.B(n_336),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_419),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_412),
.B(n_379),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_420),
.B(n_332),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_425),
.B(n_379),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_439),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_439),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_406),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_R g487 ( 
.A(n_390),
.B(n_23),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g488 ( 
.A(n_436),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_424),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_379),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_423),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_427),
.A2(n_348),
.B(n_345),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_422),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_396),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_383),
.B(n_47),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_431),
.A2(n_348),
.B(n_345),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_401),
.B(n_23),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_396),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_426),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_415),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_403),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_421),
.B(n_379),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_413),
.B(n_379),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_395),
.B(n_350),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_438),
.B(n_377),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

BUFx5_ASAP7_75t_L g511 ( 
.A(n_411),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_382),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_382),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_382),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_382),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_SL g517 ( 
.A(n_433),
.B(n_367),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_453),
.B(n_356),
.Y(n_518)
);

AND2x2_ASAP7_75t_SL g519 ( 
.A(n_466),
.B(n_369),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_453),
.A2(n_362),
.B(n_350),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_471),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g522 ( 
.A(n_503),
.B(n_380),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_451),
.B(n_380),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_449),
.B(n_376),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_442),
.B(n_376),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_442),
.B(n_369),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_493),
.A2(n_362),
.B(n_350),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_489),
.B(n_369),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_441),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_447),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_447),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_457),
.Y(n_535)
);

HB1xp67_ASAP7_75t_L g536 ( 
.A(n_471),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_476),
.B(n_369),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_478),
.B(n_369),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_458),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_483),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_492),
.B(n_484),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_478),
.B(n_501),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_450),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_503),
.B(n_350),
.Y(n_545)
);

NAND2x1p5_ASAP7_75t_L g546 ( 
.A(n_501),
.B(n_444),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_500),
.Y(n_547)
);

BUFx5_ASAP7_75t_L g548 ( 
.A(n_478),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_461),
.B(n_372),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_456),
.B(n_372),
.Y(n_550)
);

AND2x2_ASAP7_75t_SL g551 ( 
.A(n_466),
.B(n_372),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_478),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_455),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_467),
.B(n_350),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_471),
.B(n_372),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

AND2x2_ASAP7_75t_SL g558 ( 
.A(n_467),
.B(n_372),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_490),
.B(n_376),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_478),
.Y(n_560)
);

OR2x2_ASAP7_75t_SL g561 ( 
.A(n_508),
.B(n_376),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_495),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_502),
.B(n_376),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_459),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_498),
.B(n_350),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_477),
.A2(n_362),
.B(n_328),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_507),
.B(n_24),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_485),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_R g569 ( 
.A(n_487),
.B(n_49),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_446),
.B(n_362),
.Y(n_570)
);

OAI21x1_ASAP7_75t_L g571 ( 
.A1(n_444),
.A2(n_362),
.B(n_328),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_460),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_448),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_510),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_487),
.B(n_50),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_481),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_509),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_481),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_454),
.B(n_486),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_512),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_513),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_488),
.B(n_329),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_514),
.B(n_362),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_515),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_496),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_516),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_511),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_511),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_507),
.B(n_506),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_463),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_474),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_488),
.B(n_329),
.Y(n_593)
);

AND2x2_ASAP7_75t_SL g594 ( 
.A(n_504),
.B(n_469),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_511),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_464),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_509),
.B(n_329),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_465),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_511),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_504),
.B(n_325),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_491),
.B(n_51),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_511),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_474),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_468),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_325),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_531),
.B(n_505),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_526),
.B(n_480),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_540),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_592),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_526),
.B(n_594),
.Y(n_610)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_531),
.B(n_497),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_580),
.B(n_494),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_594),
.B(n_480),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_580),
.B(n_586),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_568),
.B(n_508),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_524),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_532),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_588),
.Y(n_619)
);

NAND2x1p5_ASAP7_75t_L g620 ( 
.A(n_552),
.B(n_496),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_580),
.B(n_469),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_552),
.B(n_472),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_523),
.B(n_499),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_533),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_523),
.B(n_530),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_519),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_549),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_577),
.B(n_517),
.Y(n_629)
);

BUFx12f_ASAP7_75t_L g630 ( 
.A(n_562),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_583),
.B(n_473),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_533),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_534),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_534),
.Y(n_634)
);

NOR2xp67_ASAP7_75t_L g635 ( 
.A(n_547),
.B(n_475),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_586),
.B(n_479),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_590),
.B(n_517),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_519),
.B(n_482),
.Y(n_638)
);

OR2x6_ASAP7_75t_L g639 ( 
.A(n_521),
.B(n_25),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_522),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_556),
.B(n_52),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_553),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_556),
.B(n_54),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_592),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_549),
.B(n_550),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g646 ( 
.A(n_522),
.B(n_597),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_536),
.B(n_25),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_551),
.B(n_26),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_576),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_547),
.Y(n_650)
);

INVx6_ASAP7_75t_L g651 ( 
.A(n_583),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_535),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_593),
.B(n_55),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_550),
.B(n_26),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_540),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_597),
.B(n_56),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g657 ( 
.A(n_558),
.B(n_567),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_593),
.B(n_28),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_525),
.Y(n_659)
);

AOI21x1_ASAP7_75t_L g660 ( 
.A1(n_518),
.A2(n_346),
.B(n_328),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_576),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_576),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_535),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_548),
.B(n_325),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_559),
.B(n_28),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_560),
.B(n_565),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_561),
.B(n_29),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_539),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_563),
.B(n_30),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_539),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_554),
.B(n_57),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_659),
.Y(n_673)
);

BUFx2_ASAP7_75t_SL g674 ( 
.A(n_650),
.Y(n_674)
);

INVxp67_ASAP7_75t_SL g675 ( 
.A(n_659),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_615),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_652),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_665),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_630),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_645),
.B(n_610),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_609),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_657),
.A2(n_603),
.B1(n_558),
.B2(n_551),
.Y(n_682)
);

INVxp67_ASAP7_75t_SL g683 ( 
.A(n_615),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_663),
.Y(n_684)
);

BUFx5_ASAP7_75t_L g685 ( 
.A(n_667),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_644),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_669),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_610),
.B(n_548),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_651),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_661),
.Y(n_690)
);

CKINVDCx8_ASAP7_75t_R g691 ( 
.A(n_608),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_661),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_624),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_619),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_671),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_661),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_667),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_619),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_629),
.Y(n_699)
);

INVx6_ASAP7_75t_L g700 ( 
.A(n_651),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_619),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_617),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_639),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_637),
.B(n_563),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_618),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_608),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_619),
.Y(n_707)
);

CKINVDCx6p67_ASAP7_75t_R g708 ( 
.A(n_639),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_612),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

BUFx8_ASAP7_75t_L g711 ( 
.A(n_608),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_611),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_632),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_622),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_657),
.A2(n_603),
.B1(n_560),
.B2(n_527),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_637),
.Y(n_716)
);

INVx5_ASAP7_75t_L g717 ( 
.A(n_667),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_655),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_625),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_639),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_626),
.B(n_525),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_662),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_662),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_655),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_662),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_634),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_633),
.Y(n_727)
);

INVx6_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_716),
.A2(n_614),
.B1(n_651),
.B2(n_627),
.Y(n_729)
);

BUFx2_ASAP7_75t_SL g730 ( 
.A(n_691),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_709),
.Y(n_731)
);

AOI22xp33_ASAP7_75t_L g732 ( 
.A1(n_704),
.A2(n_648),
.B1(n_614),
.B2(n_666),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_677),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_716),
.A2(n_627),
.B1(n_607),
.B2(n_646),
.Y(n_734)
);

BUFx8_ASAP7_75t_L g735 ( 
.A(n_678),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_693),
.A2(n_648),
.B1(n_621),
.B2(n_606),
.Y(n_736)
);

CKINVDCx11_ASAP7_75t_R g737 ( 
.A(n_681),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_711),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_684),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_690),
.Y(n_740)
);

BUFx4_ASAP7_75t_R g741 ( 
.A(n_679),
.Y(n_741)
);

BUFx4f_ASAP7_75t_SL g742 ( 
.A(n_711),
.Y(n_742)
);

CKINVDCx11_ASAP7_75t_R g743 ( 
.A(n_681),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_682),
.A2(n_607),
.B1(n_621),
.B2(n_640),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_691),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_686),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_698),
.A2(n_599),
.B(n_588),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_710),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_680),
.A2(n_606),
.B1(n_643),
.B2(n_641),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_680),
.A2(n_643),
.B1(n_641),
.B2(n_569),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_704),
.A2(n_699),
.B1(n_575),
.B2(n_712),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_L g752 ( 
.A1(n_721),
.A2(n_656),
.B1(n_672),
.B2(n_654),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_L g753 ( 
.A1(n_688),
.A2(n_656),
.B1(n_672),
.B2(n_668),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_715),
.A2(n_628),
.B1(n_647),
.B2(n_543),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_690),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_687),
.Y(n_756)
);

CKINVDCx11_ASAP7_75t_R g757 ( 
.A(n_686),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_683),
.B(n_628),
.Y(n_758)
);

CKINVDCx20_ASAP7_75t_R g759 ( 
.A(n_679),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_695),
.A2(n_670),
.B1(n_658),
.B2(n_642),
.Y(n_760)
);

BUFx2_ASAP7_75t_SL g761 ( 
.A(n_706),
.Y(n_761)
);

BUFx2_ASAP7_75t_SL g762 ( 
.A(n_706),
.Y(n_762)
);

BUFx12f_ASAP7_75t_L g763 ( 
.A(n_703),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_702),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_SL g765 ( 
.A1(n_720),
.A2(n_548),
.B1(n_647),
.B2(n_703),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_690),
.Y(n_766)
);

OAI21xp33_ASAP7_75t_L g767 ( 
.A1(n_673),
.A2(n_647),
.B(n_557),
.Y(n_767)
);

INVx2_ASAP7_75t_SL g768 ( 
.A(n_718),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_709),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_705),
.A2(n_548),
.B1(n_555),
.B2(n_638),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_697),
.A2(n_638),
.B1(n_546),
.B2(n_655),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_714),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_719),
.A2(n_548),
.B1(n_581),
.B2(n_587),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_697),
.B(n_649),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_697),
.A2(n_717),
.B1(n_700),
.B2(n_546),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_675),
.B(n_541),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_727),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_737),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_728),
.A2(n_720),
.B1(n_548),
.B2(n_674),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_767),
.A2(n_708),
.B1(n_582),
.B2(n_585),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_732),
.A2(n_548),
.B1(n_557),
.B2(n_554),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_732),
.A2(n_734),
.B1(n_744),
.B2(n_754),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_748),
.B(n_746),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_750),
.A2(n_561),
.B1(n_635),
.B2(n_697),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_751),
.B(n_724),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_754),
.A2(n_765),
.B1(n_736),
.B2(n_729),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_765),
.B(n_676),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_R g788 ( 
.A(n_743),
.B(n_718),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_760),
.A2(n_548),
.B1(n_587),
.B2(n_581),
.Y(n_789)
);

BUFx4f_ASAP7_75t_SL g790 ( 
.A(n_735),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_752),
.A2(n_708),
.B1(n_585),
.B2(n_582),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_731),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_733),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_745),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_739),
.B(n_676),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_758),
.Y(n_796)
);

AND2x6_ASAP7_75t_L g797 ( 
.A(n_776),
.B(n_694),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_SL g798 ( 
.A1(n_728),
.A2(n_697),
.B1(n_717),
.B2(n_667),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_760),
.A2(n_573),
.B1(n_596),
.B2(n_591),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_749),
.B(n_689),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_756),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_753),
.A2(n_574),
.B1(n_601),
.B2(n_573),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_764),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_770),
.A2(n_574),
.B1(n_601),
.B2(n_688),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_772),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_777),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_766),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_L g809 ( 
.A1(n_742),
.A2(n_717),
.B1(n_631),
.B2(n_653),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_775),
.Y(n_810)
);

BUFx5_ASAP7_75t_L g811 ( 
.A(n_747),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_770),
.A2(n_601),
.B1(n_578),
.B2(n_572),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_773),
.A2(n_717),
.B1(n_700),
.B2(n_653),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_730),
.B(n_689),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_766),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_735),
.B(n_604),
.C(n_598),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_757),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_740),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_740),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_740),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_728),
.A2(n_564),
.B1(n_542),
.B2(n_667),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_742),
.A2(n_596),
.B1(n_591),
.B2(n_544),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_755),
.Y(n_823)
);

AOI222xp33_ASAP7_75t_L g824 ( 
.A1(n_763),
.A2(n_613),
.B1(n_544),
.B2(n_565),
.C1(n_631),
.C2(n_542),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_768),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_738),
.A2(n_717),
.B1(n_685),
.B2(n_538),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_774),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_771),
.A2(n_520),
.B(n_528),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_761),
.B(n_613),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_741),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_762),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_773),
.A2(n_726),
.B1(n_713),
.B2(n_553),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_759),
.A2(n_700),
.B1(n_546),
.B2(n_620),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_793),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_824),
.A2(n_700),
.B1(n_636),
.B2(n_529),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_782),
.A2(n_636),
.B1(n_537),
.B2(n_600),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_806),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_782),
.A2(n_600),
.B1(n_545),
.B2(n_726),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_786),
.A2(n_713),
.B1(n_620),
.B2(n_685),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_816),
.A2(n_623),
.B1(n_774),
.B2(n_698),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_786),
.A2(n_685),
.B1(n_576),
.B2(n_579),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_SL g842 ( 
.A1(n_779),
.A2(n_623),
.B(n_725),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_785),
.A2(n_685),
.B1(n_579),
.B2(n_576),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_787),
.A2(n_685),
.B1(n_579),
.B2(n_755),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_801),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_784),
.A2(n_685),
.B1(n_579),
.B2(n_755),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_796),
.B(n_725),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_SL g848 ( 
.A1(n_791),
.A2(n_725),
.B(n_566),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_810),
.A2(n_685),
.B1(n_579),
.B2(n_541),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_822),
.A2(n_698),
.B1(n_707),
.B2(n_701),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_803),
.A2(n_584),
.B(n_570),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_809),
.B(n_796),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_783),
.B(n_690),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_810),
.A2(n_541),
.B1(n_649),
.B2(n_723),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_822),
.A2(n_707),
.B1(n_701),
.B2(n_694),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_800),
.A2(n_541),
.B1(n_722),
.B2(n_723),
.Y(n_856)
);

OA21x2_ASAP7_75t_L g857 ( 
.A1(n_828),
.A2(n_781),
.B(n_789),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_795),
.B(n_792),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_799),
.A2(n_707),
.B1(n_701),
.B2(n_694),
.Y(n_859)
);

OAI221xp5_ASAP7_75t_SL g860 ( 
.A1(n_789),
.A2(n_781),
.B1(n_780),
.B2(n_799),
.C(n_812),
.Y(n_860)
);

AOI221xp5_ASAP7_75t_L g861 ( 
.A1(n_809),
.A2(n_696),
.B1(n_692),
.B2(n_723),
.C(n_722),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_794),
.A2(n_541),
.B1(n_722),
.B2(n_692),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_833),
.A2(n_778),
.B1(n_830),
.B2(n_817),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_797),
.A2(n_541),
.B1(n_692),
.B2(n_696),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_797),
.A2(n_696),
.B1(n_692),
.B2(n_664),
.Y(n_865)
);

AOI222xp33_ASAP7_75t_SL g866 ( 
.A1(n_804),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.C1(n_34),
.C2(n_35),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_831),
.A2(n_696),
.B1(n_664),
.B2(n_595),
.Y(n_867)
);

OAI22xp33_ASAP7_75t_SL g868 ( 
.A1(n_807),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_797),
.A2(n_595),
.B1(n_589),
.B2(n_602),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_821),
.A2(n_589),
.B1(n_602),
.B2(n_588),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_797),
.A2(n_599),
.B1(n_571),
.B2(n_605),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_SL g872 ( 
.A1(n_813),
.A2(n_599),
.B(n_140),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_814),
.A2(n_660),
.B1(n_346),
.B2(n_328),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_797),
.A2(n_571),
.B1(n_346),
.B2(n_328),
.Y(n_874)
);

AOI22xp33_ASAP7_75t_L g875 ( 
.A1(n_790),
.A2(n_346),
.B1(n_328),
.B2(n_325),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_790),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_788),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_802),
.B(n_40),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_852),
.B(n_826),
.Y(n_879)
);

OAI21xp33_ASAP7_75t_L g880 ( 
.A1(n_877),
.A2(n_829),
.B(n_805),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_858),
.B(n_837),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_837),
.B(n_825),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_863),
.A2(n_815),
.B1(n_808),
.B2(n_827),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_847),
.B(n_832),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_876),
.A2(n_798),
.B1(n_823),
.B2(n_820),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_834),
.B(n_832),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_836),
.A2(n_819),
.B1(n_818),
.B2(n_811),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_834),
.B(n_811),
.Y(n_888)
);

NAND3xp33_ASAP7_75t_L g889 ( 
.A(n_866),
.B(n_346),
.C(n_325),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_845),
.B(n_811),
.Y(n_890)
);

AOI221xp5_ASAP7_75t_L g891 ( 
.A1(n_868),
.A2(n_346),
.B1(n_325),
.B2(n_61),
.C(n_62),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_SL g892 ( 
.A(n_853),
.B(n_811),
.C(n_59),
.Y(n_892)
);

AND2x2_ASAP7_75t_SL g893 ( 
.A(n_857),
.B(n_811),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_845),
.B(n_811),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_852),
.B(n_58),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_878),
.B(n_64),
.Y(n_896)
);

OAI221xp5_ASAP7_75t_L g897 ( 
.A1(n_835),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.C(n_68),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_839),
.B(n_70),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_857),
.A2(n_71),
.B1(n_74),
.B2(n_75),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_844),
.B(n_76),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_857),
.B(n_846),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_865),
.B(n_79),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_864),
.B(n_80),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_843),
.B(n_82),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_841),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_860),
.B(n_90),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_869),
.B(n_91),
.Y(n_907)
);

OAI221xp5_ASAP7_75t_L g908 ( 
.A1(n_872),
.A2(n_92),
.B1(n_94),
.B2(n_97),
.C(n_98),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_838),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_909)
);

NAND4xp25_ASAP7_75t_SL g910 ( 
.A(n_872),
.B(n_861),
.C(n_862),
.D(n_856),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_842),
.B(n_107),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_908),
.B(n_840),
.C(n_848),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_906),
.B(n_854),
.C(n_849),
.Y(n_913)
);

NAND4xp25_ASAP7_75t_L g914 ( 
.A(n_891),
.B(n_875),
.C(n_871),
.D(n_855),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_881),
.B(n_859),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_895),
.B(n_851),
.C(n_850),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_897),
.B(n_873),
.C(n_867),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_879),
.B(n_874),
.C(n_870),
.Y(n_918)
);

OR2x2_ASAP7_75t_L g919 ( 
.A(n_890),
.B(n_108),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_SL g920 ( 
.A1(n_911),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_884),
.B(n_113),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_888),
.B(n_882),
.Y(n_922)
);

XOR2x2_ASAP7_75t_L g923 ( 
.A(n_885),
.B(n_879),
.Y(n_923)
);

NAND3xp33_ASAP7_75t_L g924 ( 
.A(n_892),
.B(n_114),
.C(n_115),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_909),
.A2(n_119),
.B(n_120),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_894),
.B(n_123),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_SL g927 ( 
.A(n_910),
.B(n_125),
.Y(n_927)
);

NOR2x1_ASAP7_75t_L g928 ( 
.A(n_883),
.B(n_888),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_901),
.B(n_126),
.Y(n_929)
);

OA211x2_ASAP7_75t_L g930 ( 
.A1(n_899),
.A2(n_127),
.B(n_128),
.C(n_129),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_901),
.B(n_130),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_927),
.A2(n_880),
.B1(n_909),
.B2(n_902),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_922),
.Y(n_933)
);

XNOR2xp5_ASAP7_75t_L g934 ( 
.A(n_923),
.B(n_902),
.Y(n_934)
);

XNOR2xp5_ASAP7_75t_L g935 ( 
.A(n_913),
.B(n_903),
.Y(n_935)
);

XOR2x2_ASAP7_75t_L g936 ( 
.A(n_925),
.B(n_896),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_928),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_915),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_929),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_919),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_926),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_921),
.B(n_880),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_931),
.Y(n_943)
);

XNOR2x1_ASAP7_75t_L g944 ( 
.A(n_931),
.B(n_903),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_912),
.B(n_893),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_916),
.Y(n_946)
);

XOR2xp5_ASAP7_75t_L g947 ( 
.A(n_934),
.B(n_935),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_933),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_937),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_938),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_940),
.Y(n_951)
);

XNOR2xp5_ASAP7_75t_L g952 ( 
.A(n_944),
.B(n_920),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_946),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_946),
.Y(n_954)
);

OA22x2_ASAP7_75t_L g955 ( 
.A1(n_947),
.A2(n_945),
.B1(n_932),
.B2(n_943),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_953),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_950),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_952),
.Y(n_958)
);

OA22x2_ASAP7_75t_L g959 ( 
.A1(n_949),
.A2(n_945),
.B1(n_939),
.B2(n_941),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_954),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_953),
.A2(n_942),
.B1(n_936),
.B2(n_954),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_948),
.A2(n_942),
.B1(n_940),
.B2(n_930),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_957),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_956),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_960),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_959),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_961),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_963),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_965),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_964),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_964),
.Y(n_971)
);

AOI22xp5_ASAP7_75t_L g972 ( 
.A1(n_967),
.A2(n_955),
.B1(n_962),
.B2(n_958),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_969),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_SL g974 ( 
.A1(n_970),
.A2(n_966),
.B(n_951),
.C(n_905),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_972),
.A2(n_924),
.B1(n_918),
.B2(n_930),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_968),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_971),
.A2(n_917),
.B(n_914),
.C(n_900),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_975),
.B(n_893),
.Y(n_978)
);

AO22x1_ASAP7_75t_L g979 ( 
.A1(n_973),
.A2(n_904),
.B1(n_907),
.B2(n_898),
.Y(n_979)
);

AO22x2_ASAP7_75t_L g980 ( 
.A1(n_976),
.A2(n_904),
.B1(n_889),
.B2(n_907),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_977),
.B(n_886),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_974),
.B(n_131),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_973),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_973),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_983),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_984),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_980),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_982),
.Y(n_988)
);

INVxp67_ASAP7_75t_SL g989 ( 
.A(n_978),
.Y(n_989)
);

NOR3xp33_ASAP7_75t_L g990 ( 
.A(n_981),
.B(n_132),
.C(n_133),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_979),
.A2(n_887),
.B1(n_136),
.B2(n_138),
.Y(n_991)
);

BUFx4f_ASAP7_75t_SL g992 ( 
.A(n_985),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_987),
.Y(n_993)
);

HB1xp67_ASAP7_75t_L g994 ( 
.A(n_986),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_989),
.A2(n_134),
.B1(n_139),
.B2(n_142),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_988),
.Y(n_996)
);

OR3x2_ASAP7_75t_L g997 ( 
.A(n_990),
.B(n_143),
.C(n_144),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_991),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_989),
.A2(n_145),
.B1(n_147),
.B2(n_153),
.Y(n_999)
);

OAI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_988),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_162),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_994),
.B(n_164),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_993),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_996),
.Y(n_1004)
);

INVxp67_ASAP7_75t_SL g1005 ( 
.A(n_995),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_998),
.B(n_166),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_999),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_997),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1000),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_1003),
.A2(n_167),
.B1(n_168),
.B2(n_173),
.Y(n_1010)
);

AO22x2_ASAP7_75t_L g1011 ( 
.A1(n_1008),
.A2(n_222),
.B1(n_175),
.B2(n_176),
.Y(n_1011)
);

AOI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_1009),
.A2(n_174),
.B1(n_180),
.B2(n_183),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_L g1013 ( 
.A1(n_1004),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1005),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1002),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_1007),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_1011),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_1015),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_1012),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_1016),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_1018),
.A2(n_1006),
.B1(n_1001),
.B2(n_1002),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_1017),
.A2(n_1014),
.B1(n_1010),
.B2(n_1013),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1021),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1022),
.Y(n_1024)
);

OA22x2_ASAP7_75t_L g1025 ( 
.A1(n_1024),
.A2(n_1019),
.B1(n_1020),
.B2(n_202),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1023),
.A2(n_1020),
.B(n_199),
.Y(n_1026)
);

INVxp67_ASAP7_75t_SL g1027 ( 
.A(n_1025),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1026),
.Y(n_1028)
);

AOI221xp5_ASAP7_75t_L g1029 ( 
.A1(n_1027),
.A2(n_196),
.B1(n_204),
.B2(n_209),
.C(n_210),
.Y(n_1029)
);

AOI211xp5_ASAP7_75t_L g1030 ( 
.A1(n_1029),
.A2(n_1028),
.B(n_215),
.C(n_216),
.Y(n_1030)
);


endmodule