module real_jpeg_17613_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_1),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_1),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_1),
.B(n_319),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_2),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_3),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_3),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_4),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_4),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_4),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_4),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_4),
.B(n_366),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_5),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_5),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_5),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_5),
.B(n_183),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_5),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_6),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_6),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_6),
.B(n_34),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_6),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_6),
.B(n_158),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_128),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_6),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_7),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_7),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_7),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_7),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_7),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_7),
.B(n_253),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_7),
.Y(n_360)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_8),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_9),
.Y(n_201)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_9),
.Y(n_326)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_10),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_10),
.Y(n_350)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_11),
.Y(n_75)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_12),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_12),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_12),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_12),
.B(n_31),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_12),
.B(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_13),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_14),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g151 ( 
.A(n_14),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_16),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_16),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_16),
.B(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_113),
.B(n_347),
.C(n_417),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_40),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_24),
.A2(n_25),
.B1(n_67),
.B2(n_77),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_33),
.C(n_37),
.Y(n_25)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_26),
.A2(n_47),
.B1(n_63),
.B2(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_26),
.B(n_190),
.C(n_194),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_26),
.A2(n_47),
.B1(n_190),
.B2(n_191),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

NAND2x1_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_27),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_103),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_27),
.B(n_130),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_27),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_27),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

OR2x2_ASAP7_75t_SL g63 ( 
.A(n_28),
.B(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_32),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_33),
.A2(n_74),
.B(n_76),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_33),
.B(n_74),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_33),
.A2(n_49),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_33),
.B(n_170),
.C(n_173),
.Y(n_214)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_37),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

INVxp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_37),
.B(n_364),
.Y(n_363)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_38),
.Y(n_193)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_78),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_41),
.B(n_78),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_66),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.C(n_56),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_43),
.B(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_44),
.B(n_194),
.C(n_368),
.Y(n_384)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_57),
.C(n_63),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_51),
.B1(n_56),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_54),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_102),
.C(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_63),
.B(n_154),
.C(n_157),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_63),
.A2(n_102),
.B1(n_112),
.B2(n_314),
.Y(n_380)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_68),
.A2(n_69),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_84),
.C(n_89),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_69),
.B(n_76),
.Y(n_417)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_74),
.B(n_218),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_74),
.B(n_187),
.C(n_221),
.Y(n_345)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.C(n_97),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_79),
.B(n_82),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_92),
.C(n_96),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_85),
.B(n_89),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_86),
.B(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_89),
.B(n_198),
.C(n_203),
.Y(n_212)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_90),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_96),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_96),
.A2(n_100),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_96),
.A2(n_100),
.B1(n_347),
.B2(n_351),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_97),
.B(n_405),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.C(n_110),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_98),
.B(n_399),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_100),
.B(n_211),
.C(n_212),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_100),
.B(n_347),
.C(n_394),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_101),
.B(n_110),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_102),
.B(n_259),
.C(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_102),
.A2(n_259),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_102),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_102),
.A2(n_219),
.B1(n_221),
.B2(n_314),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_102),
.Y(n_383)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_106),
.B(n_380),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_108),
.Y(n_292)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_112),
.B(n_282),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_370),
.B(n_411),
.C(n_416),
.Y(n_113)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_274),
.B(n_330),
.C(n_331),
.D(n_369),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_240),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_117),
.B(n_240),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_177),
.Y(n_117)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_118),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_152),
.C(n_167),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_120),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_133),
.C(n_140),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_121),
.B(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_125),
.C(n_129),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_133),
.A2(n_134),
.B1(n_140),
.B2(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_134),
.A2(n_135),
.B(n_137),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_140),
.Y(n_296)
);

MAJx3_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.C(n_148),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_141),
.B(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_143),
.Y(n_367)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_146),
.B(n_148),
.Y(n_248)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_152),
.A2(n_168),
.B1(n_169),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_152),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.C(n_162),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_153),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_154),
.B(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_157),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_160),
.B(n_162),
.Y(n_266)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_166),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_166),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_216),
.B1(n_238),
.B2(n_239),
.Y(n_177)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_207),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_179),
.B(n_213),
.C(n_337),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.C(n_197),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_180),
.B(n_189),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g224 ( 
.A1(n_181),
.A2(n_186),
.B(n_187),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_185),
.A2(n_186),
.B1(n_251),
.B2(n_252),
.Y(n_315)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_187),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_188),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_194),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_194),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_194),
.A2(n_270),
.B1(n_365),
.B2(n_368),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_196),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_197),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_207)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_208),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_216),
.B(n_238),
.C(n_334),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_217),
.B(n_223),
.C(n_226),
.Y(n_341)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_SL g382 ( 
.A(n_221),
.B(n_355),
.C(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_225),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_227)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_233),
.B(n_236),
.C(n_282),
.Y(n_362)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_245),
.C(n_271),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_242),
.B(n_271),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_265),
.C(n_267),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_249),
.C(n_258),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_247),
.B(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_249),
.A2(n_250),
.B1(n_258),
.B2(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx5_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_258),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_259),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_260),
.B(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_267),
.Y(n_278)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_299),
.B(n_329),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_297),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_276),
.B(n_297),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.C(n_293),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_301),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_294),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_283),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.C(n_289),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_310),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.C(n_316),
.Y(n_310)
);

MAJx2_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_321),
.C(n_327),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_320),
.Y(n_359)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_333),
.B(n_335),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_352),
.C(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_352),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_340),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_343),
.C(n_344),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_345),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_347),
.Y(n_351)
);

INVx3_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2x2_ASAP7_75t_SL g352 ( 
.A(n_353),
.B(n_361),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_353),
.B(n_362),
.C(n_363),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_365),
.Y(n_368)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_396),
.C(n_406),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_374),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_372),
.B(n_374),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_375),
.B(n_378),
.C(n_385),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_385),
.B2(n_386),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2x2_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_381),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_382),
.C(n_384),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_395),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_392),
.B2(n_393),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_393),
.C(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_395),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_396),
.A2(n_412),
.B(n_415),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_404),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_404),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.C(n_401),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_400),
.Y(n_409)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_409),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_407),
.A2(n_413),
.B(n_414),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_SL g407 ( 
.A(n_408),
.B(n_410),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_410),
.Y(n_414)
);


endmodule