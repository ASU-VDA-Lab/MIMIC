module fake_aes_1534_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx1_ASAP7_75t_SL g3 ( .A(n_2), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_4), .Y(n_6) );
INVx3_ASAP7_75t_SL g7 ( .A(n_4), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_7), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_8), .B(n_7), .Y(n_10) );
OAI21xp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_9), .B(n_3), .Y(n_11) );
NAND5xp2_ASAP7_75t_L g12 ( .A(n_11), .B(n_0), .C(n_5), .D(n_4), .E(n_7), .Y(n_12) );
AOI21xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B(n_11), .Y(n_13) );
NAND2x1p5_ASAP7_75t_L g14 ( .A(n_13), .B(n_0), .Y(n_14) );
endmodule