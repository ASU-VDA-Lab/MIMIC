module fake_jpeg_22834_n_53 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_53);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_53;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_7),
.B(n_3),
.Y(n_8)
);

INVx6_ASAP7_75t_SL g9 ( 
.A(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_17),
.B(n_21),
.Y(n_25)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_19),
.Y(n_28)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_15),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_10),
.B1(n_13),
.B2(n_15),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_10),
.B1(n_19),
.B2(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_37),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_21),
.C(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.C(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_28),
.B(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_9),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_33),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_32),
.C(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_39),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_44),
.C(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_49),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_11),
.C(n_9),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_2),
.B(n_4),
.Y(n_51)
);

A2O1A1O1Ixp25_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_11),
.B(n_2),
.C(n_5),
.D(n_0),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_0),
.Y(n_53)
);


endmodule