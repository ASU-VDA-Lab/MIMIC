module fake_jpeg_9064_n_280 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_280);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_280;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_35),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_0),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_37),
.B(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_14),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_22),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_53),
.A2(n_24),
.B1(n_14),
.B2(n_17),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_25),
.Y(n_73)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_48),
.B1(n_17),
.B2(n_53),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_15),
.B1(n_34),
.B2(n_31),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_73),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_68),
.B(n_77),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_31),
.C(n_34),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_49),
.C(n_38),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_79),
.A2(n_58),
.B1(n_61),
.B2(n_78),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_91),
.CI(n_96),
.CON(n_110),
.SN(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_82),
.B(n_83),
.Y(n_108)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_30),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_92),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_29),
.C(n_35),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

BUFx4f_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_29),
.C(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_98),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_99),
.A2(n_58),
.B1(n_82),
.B2(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_48),
.B1(n_53),
.B2(n_76),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_103),
.B1(n_109),
.B2(n_111),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_117),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_91),
.A2(n_86),
.B1(n_84),
.B2(n_81),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_121),
.B1(n_27),
.B2(n_25),
.Y(n_142)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_119),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_91),
.A2(n_42),
.B1(n_50),
.B2(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_55),
.B1(n_17),
.B2(n_43),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_113),
.B(n_44),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_46),
.Y(n_116)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_59),
.B1(n_27),
.B2(n_16),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_64),
.B1(n_27),
.B2(n_16),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_135),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_112),
.A2(n_96),
.B(n_94),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_140),
.B(n_143),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_44),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_138),
.C(n_144),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_113),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_117),
.B1(n_119),
.B2(n_64),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_120),
.B(n_97),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_23),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_23),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_141),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_44),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_28),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_104),
.A2(n_25),
.B(n_18),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_145),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_0),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_88),
.Y(n_145)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_1),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_110),
.B(n_114),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_165),
.B(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_139),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_160),
.Y(n_190)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_46),
.B1(n_106),
.B2(n_52),
.Y(n_180)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_110),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_18),
.B(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_9),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_118),
.C(n_106),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_138),
.C(n_129),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_21),
.B(n_118),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_184),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_158),
.A2(n_129),
.B1(n_124),
.B2(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_162),
.B1(n_146),
.B2(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_136),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_182),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_142),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_177),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_166),
.B(n_124),
.C(n_118),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_106),
.C(n_57),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_180),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_70),
.C(n_98),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_70),
.C(n_98),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_189),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_155),
.A2(n_21),
.B(n_67),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_67),
.C(n_46),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

AO22x1_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_163),
.B1(n_160),
.B2(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_198),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_183),
.C(n_169),
.Y(n_218)
);

XOR2x2_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_151),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_196),
.A2(n_210),
.B1(n_176),
.B2(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_179),
.Y(n_198)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_159),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_207),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_153),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_177),
.B(n_146),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_188),
.B1(n_153),
.B2(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_216),
.C(n_222),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_170),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_220),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_178),
.C(n_174),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_223),
.C(n_224),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_147),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_152),
.C(n_181),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_165),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_150),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_194),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_150),
.C(n_173),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_149),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_213),
.B1(n_192),
.B2(n_219),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_232),
.C(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_229),
.B(n_234),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_226),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_231),
.Y(n_246)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_193),
.B(n_203),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_223),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_221),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_201),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_7),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_8),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g240 ( 
.A1(n_221),
.A2(n_214),
.A3(n_173),
.B1(n_19),
.B2(n_28),
.C1(n_21),
.C2(n_6),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_19),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_245),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_8),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_249),
.B(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_252),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_19),
.C(n_28),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_19),
.C(n_28),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_1),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_7),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_241),
.B(n_7),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_8),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_237),
.B(n_232),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_259),
.B(n_260),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_246),
.A2(n_241),
.B(n_235),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_6),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_251),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_265),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_6),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_261),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_10),
.B(n_11),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_254),
.B(n_9),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_269),
.A2(n_272),
.B(n_11),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_270),
.A2(n_264),
.B1(n_13),
.B2(n_3),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_274),
.B(n_271),
.Y(n_275)
);

OAI311xp33_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_13),
.A3(n_2),
.B1(n_3),
.C1(n_4),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_276),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_1),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_278),
.A2(n_2),
.B(n_3),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_2),
.Y(n_280)
);


endmodule