module fake_jpeg_7120_n_37 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_6),
.B(n_5),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_5),
.B(n_3),
.C(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_21),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_4),
.B(n_10),
.C(n_14),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_29)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_13),
.Y(n_27)
);

AOI322xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_12),
.A3(n_13),
.B1(n_16),
.B2(n_17),
.C1(n_20),
.C2(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_20),
.B1(n_22),
.B2(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_29),
.B(n_24),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_23),
.C(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_34),
.Y(n_37)
);


endmodule