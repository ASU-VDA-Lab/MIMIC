module fake_jpeg_13166_n_30 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_30);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_30;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_29;
wire n_12;
wire n_15;

BUFx4f_ASAP7_75t_SL g10 ( 
.A(n_9),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_9),
.B(n_1),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g16 ( 
.A(n_14),
.B(n_1),
.C(n_2),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_11),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_12),
.B1(n_11),
.B2(n_13),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_20),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_10),
.B(n_17),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_10),
.C(n_4),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_23),
.C(n_5),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_3),
.Y(n_27)
);

AOI321xp33_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C(n_23),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_6),
.B(n_10),
.Y(n_30)
);


endmodule