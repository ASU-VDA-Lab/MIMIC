module fake_jpeg_19196_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_0),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_0),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_57),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_55),
.B1(n_56),
.B2(n_46),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_57),
.B1(n_45),
.B2(n_63),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_44),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_64),
.B1(n_50),
.B2(n_49),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_84),
.A2(n_85),
.B1(n_42),
.B2(n_53),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_64),
.B1(n_61),
.B2(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_86),
.Y(n_91)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_97),
.B1(n_99),
.B2(n_62),
.Y(n_101)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_59),
.C(n_60),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_109),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_47),
.B(n_52),
.C(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_110),
.Y(n_126)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_114),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_90),
.B(n_99),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_112),
.B(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_96),
.B(n_47),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g113 ( 
.A1(n_91),
.A2(n_2),
.B(n_3),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_5),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_66),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_43),
.C(n_68),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_101),
.C(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_120),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_104),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_10),
.B(n_13),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_14),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_123),
.B(n_111),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_128),
.A2(n_129),
.B(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

INVx13_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_119),
.B1(n_132),
.B2(n_126),
.Y(n_136)
);

AO221x1_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_128),
.B1(n_124),
.B2(n_133),
.C(n_117),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_130),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_135),
.B1(n_19),
.B2(n_25),
.Y(n_139)
);

INVxp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_102),
.B(n_26),
.Y(n_141)
);

AOI21x1_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_17),
.B(n_28),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_143),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_33),
.Y(n_146)
);


endmodule