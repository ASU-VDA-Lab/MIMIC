module fake_jpeg_3610_n_95 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_0),
.Y(n_54)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_1),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_40),
.B1(n_37),
.B2(n_36),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_35),
.B1(n_34),
.B2(n_28),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_27),
.B(n_30),
.C(n_31),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_48),
.B(n_35),
.C(n_4),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_36),
.C(n_30),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_55),
.C(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_35),
.C(n_28),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_1),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_47),
.B(n_14),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_57),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_47),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_12),
.B1(n_24),
.B2(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_68),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_2),
.B(n_3),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_49),
.B1(n_3),
.B2(n_5),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_77),
.B(n_78),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_11),
.C(n_21),
.Y(n_75)
);

A2O1A1O1Ixp25_ASAP7_75t_L g85 ( 
.A1(n_75),
.A2(n_78),
.B(n_9),
.C(n_18),
.D(n_19),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_10),
.C(n_20),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_76),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_87),
.C(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

OAI31xp33_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_82),
.A3(n_86),
.B(n_72),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_70),
.C(n_81),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_81),
.B(n_75),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_85),
.B1(n_25),
.B2(n_7),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_2),
.Y(n_95)
);


endmodule