module fake_jpeg_1512_n_26 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_7),
.A2(n_5),
.B1(n_0),
.B2(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_2),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_9),
.A2(n_4),
.B1(n_6),
.B2(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_19),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_9),
.A2(n_2),
.B(n_4),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_6),
.Y(n_18)
);

OAI22x1_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_10),
.B1(n_8),
.B2(n_12),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_SL g23 ( 
.A(n_22),
.B(n_19),
.C(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_20),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_25),
.B(n_24),
.Y(n_26)
);


endmodule