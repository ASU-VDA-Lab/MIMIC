module real_aes_15848_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_239;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1346;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_238;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_246;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_247;
wire n_264;
wire n_237;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_235;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_245;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_248;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_249;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_243;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1343;
wire n_719;
wire n_465;
wire n_1156;
wire n_988;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_241;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_236;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_244;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_314;
wire n_283;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_240;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_0), .A2(n_175), .B1(n_1111), .B2(n_1115), .Y(n_1167) );
AOI22xp33_ASAP7_75t_SL g813 ( .A1(n_1), .A2(n_65), .B1(n_808), .B2(n_809), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_1), .A2(n_213), .B1(n_644), .B2(n_647), .Y(n_825) );
INVx1_ASAP7_75t_L g819 ( .A(n_2), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_3), .A2(n_106), .B1(n_619), .B2(n_621), .Y(n_618) );
AOI22xp33_ASAP7_75t_SL g643 ( .A1(n_3), .A2(n_110), .B1(n_644), .B2(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_4), .A2(n_48), .B1(n_1111), .B2(n_1115), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_5), .A2(n_67), .B1(n_809), .B2(n_1064), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_5), .A2(n_47), .B1(n_1083), .B2(n_1084), .Y(n_1082) );
INVx1_ASAP7_75t_L g248 ( .A(n_6), .Y(n_248) );
AND2x2_ASAP7_75t_L g269 ( .A(n_6), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_6), .B(n_196), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_6), .B(n_258), .Y(n_580) );
INVx1_ASAP7_75t_L g685 ( .A(n_7), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g810 ( .A1(n_8), .A2(n_130), .B1(n_805), .B2(n_811), .C(n_812), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_8), .A2(n_57), .B1(n_647), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g615 ( .A1(n_9), .A2(n_143), .B1(n_616), .B2(n_617), .Y(n_615) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_9), .A2(n_14), .B1(n_328), .B2(n_637), .C(n_639), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g1014 ( .A1(n_10), .A2(n_117), .B1(n_402), .B2(n_863), .Y(n_1014) );
INVxp67_ASAP7_75t_SL g1041 ( .A(n_10), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_11), .A2(n_133), .B1(n_303), .B2(n_306), .Y(n_302) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_11), .A2(n_217), .B1(n_402), .B2(n_426), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g801 ( .A(n_12), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_13), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g625 ( .A1(n_14), .A2(n_30), .B1(n_460), .B2(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g1114 ( .A(n_15), .Y(n_1114) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_15), .B(n_93), .Y(n_1116) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_15), .B(n_1120), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1019 ( .A1(n_16), .A2(n_208), .B1(n_863), .B2(n_1020), .Y(n_1019) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_16), .A2(n_117), .B1(n_637), .B2(n_1031), .C(n_1032), .Y(n_1030) );
INVx1_ASAP7_75t_L g613 ( .A(n_17), .Y(n_613) );
OAI22xp33_ASAP7_75t_L g627 ( .A1(n_18), .A2(n_184), .B1(n_477), .B2(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g652 ( .A(n_18), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_19), .A2(n_29), .B1(n_1118), .B2(n_1121), .Y(n_1144) );
XNOR2xp5_ASAP7_75t_L g902 ( .A(n_20), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g876 ( .A(n_21), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_22), .A2(n_201), .B1(n_362), .B2(n_373), .Y(n_1026) );
XOR2x2_ASAP7_75t_L g672 ( .A(n_23), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g286 ( .A(n_24), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_24), .A2(n_206), .B1(n_362), .B2(n_373), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_25), .A2(n_104), .B1(n_1118), .B2(n_1121), .Y(n_1166) );
INVx1_ASAP7_75t_L g1323 ( .A(n_26), .Y(n_1323) );
OAI22xp33_ASAP7_75t_L g1340 ( .A1(n_26), .A2(n_153), .B1(n_435), .B2(n_628), .Y(n_1340) );
OAI221xp5_ASAP7_75t_L g1330 ( .A1(n_27), .A2(n_52), .B1(n_491), .B2(n_492), .C(n_1331), .Y(n_1330) );
INVx1_ASAP7_75t_L g1349 ( .A(n_27), .Y(n_1349) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_28), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g655 ( .A1(n_30), .A2(n_656), .B(n_657), .C(n_666), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g969 ( .A(n_31), .B(n_970), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_31), .A2(n_144), .B1(n_863), .B2(n_994), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_32), .A2(n_86), .B1(n_1111), .B2(n_1205), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_33), .A2(n_144), .B1(n_288), .B2(n_305), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_33), .A2(n_210), .B1(n_626), .B2(n_863), .Y(n_989) );
INVx1_ASAP7_75t_L g700 ( .A(n_34), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g1141 ( .A1(n_35), .A2(n_81), .B1(n_1111), .B2(n_1132), .Y(n_1141) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_36), .A2(n_54), .B1(n_362), .B2(n_454), .Y(n_632) );
OAI211xp5_ASAP7_75t_L g634 ( .A1(n_36), .A2(n_480), .B(n_635), .C(n_648), .Y(n_634) );
XNOR2x2_ASAP7_75t_L g606 ( .A(n_37), .B(n_607), .Y(n_606) );
AOI21xp33_ASAP7_75t_L g918 ( .A1(n_38), .A2(n_573), .B(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g928 ( .A(n_38), .Y(n_928) );
XOR2x2_ASAP7_75t_L g1006 ( .A(n_39), .B(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_SL g1068 ( .A1(n_40), .A2(n_116), .B1(n_458), .B2(n_868), .Y(n_1068) );
INVxp67_ASAP7_75t_SL g1098 ( .A(n_40), .Y(n_1098) );
INVx1_ASAP7_75t_L g475 ( .A(n_41), .Y(n_475) );
INVx1_ASAP7_75t_L g349 ( .A(n_42), .Y(n_349) );
INVx1_ASAP7_75t_L g379 ( .A(n_42), .Y(n_379) );
INVx1_ASAP7_75t_L g952 ( .A(n_43), .Y(n_952) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_44), .A2(n_174), .B1(n_644), .B2(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g929 ( .A(n_44), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_45), .A2(n_156), .B1(n_477), .B2(n_628), .Y(n_1022) );
INVx1_ASAP7_75t_L g1035 ( .A(n_45), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1131 ( .A1(n_46), .A2(n_112), .B1(n_1111), .B2(n_1132), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_47), .A2(n_124), .B1(n_809), .B2(n_1066), .Y(n_1065) );
INVxp67_ASAP7_75t_SL g1314 ( .A(n_48), .Y(n_1314) );
AND4x1_ASAP7_75t_L g1351 ( .A(n_48), .B(n_1316), .C(n_1319), .D(n_1338), .Y(n_1351) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_48), .A2(n_1359), .B1(n_1361), .B2(n_1365), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_49), .A2(n_195), .B1(n_1118), .B2(n_1121), .Y(n_1206) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_50), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g416 ( .A1(n_50), .A2(n_115), .B1(n_417), .B2(n_419), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_51), .A2(n_110), .B1(n_621), .B2(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_51), .A2(n_106), .B1(n_659), .B2(n_662), .C(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g1350 ( .A(n_52), .Y(n_1350) );
INVx1_ASAP7_75t_L g241 ( .A(n_53), .Y(n_241) );
INVx2_ASAP7_75t_L g355 ( .A(n_55), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g907 ( .A1(n_56), .A2(n_200), .B1(n_328), .B2(n_572), .C(n_908), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_56), .A2(n_229), .B1(n_402), .B2(n_442), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_57), .A2(n_63), .B1(n_460), .B2(n_805), .C(n_806), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_58), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g393 ( .A(n_58), .Y(n_393) );
INVx1_ASAP7_75t_L g1071 ( .A(n_59), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_60), .A2(n_72), .B1(n_463), .B2(n_466), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_60), .A2(n_199), .B1(n_303), .B2(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g796 ( .A(n_61), .Y(n_796) );
INVx1_ASAP7_75t_L g795 ( .A(n_62), .Y(n_795) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_63), .A2(n_130), .B1(n_638), .B2(n_641), .C(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g996 ( .A(n_64), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g830 ( .A1(n_65), .A2(n_69), .B1(n_572), .B2(n_641), .C(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_SL g860 ( .A1(n_66), .A2(n_164), .B1(n_861), .B2(n_863), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g895 ( .A1(n_66), .A2(n_202), .B1(n_644), .B2(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g1095 ( .A(n_67), .Y(n_1095) );
INVx1_ASAP7_75t_L g558 ( .A(n_68), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_68), .A2(n_111), .B1(n_572), .B2(n_573), .C(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_69), .A2(n_213), .B1(n_808), .B2(n_809), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_70), .A2(n_182), .B1(n_362), .B2(n_373), .Y(n_1318) );
OAI211xp5_ASAP7_75t_L g1320 ( .A1(n_70), .A2(n_480), .B(n_1321), .C(n_1324), .Y(n_1320) );
AOI22xp5_ASAP7_75t_L g1117 ( .A1(n_71), .A2(n_105), .B1(n_1118), .B2(n_1121), .Y(n_1117) );
AOI21xp33_ASAP7_75t_L g499 ( .A1(n_72), .A2(n_310), .B(n_312), .Y(n_499) );
OAI211xp5_ASAP7_75t_L g737 ( .A1(n_73), .A2(n_719), .B(n_738), .C(n_740), .Y(n_737) );
INVx1_ASAP7_75t_L g783 ( .A(n_73), .Y(n_783) );
OAI22xp5_ASAP7_75t_SL g965 ( .A1(n_74), .A2(n_91), .B1(n_678), .B2(n_691), .Y(n_965) );
OAI21xp33_ASAP7_75t_L g976 ( .A1(n_74), .A2(n_977), .B(n_978), .Y(n_976) );
INVx1_ASAP7_75t_L g1057 ( .A(n_75), .Y(n_1057) );
OAI222xp33_ASAP7_75t_L g1087 ( .A1(n_75), .A2(n_108), .B1(n_492), .B2(n_1088), .C1(n_1089), .C2(n_1096), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g1152 ( .A1(n_76), .A2(n_96), .B1(n_1111), .B2(n_1115), .Y(n_1152) );
INVx1_ASAP7_75t_L g1012 ( .A(n_77), .Y(n_1012) );
OAI221xp5_ASAP7_75t_L g1037 ( .A1(n_77), .A2(n_83), .B1(n_292), .B2(n_491), .C(n_1038), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g476 ( .A1(n_78), .A2(n_80), .B1(n_429), .B2(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g488 ( .A(n_78), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_79), .A2(n_221), .B1(n_457), .B2(n_460), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g500 ( .A1(n_79), .A2(n_155), .B1(n_501), .B2(n_502), .Y(n_500) );
INVx1_ASAP7_75t_L g489 ( .A(n_80), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_82), .A2(n_226), .B1(n_896), .B2(n_1329), .Y(n_1328) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_82), .A2(n_101), .B1(n_419), .B2(n_1344), .Y(n_1345) );
INVx1_ASAP7_75t_L g1011 ( .A(n_83), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_84), .Y(n_243) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_84), .B(n_241), .Y(n_1112) );
AOI22xp33_ASAP7_75t_SL g864 ( .A1(n_85), .A2(n_233), .B1(n_417), .B2(n_865), .Y(n_864) );
AOI21xp33_ASAP7_75t_L g892 ( .A1(n_85), .A2(n_831), .B(n_893), .Y(n_892) );
CKINVDCx5p33_ASAP7_75t_R g799 ( .A(n_87), .Y(n_799) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_88), .Y(n_917) );
OAI211xp5_ASAP7_75t_L g955 ( .A1(n_89), .A2(n_956), .B(n_958), .C(n_959), .Y(n_955) );
INVxp33_ASAP7_75t_SL g979 ( .A(n_89), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_90), .A2(n_218), .B1(n_429), .B2(n_477), .Y(n_877) );
INVx1_ASAP7_75t_L g885 ( .A(n_90), .Y(n_885) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_91), .Y(n_1000) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_92), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_93), .B(n_1114), .Y(n_1113) );
INVx1_ASAP7_75t_L g1120 ( .A(n_93), .Y(n_1120) );
INVxp67_ASAP7_75t_SL g1334 ( .A(n_94), .Y(n_1334) );
AOI22xp33_ASAP7_75t_SL g1346 ( .A1(n_94), .A2(n_183), .B1(n_426), .B2(n_1347), .Y(n_1346) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_95), .A2(n_151), .B1(n_1118), .B2(n_1121), .Y(n_1130) );
CKINVDCx5p33_ASAP7_75t_R g1317 ( .A(n_97), .Y(n_1317) );
INVx1_ASAP7_75t_L g746 ( .A(n_98), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g776 ( .A1(n_98), .A2(n_682), .B(n_777), .C(n_780), .Y(n_776) );
INVxp67_ASAP7_75t_SL g317 ( .A(n_99), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_99), .A2(n_216), .B1(n_409), .B2(n_413), .Y(n_408) );
OAI211xp5_ASAP7_75t_SL g291 ( .A1(n_100), .A2(n_292), .B(n_297), .C(n_314), .Y(n_291) );
INVx1_ASAP7_75t_L g388 ( .A(n_100), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g1335 ( .A1(n_101), .A2(n_190), .B1(n_483), .B2(n_831), .C(n_1336), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_102), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g383 ( .A(n_102), .Y(n_383) );
INVx1_ASAP7_75t_L g424 ( .A(n_102), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_103), .A2(n_135), .B1(n_415), .B2(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g583 ( .A(n_103), .Y(n_583) );
INVx1_ASAP7_75t_L g280 ( .A(n_107), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_107), .A2(n_227), .B1(n_429), .B2(n_435), .Y(n_428) );
INVx1_ASAP7_75t_L g1056 ( .A(n_108), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_109), .A2(n_204), .B1(n_1118), .B2(n_1121), .Y(n_1153) );
AOI221xp5_ASAP7_75t_L g547 ( .A1(n_111), .A2(n_211), .B1(n_405), .B2(n_548), .C(n_549), .Y(n_547) );
XNOR2xp5_ASAP7_75t_L g512 ( .A(n_112), .B(n_513), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g1110 ( .A1(n_113), .A2(n_114), .B1(n_1111), .B2(n_1115), .Y(n_1110) );
INVxp67_ASAP7_75t_SL g298 ( .A(n_115), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g1077 ( .A1(n_116), .A2(n_224), .B1(n_1078), .B2(n_1079), .C(n_1081), .Y(n_1077) );
INVx1_ASAP7_75t_L g677 ( .A(n_118), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_119), .A2(n_199), .B1(n_466), .B2(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g495 ( .A(n_119), .Y(n_495) );
INVx1_ASAP7_75t_L g699 ( .A(n_120), .Y(n_699) );
INVx1_ASAP7_75t_L g914 ( .A(n_121), .Y(n_914) );
INVxp67_ASAP7_75t_SL g858 ( .A(n_122), .Y(n_858) );
OAI211xp5_ASAP7_75t_L g879 ( .A1(n_122), .A2(n_880), .B(n_881), .C(n_884), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g866 ( .A1(n_123), .A2(n_214), .B1(n_417), .B2(n_865), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_123), .A2(n_233), .B1(n_501), .B2(n_647), .Y(n_883) );
INVx1_ASAP7_75t_L g1091 ( .A(n_124), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_125), .A2(n_128), .B1(n_1118), .B2(n_1121), .Y(n_1134) );
XOR2xp5_ASAP7_75t_L g1362 ( .A(n_126), .B(n_1363), .Y(n_1362) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_127), .A2(n_225), .B1(n_525), .B2(n_528), .Y(n_524) );
INVxp33_ASAP7_75t_SL g602 ( .A(n_127), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_129), .A2(n_229), .B1(n_288), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g938 ( .A1(n_129), .A2(n_200), .B1(n_402), .B2(n_811), .Y(n_938) );
INVx1_ASAP7_75t_L g913 ( .A(n_131), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_132), .A2(n_223), .B1(n_419), .B2(n_1016), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_132), .A2(n_169), .B1(n_646), .B2(n_921), .Y(n_1033) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_133), .A2(n_158), .B1(n_402), .B2(n_404), .Y(n_401) );
BUFx3_ASAP7_75t_L g348 ( .A(n_134), .Y(n_348) );
INVx1_ASAP7_75t_L g575 ( .A(n_135), .Y(n_575) );
INVx1_ASAP7_75t_L g853 ( .A(n_136), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g887 ( .A1(n_136), .A2(n_137), .B1(n_331), .B2(n_493), .C(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g856 ( .A(n_137), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_138), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_139), .A2(n_202), .B1(n_863), .B2(n_868), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g882 ( .A1(n_139), .A2(n_164), .B1(n_328), .B2(n_573), .C(n_638), .Y(n_882) );
AOI22xp5_ASAP7_75t_L g1142 ( .A1(n_140), .A2(n_142), .B1(n_1118), .B2(n_1121), .Y(n_1142) );
INVx1_ASAP7_75t_L g544 ( .A(n_141), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_141), .A2(n_173), .B1(n_572), .B2(n_573), .C(n_574), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_143), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_L g444 ( .A(n_145), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g1145 ( .A1(n_145), .A2(n_198), .B1(n_1111), .B2(n_1115), .Y(n_1145) );
OAI21xp33_ASAP7_75t_L g1069 ( .A1(n_146), .A2(n_362), .B(n_1070), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_147), .A2(n_155), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_147), .A2(n_221), .B1(n_327), .B2(n_328), .C(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_148), .Y(n_255) );
INVx1_ASAP7_75t_L g517 ( .A(n_149), .Y(n_517) );
INVx1_ASAP7_75t_L g820 ( .A(n_150), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_152), .Y(n_536) );
INVx1_ASAP7_75t_L g1322 ( .A(n_153), .Y(n_1322) );
OAI21xp5_ASAP7_75t_SL g834 ( .A1(n_154), .A2(n_835), .B(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g1036 ( .A(n_156), .Y(n_1036) );
INVx1_ASAP7_75t_L g555 ( .A(n_157), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_158), .A2(n_217), .B1(n_325), .B2(n_327), .C(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g1072 ( .A(n_159), .Y(n_1072) );
INVx1_ASAP7_75t_L g449 ( .A(n_160), .Y(n_449) );
OAI221xp5_ASAP7_75t_SL g490 ( .A1(n_160), .A2(n_219), .B1(n_491), .B2(n_492), .C(n_494), .Y(n_490) );
XOR2x2_ASAP7_75t_L g262 ( .A(n_161), .B(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g1060 ( .A(n_162), .Y(n_1060) );
INVx1_ASAP7_75t_L g693 ( .A(n_163), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g750 ( .A1(n_165), .A2(n_180), .B1(n_751), .B2(n_754), .Y(n_750) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_165), .A2(n_180), .B1(n_763), .B2(n_764), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g915 ( .A1(n_166), .A2(n_203), .B1(n_331), .B2(n_493), .C(n_916), .Y(n_915) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_166), .A2(n_203), .B1(n_855), .B2(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g680 ( .A(n_167), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g973 ( .A1(n_168), .A2(n_312), .B(n_573), .Y(n_973) );
INVx1_ASAP7_75t_L g987 ( .A(n_168), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_169), .A2(n_232), .B1(n_419), .B2(n_1016), .Y(n_1015) );
INVxp67_ASAP7_75t_SL g1332 ( .A(n_170), .Y(n_1332) );
AOI22xp33_ASAP7_75t_SL g1342 ( .A1(n_170), .A2(n_189), .B1(n_404), .B2(n_626), .Y(n_1342) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_171), .Y(n_254) );
INVx1_ASAP7_75t_L g741 ( .A(n_172), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g561 ( .A1(n_173), .A2(n_410), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g937 ( .A(n_174), .Y(n_937) );
XOR2x2_ASAP7_75t_L g947 ( .A(n_175), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g360 ( .A(n_176), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_177), .Y(n_631) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_178), .A2(n_215), .B1(n_288), .B2(n_829), .Y(n_968) );
INVx1_ASAP7_75t_L g988 ( .A(n_178), .Y(n_988) );
INVx1_ASAP7_75t_L g688 ( .A(n_179), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_181), .B(n_849), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g872 ( .A1(n_181), .A2(n_873), .B1(n_874), .B2(n_897), .Y(n_872) );
INVx1_ASAP7_75t_L g899 ( .A(n_181), .Y(n_899) );
AOI221xp5_ASAP7_75t_L g1325 ( .A1(n_183), .A2(n_189), .B1(n_325), .B2(n_1081), .C(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g649 ( .A(n_184), .Y(n_649) );
INVx1_ASAP7_75t_L g694 ( .A(n_185), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_186), .A2(n_197), .B1(n_729), .B2(n_733), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g767 ( .A1(n_186), .A2(n_197), .B1(n_768), .B2(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g611 ( .A(n_187), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_188), .A2(n_230), .B1(n_373), .B2(n_835), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_190), .A2(n_226), .B1(n_419), .B2(n_1344), .Y(n_1343) );
AOI22xp33_ASAP7_75t_SL g1062 ( .A1(n_191), .A2(n_224), .B1(n_811), .B2(n_861), .Y(n_1062) );
INVxp67_ASAP7_75t_SL g1097 ( .A(n_191), .Y(n_1097) );
OAI211xp5_ASAP7_75t_SL g530 ( .A1(n_192), .A2(n_531), .B(n_533), .C(n_538), .Y(n_530) );
INVx1_ASAP7_75t_L g588 ( .A(n_192), .Y(n_588) );
INVx1_ASAP7_75t_L g942 ( .A(n_193), .Y(n_942) );
CKINVDCx5p33_ASAP7_75t_R g961 ( .A(n_194), .Y(n_961) );
BUFx3_ASAP7_75t_L g258 ( .A(n_196), .Y(n_258) );
INVx1_ASAP7_75t_L g270 ( .A(n_196), .Y(n_270) );
OAI211xp5_ASAP7_75t_L g1028 ( .A1(n_201), .A2(n_880), .B(n_1029), .C(n_1034), .Y(n_1028) );
INVx2_ASAP7_75t_L g340 ( .A(n_205), .Y(n_340) );
INVx1_ASAP7_75t_L g353 ( .A(n_205), .Y(n_353) );
INVx1_ASAP7_75t_L g358 ( .A(n_205), .Y(n_358) );
XNOR2x1_ASAP7_75t_L g791 ( .A(n_207), .B(n_792), .Y(n_791) );
INVxp67_ASAP7_75t_SL g1044 ( .A(n_208), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_209), .Y(n_1025) );
NAND2xp5_ASAP7_75t_SL g967 ( .A(n_210), .B(n_573), .Y(n_967) );
INVx1_ASAP7_75t_L g576 ( .A(n_211), .Y(n_576) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_212), .Y(n_452) );
OAI211xp5_ASAP7_75t_SL g479 ( .A1(n_212), .A2(n_480), .B(n_481), .C(n_487), .Y(n_479) );
INVx1_ASAP7_75t_L g889 ( .A(n_214), .Y(n_889) );
INVxp67_ASAP7_75t_SL g992 ( .A(n_215), .Y(n_992) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_216), .A2(n_308), .B(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g886 ( .A(n_218), .Y(n_886) );
INVx1_ASAP7_75t_L g450 ( .A(n_219), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g546 ( .A(n_220), .Y(n_546) );
INVx1_ASAP7_75t_L g1100 ( .A(n_222), .Y(n_1100) );
AOI221xp5_ASAP7_75t_L g1045 ( .A1(n_223), .A2(n_232), .B1(n_831), .B2(n_1046), .C(n_1047), .Y(n_1045) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_225), .Y(n_522) );
INVx1_ASAP7_75t_L g274 ( .A(n_227), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g960 ( .A(n_228), .Y(n_960) );
OAI211xp5_ASAP7_75t_L g905 ( .A1(n_230), .A2(n_880), .B(n_906), .C(n_912), .Y(n_905) );
INVx1_ASAP7_75t_L g972 ( .A(n_231), .Y(n_972) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_259), .B(n_1104), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_244), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_238), .B(n_247), .Y(n_1357) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_242), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g1360 ( .A(n_240), .B(n_243), .Y(n_1360) );
INVx1_ASAP7_75t_L g1366 ( .A(n_240), .Y(n_1366) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g1368 ( .A(n_243), .B(n_1366), .Y(n_1368) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x4_ASAP7_75t_L g788 ( .A(n_247), .B(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g313 ( .A(n_248), .B(n_257), .Y(n_313) );
AND2x4_ASAP7_75t_L g329 ( .A(n_248), .B(n_258), .Y(n_329) );
INVx1_ASAP7_75t_L g763 ( .A(n_249), .Y(n_763) );
AND2x4_ASAP7_75t_SL g1356 ( .A(n_249), .B(n_1357), .Y(n_1356) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVxp67_ASAP7_75t_L g665 ( .A(n_251), .Y(n_665) );
OR2x6_ASAP7_75t_L g769 ( .A(n_251), .B(n_766), .Y(n_769) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_L g316 ( .A(n_252), .Y(n_316) );
BUFx4f_ASAP7_75t_L g957 ( .A(n_252), .Y(n_957) );
INVx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g272 ( .A(n_254), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g277 ( .A(n_254), .B(n_255), .Y(n_277) );
INVx2_ASAP7_75t_L g284 ( .A(n_254), .Y(n_284) );
INVx2_ASAP7_75t_L g290 ( .A(n_254), .Y(n_290) );
NAND2x1_ASAP7_75t_L g301 ( .A(n_254), .B(n_255), .Y(n_301) );
INVx1_ASAP7_75t_L g366 ( .A(n_254), .Y(n_366) );
INVx2_ASAP7_75t_L g273 ( .A(n_255), .Y(n_273) );
INVx1_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
AND2x2_ASAP7_75t_L g289 ( .A(n_255), .B(n_290), .Y(n_289) );
BUFx2_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_255), .B(n_290), .Y(n_322) );
OR2x2_ASAP7_75t_L g679 ( .A(n_255), .B(n_284), .Y(n_679) );
INVxp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g779 ( .A(n_257), .Y(n_779) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
BUFx2_ASAP7_75t_L g775 ( .A(n_258), .Y(n_775) );
AND2x4_ASAP7_75t_L g786 ( .A(n_258), .B(n_365), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_842), .B1(n_1102), .B2(n_1103), .Y(n_259) );
INVx1_ASAP7_75t_L g1102 ( .A(n_260), .Y(n_1102) );
XNOR2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_508), .Y(n_260) );
XNOR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_443), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_341), .C(n_385), .Y(n_263) );
OAI31xp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_291), .A3(n_330), .B(n_335), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_279), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_274), .B(n_275), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_267), .A2(n_281), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_267), .A2(n_650), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1321 ( .A1(n_267), .A2(n_281), .B1(n_1322), .B2(n_1323), .Y(n_1321) );
BUFx6f_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g654 ( .A(n_268), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g818 ( .A1(n_268), .A2(n_281), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_268), .A2(n_281), .B1(n_885), .B2(n_886), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_268), .A2(n_282), .B1(n_913), .B2(n_914), .Y(n_912) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_268), .A2(n_650), .B1(n_1071), .B2(n_1072), .Y(n_1075) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
AND2x2_ASAP7_75t_L g282 ( .A(n_269), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g287 ( .A(n_269), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_SL g334 ( .A(n_269), .B(n_276), .Y(n_334) );
AND2x2_ASAP7_75t_L g521 ( .A(n_269), .B(n_271), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_269), .B(n_358), .Y(n_570) );
AND2x2_ASAP7_75t_L g822 ( .A(n_269), .B(n_485), .Y(n_822) );
BUFx2_ASAP7_75t_L g964 ( .A(n_269), .Y(n_964) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_270), .Y(n_766) );
INVx2_ASAP7_75t_L g642 ( .A(n_271), .Y(n_642) );
INVx1_ASAP7_75t_L g909 ( .A(n_271), .Y(n_909) );
BUFx6f_ASAP7_75t_L g1080 ( .A(n_271), .Y(n_1080) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g311 ( .A(n_272), .Y(n_311) );
BUFx3_ASAP7_75t_L g573 ( .A(n_272), .Y(n_573) );
AND2x4_ASAP7_75t_L g765 ( .A(n_272), .B(n_766), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_275), .A2(n_482), .B(n_484), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_275), .A2(n_636), .B(n_643), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_275), .A2(n_795), .B1(n_822), .B2(n_823), .C(n_825), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_275), .A2(n_882), .B(n_883), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g906 ( .A1(n_275), .A2(n_907), .B(n_910), .Y(n_906) );
AOI21xp5_ASAP7_75t_SL g1029 ( .A1(n_275), .A2(n_1030), .B(n_1033), .Y(n_1029) );
AOI21xp5_ASAP7_75t_L g1076 ( .A1(n_275), .A2(n_1077), .B(n_1082), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1324 ( .A1(n_275), .A2(n_1325), .B(n_1328), .Y(n_1324) );
AND2x6_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
BUFx3_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
BUFx3_ASAP7_75t_L g572 ( .A(n_276), .Y(n_572) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_276), .Y(n_638) );
AND2x2_ASAP7_75t_L g778 ( .A(n_276), .B(n_779), .Y(n_778) );
BUFx3_ASAP7_75t_L g970 ( .A(n_276), .Y(n_970) );
BUFx3_ASAP7_75t_L g1046 ( .A(n_276), .Y(n_1046) );
INVx1_ASAP7_75t_L g1327 ( .A(n_276), .Y(n_1327) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g661 ( .A(n_277), .Y(n_661) );
INVx1_ASAP7_75t_L g296 ( .A(n_278), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_278), .B(n_283), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_278), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_278), .B(n_340), .Y(n_594) );
AND2x2_ASAP7_75t_L g832 ( .A(n_278), .B(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_281), .B1(n_286), .B2(n_287), .Y(n_279) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g515 ( .A(n_282), .B(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g651 ( .A(n_282), .Y(n_651) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_283), .Y(n_305) );
INVx3_ASAP7_75t_L g645 ( .A(n_283), .Y(n_645) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
HB1xp67_ASAP7_75t_L g963 ( .A(n_284), .Y(n_963) );
INVx3_ASAP7_75t_L g480 ( .A(n_287), .Y(n_480) );
INVx2_ASAP7_75t_SL g880 ( .A(n_287), .Y(n_880) );
NAND2xp5_ASAP7_75t_R g1086 ( .A(n_287), .B(n_1060), .Y(n_1086) );
BUFx2_ASAP7_75t_L g306 ( .A(n_288), .Y(n_306) );
INVx1_ASAP7_75t_L g503 ( .A(n_288), .Y(n_503) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g486 ( .A(n_289), .Y(n_486) );
BUFx3_ASAP7_75t_L g647 ( .A(n_289), .Y(n_647) );
BUFx3_ASAP7_75t_L g911 ( .A(n_289), .Y(n_911) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g493 ( .A(n_293), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_293), .A2(n_332), .B1(n_611), .B2(n_613), .Y(n_666) );
NOR2x1_ASAP7_75t_L g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g596 ( .A(n_295), .Y(n_596) );
AND2x4_ASAP7_75t_L g782 ( .A(n_295), .B(n_775), .Y(n_782) );
BUFx2_ASAP7_75t_L g833 ( .A(n_295), .Y(n_833) );
INVx1_ASAP7_75t_L g954 ( .A(n_296), .Y(n_954) );
OAI211xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_302), .C(n_307), .Y(n_297) );
BUFx4f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x6_ASAP7_75t_L g604 ( .A(n_300), .B(n_605), .Y(n_604) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_300), .Y(n_682) );
INVx4_ASAP7_75t_L g891 ( .A(n_300), .Y(n_891) );
BUFx4f_ASAP7_75t_L g1090 ( .A(n_300), .Y(n_1090) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx3_ASAP7_75t_L g498 ( .A(n_301), .Y(n_498) );
INVx2_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_305), .Y(n_501) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g1047 ( .A(n_309), .Y(n_1047) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g326 ( .A(n_310), .Y(n_326) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_310), .Y(n_662) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g483 ( .A(n_311), .Y(n_483) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g663 ( .A(n_313), .Y(n_663) );
INVx2_ASAP7_75t_L g831 ( .A(n_313), .Y(n_831) );
INVx1_ASAP7_75t_L g919 ( .A(n_313), .Y(n_919) );
OAI221xp5_ASAP7_75t_L g1089 ( .A1(n_313), .A2(n_1090), .B1(n_1091), .B2(n_1092), .C(n_1095), .Y(n_1089) );
OAI221xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B1(n_318), .B2(n_323), .C(n_324), .Y(n_314) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_316), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
OAI22x1_ASAP7_75t_SL g582 ( .A1(n_316), .A2(n_546), .B1(n_577), .B2(n_583), .Y(n_582) );
INVx2_ASAP7_75t_SL g687 ( .A(n_316), .Y(n_687) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g577 ( .A(n_320), .Y(n_577) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_320), .Y(n_656) );
INVx4_ASAP7_75t_L g691 ( .A(n_320), .Y(n_691) );
INVx2_ASAP7_75t_L g1043 ( .A(n_320), .Y(n_1043) );
INVx8_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g774 ( .A(n_321), .B(n_775), .Y(n_774) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
HB1xp67_ASAP7_75t_SL g1032 ( .A(n_328), .Y(n_1032) );
INVx4_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g584 ( .A(n_329), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_329), .B(n_585), .Y(n_697) );
INVx4_ASAP7_75t_L g824 ( .A(n_329), .Y(n_824) );
NAND4xp25_ASAP7_75t_L g966 ( .A(n_329), .B(n_967), .C(n_968), .D(n_969), .Y(n_966) );
INVx1_ASAP7_75t_SL g1081 ( .A(n_329), .Y(n_1081) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g491 ( .A(n_332), .Y(n_491) );
INVx1_ASAP7_75t_L g1088 ( .A(n_332), .Y(n_1088) );
INVx4_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx3_ASAP7_75t_L g827 ( .A(n_334), .Y(n_827) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g668 ( .A(n_337), .Y(n_668) );
HB1xp67_ASAP7_75t_L g975 ( .A(n_337), .Y(n_975) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g922 ( .A(n_338), .Y(n_922) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND3x4_ASAP7_75t_L g406 ( .A(n_339), .B(n_383), .C(n_407), .Y(n_406) );
OAI31xp33_ASAP7_75t_SL g523 ( .A1(n_339), .A2(n_524), .A3(n_530), .B(n_541), .Y(n_523) );
INVx2_ASAP7_75t_SL g1048 ( .A(n_339), .Y(n_1048) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g507 ( .A(n_340), .Y(n_507) );
AOI21xp33_ASAP7_75t_SL g341 ( .A1(n_342), .A2(n_360), .B(n_361), .Y(n_341) );
AOI211x1_ASAP7_75t_L g445 ( .A1(n_342), .A2(n_446), .B(n_447), .C(n_472), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_342), .A2(n_631), .B(n_632), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_342), .A2(n_794), .B1(n_795), .B2(n_796), .C(n_797), .Y(n_793) );
NAND2xp33_ASAP7_75t_L g870 ( .A(n_342), .B(n_871), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_342), .A2(n_942), .B(n_943), .Y(n_941) );
AOI21xp33_ASAP7_75t_SL g1024 ( .A1(n_342), .A2(n_1025), .B(n_1026), .Y(n_1024) );
AOI211x1_ASAP7_75t_L g1051 ( .A1(n_342), .A2(n_1052), .B(n_1053), .C(n_1069), .Y(n_1051) );
AOI21xp33_ASAP7_75t_L g1316 ( .A1(n_342), .A2(n_1317), .B(n_1318), .Y(n_1316) );
INVx8_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_356), .Y(n_343) );
INVx1_ASAP7_75t_L g980 ( .A(n_344), .Y(n_980) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_350), .Y(n_344) );
BUFx3_ASAP7_75t_L g545 ( .A(n_345), .Y(n_545) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_346), .Y(n_715) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_L g736 ( .A(n_347), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_348), .Y(n_372) );
INVx2_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
AND2x4_ASAP7_75t_L g405 ( .A(n_348), .B(n_399), .Y(n_405) );
OR2x2_ASAP7_75t_L g432 ( .A(n_348), .B(n_378), .Y(n_432) );
INVx1_ASAP7_75t_L g371 ( .A(n_349), .Y(n_371) );
INVx2_ASAP7_75t_L g399 ( .A(n_349), .Y(n_399) );
OR2x2_ASAP7_75t_L g368 ( .A(n_350), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g434 ( .A(n_350), .Y(n_434) );
INVx1_ASAP7_75t_L g437 ( .A(n_350), .Y(n_437) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g586 ( .A(n_351), .Y(n_586) );
OR2x2_ASAP7_75t_L g704 ( .A(n_351), .B(n_563), .Y(n_704) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_351), .Y(n_760) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g527 ( .A(n_354), .Y(n_527) );
INVx1_ASAP7_75t_L g554 ( .A(n_354), .Y(n_554) );
INVx3_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
BUFx3_ASAP7_75t_L g407 ( .A(n_355), .Y(n_407) );
NAND2xp33_ASAP7_75t_SL g563 ( .A(n_355), .B(n_383), .Y(n_563) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AND2x4_ASAP7_75t_L g392 ( .A(n_357), .B(n_380), .Y(n_392) );
INVx1_ASAP7_75t_L g600 ( .A(n_357), .Y(n_600) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g423 ( .A(n_358), .Y(n_423) );
INVx1_ASAP7_75t_L g601 ( .A(n_359), .Y(n_601) );
INVx2_ASAP7_75t_L g474 ( .A(n_362), .Y(n_474) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_368), .Y(n_362) );
INVx2_ASAP7_75t_SL g597 ( .A(n_363), .Y(n_597) );
AND2x4_ASAP7_75t_L g835 ( .A(n_363), .B(n_368), .Y(n_835) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVxp67_ASAP7_75t_L g384 ( .A(n_367), .Y(n_384) );
INVx1_ASAP7_75t_L g516 ( .A(n_367), .Y(n_516) );
INVx1_ASAP7_75t_L g789 ( .A(n_367), .Y(n_789) );
INVx2_ASAP7_75t_L g981 ( .A(n_368), .Y(n_981) );
INVx3_ASAP7_75t_L g560 ( .A(n_369), .Y(n_560) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_369), .Y(n_710) );
BUFx6f_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g539 ( .A(n_370), .Y(n_539) );
BUFx3_ASAP7_75t_L g720 ( .A(n_370), .Y(n_720) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
BUFx2_ASAP7_75t_L g749 ( .A(n_371), .Y(n_749) );
INVx2_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
AND2x4_ASAP7_75t_L g415 ( .A(n_372), .B(n_398), .Y(n_415) );
BUFx2_ASAP7_75t_L g745 ( .A(n_372), .Y(n_745) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_384), .Y(n_373) );
OR2x6_ASAP7_75t_L g454 ( .A(n_374), .B(n_384), .Y(n_454) );
INVx2_ASAP7_75t_L g532 ( .A(n_374), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_375), .B(n_380), .Y(n_374) );
INVx8_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
AND2x2_ASAP7_75t_L g553 ( .A(n_375), .B(n_554), .Y(n_553) );
BUFx3_ASAP7_75t_L g565 ( .A(n_375), .Y(n_565) );
BUFx3_ASAP7_75t_L g626 ( .A(n_375), .Y(n_626) );
HB1xp67_ASAP7_75t_L g994 ( .A(n_375), .Y(n_994) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AND2x4_ASAP7_75t_L g411 ( .A(n_376), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g412 ( .A(n_379), .Y(n_412) );
AND2x6_ASAP7_75t_L g535 ( .A(n_380), .B(n_390), .Y(n_535) );
AND2x2_ASAP7_75t_L g537 ( .A(n_380), .B(n_397), .Y(n_537) );
INVx1_ASAP7_75t_L g540 ( .A(n_380), .Y(n_540) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
NAND3x1_ASAP7_75t_L g422 ( .A(n_381), .B(n_423), .C(n_424), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g551 ( .A(n_381), .B(n_424), .Y(n_551) );
INVx1_ASAP7_75t_L g732 ( .A(n_381), .Y(n_732) );
OR2x6_ASAP7_75t_L g735 ( .A(n_381), .B(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g739 ( .A(n_381), .B(n_405), .Y(n_739) );
OR2x4_ASAP7_75t_L g753 ( .A(n_381), .B(n_432), .Y(n_753) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_383), .Y(n_758) );
NOR3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_428), .C(n_439), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_400), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B1(n_393), .B2(n_394), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_389), .A2(n_394), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_389), .A2(n_394), .B1(n_1349), .B2(n_1350), .Y(n_1348) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
AND2x2_ASAP7_75t_L g612 ( .A(n_390), .B(n_392), .Y(n_612) );
AND2x4_ASAP7_75t_SL g800 ( .A(n_390), .B(n_392), .Y(n_800) );
NAND2x1_ASAP7_75t_L g855 ( .A(n_390), .B(n_392), .Y(n_855) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g394 ( .A(n_392), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g441 ( .A(n_392), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_SL g802 ( .A(n_392), .B(n_395), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_394), .A2(n_611), .B1(n_612), .B2(n_613), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g852 ( .A1(n_394), .A2(n_853), .B1(n_854), .B2(n_856), .Y(n_852) );
AOI221x1_ASAP7_75t_L g982 ( .A1(n_394), .A2(n_854), .B1(n_952), .B2(n_960), .C(n_983), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_394), .A2(n_854), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
AO22x1_ASAP7_75t_L g1055 ( .A1(n_394), .A2(n_612), .B1(n_1056), .B2(n_1057), .Y(n_1055) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI33xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_406), .A3(n_408), .B1(n_416), .B2(n_420), .B3(n_425), .Y(n_400) );
BUFx2_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
INVx8_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_403), .Y(n_548) );
INVx2_ASAP7_75t_L g616 ( .A(n_403), .Y(n_616) );
INVx2_ASAP7_75t_L g805 ( .A(n_403), .Y(n_805) );
INVx3_ASAP7_75t_L g868 ( .A(n_403), .Y(n_868) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g427 ( .A(n_405), .Y(n_427) );
BUFx2_ASAP7_75t_L g442 ( .A(n_405), .Y(n_442) );
BUFx2_ASAP7_75t_L g460 ( .A(n_405), .Y(n_460) );
AND2x2_ASAP7_75t_L g556 ( .A(n_405), .B(n_554), .Y(n_556) );
BUFx3_ASAP7_75t_L g863 ( .A(n_405), .Y(n_863) );
BUFx3_ASAP7_75t_L g461 ( .A(n_406), .Y(n_461) );
INVx1_ASAP7_75t_L g812 ( .A(n_406), .Y(n_812) );
AOI33xp33_ASAP7_75t_L g859 ( .A1(n_406), .A2(n_860), .A3(n_864), .B1(n_866), .B2(n_867), .B3(n_869), .Y(n_859) );
AOI33xp33_ASAP7_75t_L g1013 ( .A1(n_406), .A2(n_420), .A3(n_1014), .B1(n_1015), .B2(n_1018), .B3(n_1019), .Y(n_1013) );
AOI33xp33_ASAP7_75t_L g1341 ( .A1(n_406), .A2(n_722), .A3(n_1342), .B1(n_1343), .B2(n_1345), .B3(n_1346), .Y(n_1341) );
INVx3_ASAP7_75t_L g744 ( .A(n_407), .Y(n_744) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_SL g418 ( .A(n_410), .Y(n_418) );
INVx3_ASAP7_75t_L g543 ( .A(n_410), .Y(n_543) );
INVx5_ASAP7_75t_L g624 ( .A(n_410), .Y(n_624) );
INVx2_ASAP7_75t_SL g986 ( .A(n_410), .Y(n_986) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx8_ASAP7_75t_L g438 ( .A(n_411), .Y(n_438) );
INVx2_ASAP7_75t_L g465 ( .A(n_411), .Y(n_465) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_411), .Y(n_713) );
INVx2_ASAP7_75t_R g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
INVx2_ASAP7_75t_L g1064 ( .A(n_414), .Y(n_1064) );
INVx5_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g419 ( .A(n_415), .Y(n_419) );
AND2x4_ASAP7_75t_L g529 ( .A(n_415), .B(n_527), .Y(n_529) );
BUFx3_ASAP7_75t_L g621 ( .A(n_415), .Y(n_621) );
BUFx12f_ASAP7_75t_L g808 ( .A(n_415), .Y(n_808) );
BUFx2_ASAP7_75t_L g865 ( .A(n_415), .Y(n_865) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI33xp33_ASAP7_75t_L g614 ( .A1(n_420), .A2(n_461), .A3(n_615), .B1(n_618), .B2(n_622), .B3(n_625), .Y(n_614) );
BUFx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g722 ( .A(n_421), .Y(n_722) );
BUFx2_ASAP7_75t_L g869 ( .A(n_421), .Y(n_869) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_421), .Y(n_1067) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g811 ( .A(n_427), .Y(n_811) );
OR2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
OR2x6_ASAP7_75t_L g628 ( .A(n_430), .B(n_433), .Y(n_628) );
INVx2_ASAP7_75t_SL g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx4f_ASAP7_75t_L g707 ( .A(n_432), .Y(n_707) );
OR2x4_ASAP7_75t_L g731 ( .A(n_432), .B(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g838 ( .A(n_434), .B(n_839), .Y(n_838) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_436), .A2(n_913), .B1(n_914), .B2(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_436), .A2(n_945), .B1(n_1071), .B2(n_1072), .Y(n_1070) );
AND2x4_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
AND2x4_ASAP7_75t_L g837 ( .A(n_437), .B(n_616), .Y(n_837) );
AND2x4_ASAP7_75t_L g945 ( .A(n_437), .B(n_616), .Y(n_945) );
INVx3_ASAP7_75t_L g469 ( .A(n_438), .Y(n_469) );
INVx2_ASAP7_75t_SL g927 ( .A(n_438), .Y(n_927) );
INVx3_ASAP7_75t_L g1017 ( .A(n_438), .Y(n_1017) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND4xp25_ASAP7_75t_SL g447 ( .A(n_440), .B(n_448), .C(n_451), .D(n_455), .Y(n_447) );
NAND4xp25_ASAP7_75t_SL g851 ( .A(n_440), .B(n_852), .C(n_857), .D(n_859), .Y(n_851) );
NAND2xp5_ASAP7_75t_SL g1058 ( .A(n_440), .B(n_1059), .Y(n_1058) );
INVx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_441), .Y(n_629) );
INVx3_ASAP7_75t_L g814 ( .A(n_441), .Y(n_814) );
NOR3xp33_ASAP7_75t_L g923 ( .A(n_441), .B(n_924), .C(n_939), .Y(n_923) );
BUFx2_ASAP7_75t_L g617 ( .A(n_442), .Y(n_617) );
XNOR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_453), .B(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_453), .B(n_1000), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_453), .B(n_1060), .Y(n_1059) );
INVx5_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g794 ( .A(n_454), .Y(n_794) );
AOI33xp33_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_461), .A3(n_462), .B1(n_467), .B2(n_470), .B3(n_471), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI33xp33_ASAP7_75t_L g1061 ( .A1(n_461), .A2(n_1062), .A3(n_1063), .B1(n_1065), .B2(n_1067), .B3(n_1068), .Y(n_1061) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
OR2x6_ASAP7_75t_SL g525 ( .A(n_465), .B(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g620 ( .A(n_465), .Y(n_620) );
INVx3_ASAP7_75t_L g839 ( .A(n_465), .Y(n_839) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_470), .Y(n_934) );
INVx2_ASAP7_75t_L g990 ( .A(n_470), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_478), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_476), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_474), .A2(n_876), .B(n_877), .Y(n_875) );
OAI21xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_490), .B(n_504), .Y(n_478) );
AND2x4_ASAP7_75t_L g589 ( .A(n_485), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g896 ( .A(n_486), .Y(n_896) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
OAI211xp5_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_499), .C(n_500), .Y(n_494) );
OAI211xp5_ASAP7_75t_L g916 ( .A1(n_496), .A2(n_917), .B(n_918), .C(n_920), .Y(n_916) );
OAI211xp5_ASAP7_75t_L g971 ( .A1(n_496), .A2(n_972), .B(n_973), .C(n_974), .Y(n_971) );
INVx5_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g569 ( .A(n_498), .B(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g816 ( .A(n_505), .Y(n_816) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g1337 ( .A(n_506), .Y(n_1337) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g579 ( .A(n_507), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g806 ( .A(n_507), .B(n_551), .Y(n_806) );
AOI22xp5_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_510), .B1(n_671), .B2(n_841), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_606), .B1(n_669), .B2(n_670), .Y(n_510) );
INVx1_ASAP7_75t_L g670 ( .A(n_511), .Y(n_670) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AOI211x1_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_517), .B(n_518), .C(n_566), .Y(n_513) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx3_ASAP7_75t_L g998 ( .A(n_515), .Y(n_998) );
AND2x4_ASAP7_75t_L g520 ( .A(n_516), .B(n_521), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_517), .A2(n_553), .B1(n_555), .B2(n_556), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_522), .Y(n_519) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B1(n_536), .B2(n_537), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g587 ( .A1(n_534), .A2(n_555), .B1(n_588), .B2(n_589), .C1(n_591), .C2(n_597), .Y(n_587) );
AOI222xp33_ASAP7_75t_L g567 ( .A1(n_536), .A2(n_568), .B1(n_571), .B2(n_578), .C1(n_581), .C2(n_584), .Y(n_567) );
OR2x6_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_552), .C(n_557), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_545), .B2(n_546), .C(n_547), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g991 ( .A1(n_545), .A2(n_624), .B1(n_972), .B2(n_992), .C(n_993), .Y(n_991) );
INVx3_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
OAI211xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_561), .C(n_564), .Y(n_557) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g1347 ( .A(n_565), .Y(n_1347) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_567), .B(n_587), .C(n_598), .Y(n_566) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g590 ( .A(n_570), .Y(n_590) );
INVx1_ASAP7_75t_L g894 ( .A(n_573), .Y(n_894) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g683 ( .A(n_579), .Y(n_683) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx1_ASAP7_75t_L g605 ( .A(n_593), .Y(n_605) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_602), .B(n_603), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g669 ( .A(n_606), .Y(n_669) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_630), .C(n_633), .Y(n_607) );
NOR3xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_627), .C(n_629), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_614), .Y(n_609) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx8_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_SL g862 ( .A(n_626), .Y(n_862) );
INVx1_ASAP7_75t_L g1021 ( .A(n_626), .Y(n_1021) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_628), .B(n_998), .Y(n_997) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_655), .B(n_667), .Y(n_633) );
BUFx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
HB1xp67_ASAP7_75t_L g1031 ( .A(n_641), .Y(n_1031) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g829 ( .A(n_645), .Y(n_829) );
INVx2_ASAP7_75t_SL g921 ( .A(n_645), .Y(n_921) );
INVx2_ASAP7_75t_L g1083 ( .A(n_645), .Y(n_1083) );
INVx2_ASAP7_75t_L g1329 ( .A(n_645), .Y(n_1329) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g1085 ( .A(n_647), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_648) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx5_ASAP7_75t_L g1099 ( .A(n_656), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_664), .Y(n_657) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1078 ( .A(n_660), .Y(n_1078) );
BUFx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g841 ( .A(n_671), .Y(n_841) );
AO22x1_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_790), .B1(n_791), .B2(n_840), .Y(n_671) );
INVx1_ASAP7_75t_L g840 ( .A(n_672), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_727), .C(n_761), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_701), .Y(n_674) );
OAI33xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_683), .A3(n_684), .B1(n_692), .B2(n_695), .B3(n_698), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_680), .B2(n_681), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_677), .A2(n_693), .B1(n_712), .B2(n_714), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_678), .A2(n_689), .B1(n_699), .B2(n_700), .Y(n_698) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx2_ASAP7_75t_L g1094 ( .A(n_679), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_680), .A2(n_694), .B1(n_717), .B2(n_719), .Y(n_716) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g692 ( .A1(n_682), .A2(n_686), .B1(n_693), .B2(n_694), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_686), .B1(n_688), .B2(n_689), .Y(n_684) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_685), .A2(n_699), .B1(n_706), .B2(n_708), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g1331 ( .A1(n_686), .A2(n_1332), .B1(n_1333), .B2(n_1334), .C(n_1335), .Y(n_1331) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_688), .A2(n_700), .B1(n_724), .B2(n_726), .Y(n_723) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI33xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_705), .A3(n_711), .B1(n_716), .B2(n_721), .B3(n_723), .Y(n_701) );
BUFx3_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
BUFx4f_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx8_ASAP7_75t_L g925 ( .A(n_704), .Y(n_925) );
BUFx2_ASAP7_75t_L g984 ( .A(n_704), .Y(n_984) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g725 ( .A(n_707), .Y(n_725) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g1344 ( .A(n_712), .Y(n_1344) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_713), .Y(n_718) );
AND2x4_ASAP7_75t_L g755 ( .A(n_713), .B(n_732), .Y(n_755) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_713), .Y(n_809) );
INVx3_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g726 ( .A(n_715), .Y(n_726) );
CKINVDCx8_ASAP7_75t_R g936 ( .A(n_715), .Y(n_936) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g985 ( .A1(n_726), .A2(n_986), .B1(n_987), .B2(n_988), .C(n_989), .Y(n_985) );
OAI31xp33_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_737), .A3(n_750), .B(n_756), .Y(n_727) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g932 ( .A(n_736), .Y(n_932) );
CKINVDCx8_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_746), .B2(n_747), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_741), .A2(n_781), .B1(n_783), .B2(n_784), .Y(n_780) );
BUFx3_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
AND2x4_ASAP7_75t_L g748 ( .A(n_744), .B(n_749), .Y(n_748) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_SL g756 ( .A(n_757), .B(n_759), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI31xp33_ASAP7_75t_SL g761 ( .A1(n_762), .A2(n_767), .A3(n_776), .B(n_787), .Y(n_761) );
INVx3_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx3_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx3_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
BUFx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_815), .Y(n_792) );
NAND3xp33_ASAP7_75t_SL g797 ( .A(n_798), .B(n_803), .C(n_814), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B1(n_801), .B2(n_802), .Y(n_798) );
AOI222xp33_ASAP7_75t_L g826 ( .A1(n_799), .A2(n_801), .B1(n_827), .B2(n_828), .C1(n_830), .C2(n_832), .Y(n_826) );
INVx1_ASAP7_75t_L g940 ( .A(n_802), .Y(n_940) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B1(n_810), .B2(n_813), .Y(n_803) );
BUFx2_ASAP7_75t_L g1066 ( .A(n_808), .Y(n_1066) );
AND5x1_ASAP7_75t_L g948 ( .A(n_814), .B(n_949), .C(n_982), .D(n_995), .E(n_999), .Y(n_948) );
INVx2_ASAP7_75t_SL g1023 ( .A(n_814), .Y(n_1023) );
AND4x1_ASAP7_75t_L g1338 ( .A(n_814), .B(n_1339), .C(n_1341), .D(n_1348), .Y(n_1338) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B(n_834), .Y(n_815) );
OAI21xp5_ASAP7_75t_L g878 ( .A1(n_816), .A2(n_879), .B(n_887), .Y(n_878) );
OAI21xp5_ASAP7_75t_L g1073 ( .A1(n_816), .A2(n_1074), .B(n_1087), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g817 ( .A(n_818), .B(n_821), .C(n_826), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_819), .A2(n_820), .B1(n_837), .B2(n_838), .Y(n_836) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_827), .B(n_952), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_833), .A2(n_960), .B1(n_961), .B2(n_962), .Y(n_959) );
INVx2_ASAP7_75t_SL g977 ( .A(n_838), .Y(n_977) );
INVx1_ASAP7_75t_L g1103 ( .A(n_842), .Y(n_1103) );
XNOR2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_1004), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_900), .B1(n_1002), .B2(n_1003), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_SL g1002 ( .A(n_846), .Y(n_1002) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NAND2x1p5_ASAP7_75t_L g847 ( .A(n_848), .B(n_872), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_870), .Y(n_849) );
INVxp67_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
NOR2xp33_ASAP7_75t_SL g897 ( .A(n_851), .B(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_870), .B(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_878), .Y(n_874) );
OAI211xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B(n_892), .C(n_895), .Y(n_888) );
INVx2_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx2_ASAP7_75t_L g958 ( .A(n_891), .Y(n_958) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1003 ( .A(n_900), .Y(n_1003) );
OA22x2_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_946), .B1(n_947), .B2(n_1001), .Y(n_900) );
INVx1_ASAP7_75t_L g1001 ( .A(n_901), .Y(n_1001) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
AND4x1_ASAP7_75t_L g903 ( .A(n_904), .B(n_923), .C(n_941), .D(n_944), .Y(n_903) );
OAI21xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_915), .B(n_922), .Y(n_904) );
INVx2_ASAP7_75t_SL g908 ( .A(n_909), .Y(n_908) );
OAI221xp5_ASAP7_75t_L g935 ( .A1(n_917), .A2(n_927), .B1(n_936), .B2(n_937), .C(n_938), .Y(n_935) );
OAI22xp5_ASAP7_75t_SL g924 ( .A1(n_925), .A2(n_926), .B1(n_934), .B2(n_935), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_927), .A2(n_928), .B1(n_929), .B2(n_930), .C(n_933), .Y(n_926) );
INVx3_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
BUFx2_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
INVx2_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
AOI21xp5_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_975), .B(n_976), .Y(n_949) );
NAND4xp25_ASAP7_75t_L g950 ( .A(n_951), .B(n_953), .C(n_966), .D(n_971), .Y(n_950) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B1(n_964), .B2(n_965), .Y(n_953) );
INVx4_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
BUFx6f_ASAP7_75t_L g1040 ( .A(n_957), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g978 ( .A1(n_961), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
OAI22xp5_ASAP7_75t_SL g983 ( .A1(n_984), .A2(n_985), .B1(n_990), .B2(n_991), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1006), .B1(n_1049), .B2(n_1101), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1024), .C(n_1027), .Y(n_1007) );
NOR3xp33_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1022), .C(n_1023), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1013), .Y(n_1009) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
OAI21xp5_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1037), .B(n_1048), .Y(n_1027) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1041), .B1(n_1042), .B2(n_1044), .C(n_1045), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_1039), .A2(n_1097), .B1(n_1098), .B2(n_1099), .Y(n_1096) );
INVx2_ASAP7_75t_L g1039 ( .A(n_1040), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1333 ( .A(n_1042), .Y(n_1333) );
BUFx6f_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1049), .Y(n_1101) );
XOR2x2_ASAP7_75t_L g1049 ( .A(n_1050), .B(n_1100), .Y(n_1049) );
NAND2xp5_ASAP7_75t_SL g1050 ( .A(n_1051), .B(n_1073), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1061), .Y(n_1053) );
NOR2xp33_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1058), .Y(n_1054) );
NAND3xp33_ASAP7_75t_SL g1074 ( .A(n_1075), .B(n_1076), .C(n_1086), .Y(n_1074) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_SL g1084 ( .A(n_1085), .Y(n_1084) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx4_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
OAI221xp5_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1308), .B1(n_1311), .B2(n_1352), .C(n_1358), .Y(n_1104) );
NOR2xp67_ASAP7_75t_SL g1105 ( .A(n_1106), .B(n_1246), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1207), .Y(n_1106) );
A2O1A1Ixp33_ASAP7_75t_SL g1107 ( .A1(n_1108), .A2(n_1123), .B(n_1156), .C(n_1202), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1108), .B(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1108), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1244 ( .A(n_1108), .B(n_1245), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1108), .B(n_1194), .Y(n_1269) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1108), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1108), .B(n_1140), .Y(n_1305) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1109), .Y(n_1159) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1109), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1109), .B(n_1154), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1109), .B(n_1201), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1109), .B(n_1140), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1117), .Y(n_1109) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1111), .Y(n_1310) );
AND2x6_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1113), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1115 ( .A(n_1112), .B(n_1116), .Y(n_1115) );
AND2x4_ASAP7_75t_L g1118 ( .A(n_1112), .B(n_1119), .Y(n_1118) );
AND2x6_ASAP7_75t_L g1121 ( .A(n_1112), .B(n_1122), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1112), .B(n_1116), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1112), .B(n_1116), .Y(n_1205) );
OAI21xp5_ASAP7_75t_L g1365 ( .A1(n_1113), .A2(n_1366), .B(n_1367), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1114), .B(n_1120), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1139), .B1(n_1146), .B2(n_1155), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NOR2xp33_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1136), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1126), .B(n_1143), .Y(n_1256) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1127), .B(n_1165), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1220 ( .A(n_1127), .B(n_1171), .Y(n_1220) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1128), .B(n_1133), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1128), .B(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1128), .B(n_1188), .Y(n_1187) );
A2O1A1Ixp33_ASAP7_75t_L g1249 ( .A1(n_1128), .A2(n_1231), .B(n_1250), .C(n_1252), .Y(n_1249) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1129), .B(n_1138), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1129), .B(n_1133), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1129), .B(n_1165), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1129), .B(n_1281), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_1130), .B(n_1131), .Y(n_1129) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1133), .Y(n_1138) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1133), .Y(n_1155) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1133), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1133), .B(n_1171), .Y(n_1240) );
NAND2x1_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1135), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1136), .B(n_1171), .Y(n_1272) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1137), .B(n_1171), .Y(n_1170) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1143), .Y(n_1139) );
CKINVDCx5p33_ASAP7_75t_R g1154 ( .A(n_1140), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1174 ( .A(n_1140), .B(n_1151), .Y(n_1174) );
NAND2xp5_ASAP7_75t_L g1190 ( .A(n_1140), .B(n_1191), .Y(n_1190) );
OAI22xp5_ASAP7_75t_L g1270 ( .A1(n_1140), .A2(n_1234), .B1(n_1253), .B2(n_1271), .Y(n_1270) );
AND2x4_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
INVx3_ASAP7_75t_L g1148 ( .A(n_1143), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g1163 ( .A(n_1143), .Y(n_1163) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_1143), .B(n_1165), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1213 ( .A(n_1143), .B(n_1187), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1143), .B(n_1217), .Y(n_1241) );
AND2x4_ASAP7_75t_SL g1143 ( .A(n_1144), .B(n_1145), .Y(n_1143) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
NOR2xp33_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1149), .Y(n_1147) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1148), .B(n_1171), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1148), .B(n_1150), .Y(n_1201) );
NOR2xp33_ASAP7_75t_L g1259 ( .A(n_1148), .B(n_1260), .Y(n_1259) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_1148), .B(n_1180), .Y(n_1267) );
CKINVDCx14_ASAP7_75t_R g1286 ( .A(n_1148), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1148), .B(n_1169), .Y(n_1289) );
AOI211xp5_ASAP7_75t_L g1215 ( .A1(n_1149), .A2(n_1216), .B(n_1218), .C(n_1221), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1154), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1150), .B(n_1211), .Y(n_1210) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1150), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1150), .B(n_1212), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1284 ( .A(n_1150), .B(n_1285), .Y(n_1284) );
INVx2_ASAP7_75t_SL g1150 ( .A(n_1151), .Y(n_1150) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1151), .B(n_1154), .Y(n_1184) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1151), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1154), .B(n_1159), .Y(n_1158) );
NAND3xp33_ASAP7_75t_L g1258 ( .A(n_1154), .B(n_1180), .C(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1155), .B(n_1171), .Y(n_1263) );
NAND4xp25_ASAP7_75t_SL g1156 ( .A(n_1157), .B(n_1175), .C(n_1192), .D(n_1198), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1160), .B1(n_1169), .B2(n_1172), .Y(n_1157) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1159), .Y(n_1214) );
OAI211xp5_ASAP7_75t_L g1278 ( .A1(n_1159), .A2(n_1279), .B(n_1282), .C(n_1284), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1168), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
OAI21xp5_ASAP7_75t_L g1226 ( .A1(n_1162), .A2(n_1173), .B(n_1227), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1164), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1163), .B(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1219 ( .A(n_1163), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1163), .B(n_1233), .Y(n_1235) );
OR2x2_ASAP7_75t_L g1251 ( .A(n_1163), .B(n_1190), .Y(n_1251) );
NOR2xp33_ASAP7_75t_L g1252 ( .A(n_1163), .B(n_1253), .Y(n_1252) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1165), .Y(n_1171) );
OR2x2_ASAP7_75t_L g1212 ( .A(n_1165), .B(n_1213), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1165), .B(n_1188), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1273 ( .A1(n_1165), .A2(n_1274), .B1(n_1276), .B2(n_1277), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1167), .Y(n_1165) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1168), .Y(n_1176) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1199 ( .A(n_1170), .B(n_1200), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1178 ( .A(n_1171), .B(n_1179), .Y(n_1178) );
NAND2xp5_ASAP7_75t_L g1243 ( .A(n_1171), .B(n_1187), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_1171), .B(n_1267), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_1173), .B(n_1230), .Y(n_1229) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
O2A1O1Ixp33_ASAP7_75t_L g1175 ( .A1(n_1176), .A2(n_1177), .B(n_1181), .C(n_1185), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1279 ( .A1(n_1176), .A2(n_1184), .B1(n_1260), .B2(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1178), .Y(n_1177) );
AOI21xp5_ASAP7_75t_L g1185 ( .A1(n_1178), .A2(n_1186), .B(n_1190), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1196 ( .A(n_1179), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1180), .B(n_1189), .Y(n_1211) );
OAI211xp5_ASAP7_75t_L g1238 ( .A1(n_1180), .A2(n_1183), .B(n_1239), .C(n_1241), .Y(n_1238) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1183), .Y(n_1253) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
OR2x2_ASAP7_75t_L g1299 ( .A(n_1184), .B(n_1300), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1189), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1187), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1189), .Y(n_1281) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1190), .Y(n_1225) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1190), .Y(n_1245) );
INVx2_ASAP7_75t_L g1194 ( .A(n_1191), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1195), .Y(n_1192) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1194), .B(n_1217), .Y(n_1216) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_1194), .A2(n_1291), .B(n_1293), .Y(n_1290) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
A2O1A1Ixp33_ASAP7_75t_L g1222 ( .A1(n_1196), .A2(n_1223), .B(n_1224), .C(n_1226), .Y(n_1222) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1197), .Y(n_1292) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
CKINVDCx14_ASAP7_75t_R g1221 ( .A(n_1202), .Y(n_1221) );
A2O1A1Ixp33_ASAP7_75t_L g1287 ( .A1(n_1202), .A2(n_1288), .B(n_1290), .C(n_1295), .Y(n_1287) );
INVx3_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
OAI221xp5_ASAP7_75t_L g1261 ( .A1(n_1203), .A2(n_1232), .B1(n_1236), .B2(n_1262), .C(n_1264), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1206), .Y(n_1203) );
NOR5xp2_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1215), .C(n_1222), .D(n_1228), .E(n_1242), .Y(n_1207) );
AOI21xp33_ASAP7_75t_L g1208 ( .A1(n_1209), .A2(n_1212), .B(n_1214), .Y(n_1208) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1210), .Y(n_1209) );
INVxp67_ASAP7_75t_L g1223 ( .A(n_1211), .Y(n_1223) );
OR2x2_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1220), .Y(n_1218) );
INVx2_ASAP7_75t_L g1227 ( .A(n_1220), .Y(n_1227) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
AOI211xp5_ASAP7_75t_L g1254 ( .A1(n_1225), .A2(n_1255), .B(n_1257), .C(n_1261), .Y(n_1254) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1227), .B(n_1286), .Y(n_1294) );
OAI221xp5_ASAP7_75t_SL g1228 ( .A1(n_1229), .A2(n_1232), .B1(n_1234), .B2(n_1236), .C(n_1238), .Y(n_1228) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1229), .Y(n_1277) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
NOR2xp33_ASAP7_75t_L g1242 ( .A(n_1243), .B(n_1244), .Y(n_1242) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1243), .Y(n_1268) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1244), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1297), .Y(n_1246) );
OAI21xp5_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1278), .B(n_1287), .Y(n_1247) );
NAND4xp25_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1254), .C(n_1265), .D(n_1273), .Y(n_1248) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
OAI21xp5_ASAP7_75t_SL g1298 ( .A1(n_1262), .A2(n_1299), .B(n_1301), .Y(n_1298) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
O2A1O1Ixp33_ASAP7_75t_L g1265 ( .A1(n_1266), .A2(n_1268), .B(n_1269), .C(n_1270), .Y(n_1265) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_1266), .A2(n_1286), .B1(n_1298), .B2(n_1306), .Y(n_1297) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx2_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1272), .B(n_1286), .Y(n_1285) );
OAI31xp33_ASAP7_75t_L g1301 ( .A1(n_1274), .A2(n_1302), .A3(n_1304), .B(n_1305), .Y(n_1301) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
A2O1A1Ixp33_ASAP7_75t_L g1306 ( .A1(n_1275), .A2(n_1299), .B(n_1303), .C(n_1307), .Y(n_1306) );
INVxp67_ASAP7_75t_SL g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1299), .Y(n_1304) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1305), .Y(n_1307) );
CKINVDCx20_ASAP7_75t_R g1308 ( .A(n_1309), .Y(n_1308) );
CKINVDCx20_ASAP7_75t_R g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
AO21x2_ASAP7_75t_L g1313 ( .A1(n_1314), .A2(n_1315), .B(n_1351), .Y(n_1313) );
INVxp33_ASAP7_75t_L g1364 ( .A(n_1315), .Y(n_1364) );
NAND3xp33_ASAP7_75t_SL g1315 ( .A(n_1316), .B(n_1319), .C(n_1338), .Y(n_1315) );
OAI21xp5_ASAP7_75t_L g1319 ( .A1(n_1320), .A2(n_1330), .B(n_1337), .Y(n_1319) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1327), .Y(n_1336) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
CKINVDCx20_ASAP7_75t_R g1352 ( .A(n_1353), .Y(n_1352) );
CKINVDCx20_ASAP7_75t_R g1353 ( .A(n_1354), .Y(n_1353) );
INVx3_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
BUFx3_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
HB1xp67_ASAP7_75t_SL g1359 ( .A(n_1360), .Y(n_1359) );
INVxp33_ASAP7_75t_L g1361 ( .A(n_1362), .Y(n_1361) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
endmodule