module fake_jpeg_14212_n_406 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_406);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_406;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_292;
wire n_213;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_7),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_44),
.B(n_56),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_45),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_14),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_54),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_57),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

AND2x6_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_1),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_59),
.B(n_22),
.C(n_31),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_27),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_65),
.B(n_69),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_2),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_83),
.Y(n_138)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_17),
.B(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_84),
.B(n_85),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_87),
.Y(n_139)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_41),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_29),
.B1(n_24),
.B2(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_90),
.A2(n_115),
.B1(n_128),
.B2(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_93),
.B(n_116),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_122),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_32),
.B1(n_39),
.B2(n_41),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_123),
.B(n_61),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_29),
.B1(n_24),
.B2(n_39),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_53),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_46),
.A2(n_41),
.B1(n_24),
.B2(n_35),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_40),
.B1(n_82),
.B2(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_81),
.B(n_35),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_119),
.B(n_125),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_76),
.A2(n_32),
.B1(n_42),
.B2(n_28),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_31),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_37),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_126),
.B(n_129),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_52),
.A2(n_34),
.B1(n_40),
.B2(n_32),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_37),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_57),
.A2(n_40),
.B1(n_26),
.B2(n_42),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_131),
.A2(n_58),
.B1(n_45),
.B2(n_63),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_66),
.A2(n_40),
.B1(n_42),
.B2(n_33),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_143),
.A2(n_159),
.B1(n_113),
.B2(n_137),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_92),
.B(n_36),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_144),
.B(n_153),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_145),
.A2(n_173),
.B(n_181),
.Y(n_192)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_146),
.Y(n_228)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_111),
.Y(n_149)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_151),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_2),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_155),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_2),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_107),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_118),
.A2(n_77),
.B1(n_70),
.B2(n_67),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_3),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_174),
.Y(n_201)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_163),
.Y(n_209)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_79),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_164),
.B(n_169),
.Y(n_224)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_68),
.B1(n_64),
.B2(n_60),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_167),
.B1(n_180),
.B2(n_188),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

OR2x2_ASAP7_75t_SL g169 ( 
.A(n_104),
.B(n_45),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_63),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_172),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_3),
.B(n_4),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_171),
.A2(n_164),
.B(n_170),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_139),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_62),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_118),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_99),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_175),
.A2(n_136),
.B1(n_114),
.B2(n_108),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_124),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx13_ASAP7_75t_L g177 ( 
.A(n_95),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_177),
.Y(n_210)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_99),
.Y(n_178)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_10),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_106),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_102),
.B(n_11),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_11),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_189),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_12),
.Y(n_184)
);

OA21x2_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_101),
.B(n_112),
.Y(n_215)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_186),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_137),
.B1(n_98),
.B2(n_96),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_123),
.A2(n_12),
.B1(n_13),
.B2(n_110),
.Y(n_188)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_103),
.B(n_12),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_154),
.A2(n_150),
.A3(n_169),
.B1(n_185),
.B2(n_152),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_L g261 ( 
.A1(n_190),
.A2(n_218),
.B(n_156),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_108),
.B1(n_94),
.B2(n_113),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_196),
.A2(n_197),
.B1(n_149),
.B2(n_162),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_147),
.A2(n_110),
.B1(n_136),
.B2(n_94),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_204),
.A2(n_206),
.B1(n_212),
.B2(n_149),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_143),
.A2(n_112),
.B1(n_103),
.B2(n_101),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_217),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_150),
.A2(n_95),
.A3(n_96),
.B1(n_141),
.B2(n_98),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_189),
.B(n_171),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_150),
.B(n_141),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_225),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_146),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_155),
.B(n_13),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_179),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_181),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_204),
.A2(n_172),
.B1(n_170),
.B2(n_145),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_229),
.A2(n_249),
.B1(n_251),
.B2(n_260),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_231),
.A2(n_236),
.B1(n_207),
.B2(n_208),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_232),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_262),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_234),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_243),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_182),
.B1(n_175),
.B2(n_151),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_199),
.C(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_242),
.C(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_203),
.Y(n_240)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_240),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_148),
.C(n_168),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_199),
.B(n_160),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_205),
.B(n_161),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_252),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_220),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_257),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_224),
.A2(n_219),
.B(n_192),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_248),
.A2(n_250),
.B(n_255),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_184),
.B1(n_181),
.B2(n_173),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_192),
.A2(n_184),
.B(n_173),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_157),
.B1(n_158),
.B2(n_178),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_186),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_165),
.C(n_177),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_163),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_187),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_207),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_195),
.B(n_187),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_215),
.A2(n_183),
.B1(n_187),
.B2(n_156),
.Y(n_260)
);

OR2x6_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_210),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_226),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_261),
.A2(n_223),
.B(n_191),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_267),
.B(n_241),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_216),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_268),
.B(n_286),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_247),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_232),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_273),
.B(n_281),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_223),
.B(n_194),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_275),
.A2(n_284),
.B(n_255),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_236),
.A2(n_197),
.B1(n_200),
.B2(n_208),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_194),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_230),
.A2(n_200),
.B1(n_198),
.B2(n_193),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_231),
.A2(n_198),
.B1(n_193),
.B2(n_202),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_235),
.B(n_216),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_251),
.B(n_202),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_289),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_243),
.B(n_202),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_290),
.B(n_245),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_305),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_248),
.B1(n_234),
.B2(n_250),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_312),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_229),
.B1(n_262),
.B2(n_241),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_256),
.Y(n_298)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_265),
.B(n_246),
.CI(n_239),
.CON(n_299),
.SN(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_299),
.A2(n_317),
.B(n_274),
.C(n_279),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_242),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_304),
.C(n_310),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_301),
.B(n_280),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_244),
.B1(n_240),
.B2(n_238),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_270),
.B(n_239),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_275),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_269),
.Y(n_306)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_306),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_309),
.A2(n_276),
.B(n_284),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_267),
.B(n_254),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_277),
.A2(n_253),
.B1(n_255),
.B2(n_257),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_271),
.Y(n_313)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

OAI32xp33_ASAP7_75t_L g314 ( 
.A1(n_271),
.A2(n_252),
.A3(n_249),
.B1(n_237),
.B2(n_259),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_214),
.C(n_260),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

AOI22x1_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_277),
.B1(n_289),
.B2(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_273),
.B(n_214),
.Y(n_317)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_319),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_312),
.A2(n_284),
.B1(n_272),
.B2(n_282),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_292),
.A2(n_284),
.B1(n_276),
.B2(n_281),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_296),
.A2(n_284),
.B1(n_265),
.B2(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_294),
.A2(n_284),
.B1(n_311),
.B2(n_295),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_328),
.B(n_310),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_294),
.A2(n_287),
.B(n_289),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_330),
.B(n_309),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_293),
.A2(n_285),
.B1(n_291),
.B2(n_274),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_332),
.A2(n_339),
.B1(n_322),
.B2(n_337),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_335),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_293),
.A2(n_279),
.B1(n_291),
.B2(n_288),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_334),
.B(n_300),
.C(n_304),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_352),
.C(n_353),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_297),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_341),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_342),
.B(n_343),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_301),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_324),
.A2(n_305),
.B1(n_303),
.B2(n_316),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_344),
.B(n_350),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_351),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_324),
.A2(n_314),
.B1(n_299),
.B2(n_288),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_348),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_299),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_320),
.B(n_213),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_213),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_209),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_326),
.B(n_209),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_355),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_156),
.C(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);

AO221x1_ASAP7_75t_L g358 ( 
.A1(n_345),
.A2(n_329),
.B1(n_330),
.B2(n_335),
.C(n_321),
.Y(n_358)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

O2A1O1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_345),
.A2(n_347),
.B(n_318),
.C(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_349),
.B(n_339),
.Y(n_362)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_366),
.Y(n_381)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_356),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_355),
.A2(n_327),
.B1(n_318),
.B2(n_332),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_368),
.A2(n_352),
.B1(n_319),
.B2(n_353),
.Y(n_375)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_371),
.B(n_348),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_369),
.B(n_340),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_374),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_343),
.C(n_342),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_377),
.C(n_363),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_376),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_319),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_331),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_367),
.B(n_370),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_380),
.A2(n_365),
.B(n_359),
.Y(n_388)
);

AOI211xp5_ASAP7_75t_L g382 ( 
.A1(n_378),
.A2(n_367),
.B(n_366),
.C(n_358),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_382),
.B(n_371),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_383),
.B(n_376),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_363),
.C(n_359),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_385),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_379),
.A2(n_362),
.B(n_361),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_365),
.Y(n_392)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_375),
.A2(n_361),
.B(n_360),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_389),
.B(n_377),
.Y(n_391)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_391),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_392),
.B(n_395),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_393),
.B(n_394),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_387),
.B(n_384),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_381),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_398),
.Y(n_401)
);

NAND3xp33_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_396),
.C(n_399),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_402),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_403),
.A2(n_400),
.B1(n_381),
.B2(n_391),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_404),
.A2(n_386),
.B1(n_389),
.B2(n_401),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_405),
.B(n_386),
.Y(n_406)
);


endmodule