module fake_ariane_2337_n_21 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_21);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_21;

wire n_13;
wire n_20;
wire n_17;
wire n_18;
wire n_11;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_10;

AOI22xp5_ASAP7_75t_L g10 ( 
.A1(n_4),
.A2(n_0),
.B1(n_3),
.B2(n_9),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_7),
.B(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2x1_ASAP7_75t_SL g17 ( 
.A(n_16),
.B(n_11),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_13),
.C(n_10),
.Y(n_18)
);

NOR5xp2_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_16),
.C(n_15),
.D(n_11),
.E(n_5),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_0),
.Y(n_20)
);

OAI222xp33_ASAP7_75t_L g21 ( 
.A1(n_20),
.A2(n_12),
.B1(n_19),
.B2(n_5),
.C1(n_1),
.C2(n_2),
.Y(n_21)
);


endmodule