module fake_jpeg_28805_n_121 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_121);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_1),
.Y(n_60)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_15),
.B1(n_17),
.B2(n_22),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_50),
.B1(n_57),
.B2(n_49),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_43),
.A2(n_46),
.B1(n_53),
.B2(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_16),
.B1(n_33),
.B2(n_35),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_11),
.B1(n_23),
.B2(n_21),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_54),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_28),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_29),
.B(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_36),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_56)
);

NOR3xp33_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_24),
.C(n_3),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_3),
.B(n_5),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_62),
.B(n_73),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_37),
.B(n_27),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_65),
.B(n_70),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_34),
.B(n_5),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_40),
.B1(n_41),
.B2(n_24),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_74),
.B1(n_45),
.B2(n_47),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_69),
.Y(n_86)
);

FAx1_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_50),
.CI(n_42),
.CON(n_69),
.SN(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_58),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_61),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_59),
.B(n_61),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_65),
.B(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_47),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_83),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_85),
.B(n_89),
.Y(n_92)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_76),
.B1(n_69),
.B2(n_71),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_86),
.B(n_79),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_96),
.B(n_97),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_80),
.B(n_63),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_82),
.B1(n_85),
.B2(n_84),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_101),
.A2(n_106),
.B1(n_86),
.B2(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_63),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_79),
.C(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_112),
.B(n_105),
.C(n_100),
.Y(n_114)
);

NAND5xp2_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_96),
.C(n_100),
.D(n_90),
.E(n_85),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_106),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_115),
.Y(n_117)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_111),
.B(n_98),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g119 ( 
.A1(n_118),
.A2(n_116),
.A3(n_102),
.B1(n_117),
.B2(n_112),
.C1(n_110),
.C2(n_99),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_76),
.B(n_69),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_75),
.Y(n_121)
);


endmodule