module fake_jpeg_15825_n_173 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_11),
.B(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_35),
.A2(n_36),
.B1(n_40),
.B2(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_20),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_37),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_47),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_7),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_23),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_28),
.B(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_SL g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_SL g60 ( 
.A(n_56),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_32),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_57),
.A2(n_18),
.B1(n_16),
.B2(n_13),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_12),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_62),
.A2(n_64),
.B1(n_39),
.B2(n_41),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_43),
.A2(n_30),
.B1(n_27),
.B2(n_26),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_15),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_72),
.B(n_22),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_49),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_55),
.A2(n_30),
.B1(n_31),
.B2(n_21),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_71),
.B(n_79),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_47),
.B(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_35),
.B1(n_14),
.B2(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_48),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_36),
.B(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_40),
.A2(n_34),
.B1(n_25),
.B2(n_14),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_75),
.B1(n_76),
.B2(n_86),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_14),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_106),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_107),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_25),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_102),
.B(n_105),
.Y(n_131)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_22),
.B(n_38),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_104),
.A2(n_110),
.B(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_39),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_41),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_72),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_86),
.B1(n_73),
.B2(n_64),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_74),
.B1(n_63),
.B2(n_67),
.Y(n_116)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_61),
.B1(n_68),
.B2(n_93),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_113),
.B1(n_104),
.B2(n_105),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_93),
.A2(n_62),
.B(n_68),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_106),
.B(n_95),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_120),
.C(n_126),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_87),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_66),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_125),
.B(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_80),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_96),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_80),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_63),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_92),
.B(n_67),
.Y(n_133)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_112),
.B1(n_107),
.B2(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_142),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_143),
.A2(n_135),
.B1(n_132),
.B2(n_117),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_100),
.Y(n_145)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_145),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_147),
.B1(n_124),
.B2(n_128),
.Y(n_158)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_148),
.A2(n_129),
.B1(n_103),
.B2(n_61),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_151),
.A2(n_122),
.B1(n_139),
.B2(n_133),
.C(n_141),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_125),
.B1(n_128),
.B2(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_140),
.A2(n_143),
.B1(n_136),
.B2(n_138),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_140),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_130),
.C(n_121),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_164),
.B1(n_153),
.B2(n_151),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_118),
.B1(n_138),
.B2(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_157),
.B1(n_153),
.B2(n_156),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_166),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_161),
.A2(n_150),
.B1(n_154),
.B2(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_167),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_168),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_L g172 ( 
.A1(n_170),
.A2(n_98),
.A3(n_123),
.B1(n_129),
.B2(n_155),
.C(n_171),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_167),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_98),
.Y(n_173)
);


endmodule