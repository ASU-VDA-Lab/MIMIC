module fake_jpeg_27659_n_176 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx2_ASAP7_75t_SL g61 ( 
.A(n_34),
.Y(n_61)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_3),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_26),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_26),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_20),
.B1(n_30),
.B2(n_16),
.Y(n_53)
);

OAI211xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_59),
.B(n_16),
.C(n_24),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_20),
.B1(n_30),
.B2(n_24),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_57),
.B1(n_37),
.B2(n_40),
.Y(n_71)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_42),
.A2(n_32),
.B1(n_21),
.B2(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_78),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_28),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_61),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_63),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_41),
.B1(n_43),
.B2(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_55),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_34),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_49),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_84),
.B(n_23),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_102),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_88),
.A2(n_39),
.B1(n_75),
.B2(n_64),
.Y(n_116)
);

INVxp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_92),
.Y(n_118)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_25),
.A3(n_21),
.B1(n_52),
.B2(n_51),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_68),
.B(n_81),
.C(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_55),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_72),
.Y(n_100)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_34),
.C(n_35),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_62),
.C(n_44),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_14),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_71),
.A2(n_41),
.B1(n_43),
.B2(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_62),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_68),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_119),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_86),
.B(n_91),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_97),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_69),
.B(n_80),
.C(n_62),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_19),
.B(n_48),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_121),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_116),
.B1(n_122),
.B2(n_56),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_73),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_97),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_64),
.C(n_48),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_123),
.C(n_96),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_31),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_48),
.C(n_31),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_96),
.B1(n_103),
.B2(n_86),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_136),
.B1(n_3),
.B2(n_4),
.Y(n_147)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_133),
.Y(n_143)
);

XOR2x2_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_107),
.Y(n_131)
);

AOI221xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_123),
.B1(n_120),
.B2(n_110),
.C(n_117),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_96),
.B1(n_93),
.B2(n_92),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_116),
.B1(n_106),
.B2(n_5),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_93),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_90),
.Y(n_139)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_145),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_150),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_129),
.B1(n_138),
.B2(n_130),
.Y(n_157)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NAND2x1_ASAP7_75t_SL g158 ( 
.A(n_151),
.B(n_132),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_135),
.C(n_127),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_135),
.C(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_133),
.C(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_159),
.B1(n_150),
.B2(n_141),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_137),
.B1(n_12),
.B2(n_13),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_145),
.B(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_164),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_165),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_154),
.B(n_146),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_146),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_153),
.C(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_158),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_15),
.B(n_11),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.C(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_173),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_6),
.C(n_7),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_10),
.B(n_172),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);


endmodule