module fake_jpeg_4082_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx5_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx11_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

OR2x4_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_22),
.Y(n_28)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_17),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_17),
.B(n_13),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_34),
.Y(n_42)
);

AND2x6_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_27),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_16),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_18),
.C(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_49),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_14),
.B1(n_15),
.B2(n_10),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_13),
.B(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_41),
.B1(n_45),
.B2(n_21),
.Y(n_51)
);

OAI22x1_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_55),
.B1(n_25),
.B2(n_20),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_41),
.B1(n_21),
.B2(n_26),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_5),
.C(n_8),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_38),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_SL g59 ( 
.A(n_53),
.B(n_16),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_62),
.C(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_4),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_64),
.A2(n_6),
.B(n_8),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_66),
.C(n_25),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_25),
.C(n_26),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_69),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_2),
.B(n_3),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_70),
.B(n_6),
.Y(n_72)
);

AOI21x1_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_16),
.B(n_12),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_0),
.B(n_14),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_12),
.B(n_1),
.C(n_0),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_14),
.B(n_71),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.C(n_30),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_23),
.B(n_26),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_23),
.Y(n_78)
);


endmodule