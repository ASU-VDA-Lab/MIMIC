module fake_netlist_1_1667_n_18 (n_1, n_2, n_0, n_18);
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
BUFx6f_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
INVx1_ASAP7_75t_L g5 ( .A(n_2), .Y(n_5) );
AOI21xp5_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_3), .B(n_0), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_4), .Y(n_8) );
OAI22xp5_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_5), .B1(n_4), .B2(n_3), .Y(n_9) );
NAND2xp5_ASAP7_75t_L g10 ( .A(n_8), .B(n_4), .Y(n_10) );
AOI211xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_3), .B(n_1), .C(n_2), .Y(n_11) );
OAI221xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_8), .B1(n_3), .B2(n_2), .C(n_1), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_10), .B(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
AOI21xp5_ASAP7_75t_L g16 ( .A1(n_14), .A2(n_3), .B(n_1), .Y(n_16) );
AOI32xp33_ASAP7_75t_L g17 ( .A1(n_15), .A2(n_0), .A3(n_3), .B1(n_12), .B2(n_11), .Y(n_17) );
AOI221xp5_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_0), .B1(n_3), .B2(n_14), .C(n_17), .Y(n_18) );
endmodule