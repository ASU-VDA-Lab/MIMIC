module fake_jpeg_23624_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_4),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx6_ASAP7_75t_SL g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_19),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_24),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_13),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_2),
.B1(n_7),
.B2(n_12),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_16),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_23),
.A2(n_15),
.B(n_9),
.Y(n_34)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_10),
.A2(n_17),
.B1(n_8),
.B2(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_23),
.A2(n_15),
.B1(n_9),
.B2(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_21),
.C(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_21),
.B1(n_34),
.B2(n_31),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_26),
.C(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_46),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_30),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_43),
.C(n_45),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_40),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_33),
.B1(n_42),
.B2(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_53),
.B(n_33),
.Y(n_54)
);


endmodule