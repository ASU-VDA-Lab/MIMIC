module fake_netlist_1_1968_n_714 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_714);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_714;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_529;
wire n_312;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_73), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_23), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_13), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_30), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_45), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_52), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_37), .Y(n_85) );
OR2x2_ASAP7_75t_L g86 ( .A(n_70), .B(n_61), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_78), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_77), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_75), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_60), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_55), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_38), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_41), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_6), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_49), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_48), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_10), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_31), .Y(n_99) );
INVxp33_ASAP7_75t_L g100 ( .A(n_68), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_54), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_3), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_40), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_76), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_7), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_22), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_43), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_65), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_59), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_17), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_28), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_56), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_64), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_7), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_51), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_0), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_62), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_33), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_12), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_25), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_39), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_44), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_35), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_21), .Y(n_126) );
INVx2_ASAP7_75t_SL g127 ( .A(n_67), .Y(n_127) );
INVxp67_ASAP7_75t_L g128 ( .A(n_111), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_102), .Y(n_129) );
AND2x4_ASAP7_75t_SL g130 ( .A(n_99), .B(n_24), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_117), .B(n_0), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_117), .B(n_1), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_87), .A2(n_26), .B(n_72), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_87), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_100), .B(n_1), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_114), .B(n_2), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_88), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_81), .B(n_2), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_113), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_127), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_88), .A2(n_27), .B(n_71), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_81), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_127), .B(n_3), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_91), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
BUFx2_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_85), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_93), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_94), .B(n_4), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_89), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_94), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_96), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_96), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_97), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_97), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_121), .B(n_4), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_79), .B(n_5), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_80), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_83), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_82), .B(n_5), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_104), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_106), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_89), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_108), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_109), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_141), .B(n_107), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_149), .B(n_92), .Y(n_173) );
INVx8_ASAP7_75t_L g174 ( .A(n_139), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_149), .B(n_126), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_141), .B(n_119), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_128), .B(n_112), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_156), .B(n_124), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_164), .B(n_122), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_132), .B(n_95), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_144), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_156), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_129), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_164), .B(n_103), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_135), .A2(n_95), .B1(n_116), .B2(n_120), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
AO221x1_ASAP7_75t_L g195 ( .A1(n_130), .A2(n_116), .B1(n_105), .B2(n_103), .C(n_101), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_156), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_132), .A2(n_98), .B1(n_115), .B2(n_110), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_168), .B(n_115), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_168), .B(n_110), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_135), .B(n_101), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_144), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_156), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_157), .B(n_90), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_138), .B(n_90), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_150), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_153), .A2(n_86), .B(n_123), .C(n_84), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_138), .A2(n_86), .B1(n_9), .B2(n_10), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_169), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_208) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
INVx8_ASAP7_75t_L g210 ( .A(n_136), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_147), .B(n_8), .Y(n_211) );
AOI221xp5_ASAP7_75t_L g212 ( .A1(n_147), .A2(n_11), .B1(n_12), .B2(n_13), .C(n_14), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_154), .B(n_15), .Y(n_213) );
AOI221xp5_ASAP7_75t_L g214 ( .A1(n_154), .A2(n_15), .B1(n_16), .B2(n_18), .C(n_19), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_131), .Y(n_215) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_130), .A2(n_16), .B1(n_20), .B2(n_29), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_158), .B(n_32), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_158), .B(n_34), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_161), .B(n_36), .Y(n_220) );
AND2x2_ASAP7_75t_L g221 ( .A(n_161), .B(n_42), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_150), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_151), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_150), .Y(n_225) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_137), .A2(n_46), .B1(n_47), .B2(n_50), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_165), .B(n_53), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_165), .B(n_57), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_165), .B(n_58), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_171), .B(n_63), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_151), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_171), .B(n_66), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_171), .B(n_74), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_146), .A2(n_148), .B(n_162), .C(n_133), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_151), .B(n_159), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_200), .B(n_145), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_204), .B(n_163), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_174), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_174), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_210), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_191), .B(n_162), .Y(n_242) );
OR2x2_ASAP7_75t_L g243 ( .A(n_215), .B(n_166), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_177), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_198), .B(n_148), .Y(n_246) );
O2A1O1Ixp5_ASAP7_75t_L g247 ( .A1(n_183), .A2(n_152), .B(n_148), .C(n_146), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_177), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_210), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_199), .B(n_130), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_189), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_210), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_194), .B(n_203), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_186), .B(n_160), .Y(n_255) );
OR2x6_ASAP7_75t_L g256 ( .A(n_190), .B(n_142), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
BUFx8_ASAP7_75t_L g258 ( .A(n_186), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_182), .B(n_143), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_172), .B(n_143), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_173), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_175), .B(n_143), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_172), .B(n_143), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_181), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_196), .Y(n_266) );
BUFx12f_ASAP7_75t_L g267 ( .A(n_195), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_202), .A2(n_142), .B(n_134), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_184), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_180), .B(n_133), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_211), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_201), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_180), .B(n_140), .Y(n_273) );
BUFx12f_ASAP7_75t_L g274 ( .A(n_221), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_213), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_183), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_185), .Y(n_277) );
NAND2xp33_ASAP7_75t_L g278 ( .A(n_229), .B(n_151), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_197), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_184), .B(n_140), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_193), .B(n_167), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_193), .B(n_167), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_185), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_235), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g285 ( .A1(n_236), .A2(n_134), .B(n_167), .Y(n_285) );
NOR2x1_ASAP7_75t_L g286 ( .A(n_206), .B(n_167), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
INVxp67_ASAP7_75t_L g288 ( .A(n_218), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_208), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_224), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_176), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_207), .B(n_151), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_224), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_207), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_176), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_218), .B(n_170), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_220), .B(n_170), .Y(n_297) );
NOR3xp33_ASAP7_75t_L g298 ( .A(n_212), .B(n_155), .C(n_159), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g299 ( .A(n_220), .B(n_167), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_179), .Y(n_300) );
OAI22xp33_ASAP7_75t_L g301 ( .A1(n_226), .A2(n_155), .B1(n_159), .B2(n_170), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_217), .B(n_155), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_236), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_227), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_227), .B(n_170), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g306 ( .A(n_253), .B(n_134), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_269), .B(n_214), .Y(n_307) );
INVx1_ASAP7_75t_SL g308 ( .A(n_241), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_269), .B(n_234), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g310 ( .A(n_267), .B(n_230), .Y(n_310) );
NOR2xp33_ASAP7_75t_SL g311 ( .A(n_241), .B(n_234), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_294), .A2(n_167), .B1(n_170), .B2(n_159), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_255), .B(n_262), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_245), .Y(n_314) );
AOI22xp33_ASAP7_75t_SL g315 ( .A1(n_258), .A2(n_134), .B1(n_155), .B2(n_159), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_287), .A2(n_233), .B1(n_231), .B2(n_155), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_279), .A2(n_155), .B1(n_159), .B2(n_170), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_261), .B(n_232), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_253), .B(n_232), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_252), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_249), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_243), .B(n_179), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_250), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_258), .A2(n_209), .B1(n_201), .B2(n_192), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_239), .B(n_187), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_238), .A2(n_187), .B(n_188), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_240), .B(n_228), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_288), .A2(n_188), .B1(n_192), .B2(n_225), .Y(n_329) );
INVx3_ASAP7_75t_SL g330 ( .A(n_292), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_274), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_237), .B(n_205), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_244), .B(n_201), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_263), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_266), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_271), .A2(n_205), .B(n_222), .C(n_223), .Y(n_336) );
NOR3xp33_ASAP7_75t_L g337 ( .A(n_251), .B(n_222), .C(n_223), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_275), .B(n_225), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g339 ( .A(n_298), .B(n_209), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_252), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_289), .B(n_228), .Y(n_341) );
BUFx12f_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_254), .B(n_209), .Y(n_343) );
OAI21xp33_ASAP7_75t_L g344 ( .A1(n_281), .A2(n_209), .B(n_282), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_298), .A2(n_286), .B1(n_254), .B2(n_259), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_246), .A2(n_304), .B(n_288), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_260), .B(n_264), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_259), .B(n_273), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_257), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_265), .B(n_290), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_256), .B(n_247), .C(n_270), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_242), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_284), .A2(n_273), .B1(n_270), .B2(n_276), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_280), .B(n_302), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_278), .A2(n_305), .B(n_268), .Y(n_355) );
AOI21xp33_ASAP7_75t_SL g356 ( .A1(n_301), .A2(n_256), .B(n_303), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_285), .A2(n_247), .B(n_299), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_256), .B(n_302), .Y(n_358) );
OA21x2_ASAP7_75t_L g359 ( .A1(n_344), .A2(n_297), .B(n_296), .Y(n_359) );
OR2x6_ASAP7_75t_L g360 ( .A(n_358), .B(n_299), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_349), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_320), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_335), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_340), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_342), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_357), .A2(n_291), .B(n_300), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_321), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_321), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_352), .A2(n_301), .B1(n_291), .B2(n_300), .Y(n_369) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_344), .A2(n_295), .B(n_277), .Y(n_370) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_321), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_332), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_308), .B(n_290), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_323), .B(n_249), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_306), .A2(n_295), .B(n_283), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_313), .B(n_293), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_347), .B(n_249), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_341), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_314), .Y(n_380) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_356), .A2(n_249), .B(n_272), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_325), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_318), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_354), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_334), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_334), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
OAI21x1_ASAP7_75t_L g388 ( .A1(n_355), .A2(n_272), .B(n_339), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_307), .B(n_272), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_326), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_372), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_372), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_376), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_380), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_380), .B(n_330), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_380), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_388), .A2(n_351), .B(n_327), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_376), .A2(n_348), .B1(n_345), .B2(n_311), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_376), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_378), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_371), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_371), .Y(n_406) );
AO31x2_ASAP7_75t_L g407 ( .A1(n_369), .A2(n_316), .A3(n_317), .B(n_336), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_363), .B(n_353), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_362), .Y(n_409) );
INVxp67_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_371), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_377), .B(n_354), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_371), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVxp67_ASAP7_75t_SL g416 ( .A(n_369), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_377), .B(n_309), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_364), .B(n_358), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_379), .B(n_358), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_394), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_409), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_401), .B(n_364), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_400), .A2(n_360), .B1(n_379), .B2(n_384), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_417), .A2(n_391), .B1(n_360), .B2(n_310), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_401), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_401), .B(n_324), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_409), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_397), .B(n_404), .Y(n_433) );
INVxp67_ASAP7_75t_SL g434 ( .A(n_418), .Y(n_434) );
INVxp67_ASAP7_75t_L g435 ( .A(n_414), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_398), .Y(n_436) );
INVxp33_ASAP7_75t_L g437 ( .A(n_396), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_417), .B(n_382), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_392), .A2(n_360), .B1(n_365), .B2(n_382), .Y(n_440) );
BUFx2_ASAP7_75t_L g441 ( .A(n_406), .Y(n_441) );
OAI211xp5_ASAP7_75t_L g442 ( .A1(n_408), .A2(n_310), .B(n_373), .C(n_365), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_406), .Y(n_443) );
NAND4xp25_ASAP7_75t_L g444 ( .A(n_420), .B(n_315), .C(n_322), .D(n_389), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_412), .A2(n_360), .B1(n_391), .B2(n_337), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_396), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_392), .B(n_364), .Y(n_447) );
AND2x4_ASAP7_75t_L g448 ( .A(n_419), .B(n_381), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_398), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_402), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_393), .B(n_386), .Y(n_451) );
CKINVDCx8_ASAP7_75t_R g452 ( .A(n_411), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_393), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_415), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_412), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_419), .B(n_381), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_426), .B(n_400), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_438), .B(n_402), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_448), .B(n_403), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_436), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_428), .B(n_415), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_422), .Y(n_463) );
INVxp67_ASAP7_75t_L g464 ( .A(n_446), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_422), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_436), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_428), .B(n_415), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_449), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_449), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_442), .B(n_403), .C(n_356), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_404), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_452), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_450), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_426), .B(n_408), .C(n_420), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_433), .B(n_410), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_431), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_428), .B(n_416), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_437), .B(n_410), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_450), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_427), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_455), .B(n_416), .Y(n_481) );
AOI211xp5_ASAP7_75t_L g482 ( .A1(n_424), .A2(n_331), .B(n_343), .C(n_374), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_427), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_453), .Y(n_484) );
INVx1_ASAP7_75t_SL g485 ( .A(n_433), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g486 ( .A(n_441), .B(n_406), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_430), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_440), .A2(n_360), .B1(n_386), .B2(n_385), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_430), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_434), .B(n_411), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_435), .B(n_390), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_432), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_423), .B(n_399), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_432), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_423), .B(n_399), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_445), .A2(n_390), .B1(n_387), .B2(n_385), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_439), .A2(n_381), .B(n_413), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_447), .B(n_390), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_421), .B(n_407), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_451), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_439), .B(n_399), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_451), .B(n_387), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_441), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_439), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_425), .B(n_387), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_459), .B(n_456), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_485), .B(n_454), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_484), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_480), .Y(n_512) );
OR2x2_ASAP7_75t_L g513 ( .A(n_502), .B(n_456), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_506), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_459), .B(n_494), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_506), .Y(n_516) );
NAND2x1p5_ASAP7_75t_L g517 ( .A(n_472), .B(n_443), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_472), .B(n_454), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_486), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_464), .B(n_454), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_457), .A2(n_456), .B1(n_448), .B2(n_444), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_503), .B(n_456), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_498), .B(n_448), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_458), .B(n_448), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_489), .B(n_443), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g526 ( .A(n_459), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_494), .B(n_443), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_493), .B(n_443), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_471), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_466), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_491), .Y(n_531) );
NOR2x1_ASAP7_75t_L g532 ( .A(n_470), .B(n_429), .Y(n_532) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_490), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_480), .Y(n_534) );
INVxp67_ASAP7_75t_L g535 ( .A(n_471), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_496), .B(n_399), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_483), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_462), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_483), .Y(n_539) );
INVx1_ASAP7_75t_SL g540 ( .A(n_462), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_496), .B(n_399), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_477), .B(n_381), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_477), .B(n_407), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_461), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_487), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_466), .B(n_407), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_502), .B(n_407), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_478), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_487), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_481), .B(n_407), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_467), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_495), .B(n_407), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_468), .B(n_359), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_461), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_468), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g556 ( .A(n_482), .B(n_385), .C(n_386), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_469), .B(n_359), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_469), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_475), .B(n_452), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_473), .B(n_359), .Y(n_560) );
INVxp67_ASAP7_75t_SL g561 ( .A(n_463), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_473), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_460), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_479), .B(n_359), .Y(n_564) );
NOR2xp33_ASAP7_75t_SL g565 ( .A(n_472), .B(n_486), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_463), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_504), .B(n_413), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_465), .B(n_413), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_526), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_511), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_531), .B(n_474), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_556), .A2(n_488), .B1(n_475), .B2(n_505), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_524), .B(n_508), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_521), .A2(n_500), .B1(n_501), .B2(n_497), .C(n_504), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_515), .B(n_486), .Y(n_575) );
NOR2xp67_ASAP7_75t_L g576 ( .A(n_515), .B(n_507), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_509), .B(n_467), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_509), .B(n_507), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_548), .B(n_499), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_530), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_565), .B(n_519), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_529), .B(n_499), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_563), .B(n_492), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_530), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_519), .A2(n_492), .B(n_465), .Y(n_585) );
NAND2xp33_ASAP7_75t_L g586 ( .A(n_517), .B(n_476), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_514), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_512), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_534), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_520), .B(n_476), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_548), .B(n_413), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_535), .B(n_405), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_537), .B(n_405), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_538), .B(n_405), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_539), .B(n_405), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_545), .B(n_388), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_549), .B(n_388), .Y(n_597) );
INVx1_ASAP7_75t_SL g598 ( .A(n_516), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_540), .B(n_411), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_561), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_532), .B(n_411), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_522), .B(n_411), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_558), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_527), .B(n_411), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_544), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_527), .B(n_375), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_517), .B(n_371), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_523), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_525), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_528), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_510), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_566), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_517), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_513), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_513), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_559), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_546), .B(n_370), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_551), .B(n_370), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_570), .Y(n_622) );
NOR3xp33_ASAP7_75t_L g623 ( .A(n_571), .B(n_533), .C(n_518), .Y(n_623) );
NAND3xp33_ASAP7_75t_SL g624 ( .A(n_581), .B(n_518), .C(n_550), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g625 ( .A1(n_581), .A2(n_552), .B(n_550), .C(n_547), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_569), .A2(n_543), .B1(n_547), .B2(n_546), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_576), .B(n_542), .Y(n_627) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_572), .B(n_543), .C(n_542), .D(n_567), .Y(n_628) );
AOI211x1_ASAP7_75t_L g629 ( .A1(n_619), .A2(n_536), .B(n_541), .C(n_567), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_575), .B(n_536), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_610), .A2(n_541), .B1(n_564), .B2(n_553), .C(n_557), .Y(n_631) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_569), .A2(n_568), .B1(n_554), .B2(n_544), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_588), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_611), .B(n_564), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g635 ( .A(n_569), .B(n_554), .Y(n_635) );
XNOR2x2_ASAP7_75t_L g636 ( .A(n_598), .B(n_568), .Y(n_636) );
NAND2xp33_ASAP7_75t_L g637 ( .A(n_572), .B(n_560), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_589), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_612), .B(n_560), .Y(n_639) );
INVxp33_ASAP7_75t_L g640 ( .A(n_579), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g641 ( .A(n_585), .B(n_587), .C(n_579), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_600), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_604), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_617), .B(n_557), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_607), .Y(n_645) );
OAI33xp33_ASAP7_75t_L g646 ( .A1(n_618), .A2(n_329), .A3(n_327), .B1(n_553), .B2(n_367), .B3(n_368), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_580), .Y(n_647) );
NOR3xp33_ASAP7_75t_L g648 ( .A(n_591), .B(n_375), .C(n_312), .Y(n_648) );
AND3x1_ASAP7_75t_L g649 ( .A(n_591), .B(n_312), .C(n_368), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_586), .A2(n_375), .B(n_368), .Y(n_650) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_586), .B(n_367), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_584), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_613), .A2(n_328), .B1(n_350), .B2(n_319), .C(n_333), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_602), .B(n_367), .C(n_370), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_601), .B(n_370), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_573), .B(n_371), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_602), .B(n_366), .C(n_328), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_601), .B(n_366), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_640), .B(n_577), .Y(n_659) );
INVx2_ASAP7_75t_SL g660 ( .A(n_630), .Y(n_660) );
AOI222xp33_ASAP7_75t_L g661 ( .A1(n_637), .A2(n_574), .B1(n_582), .B2(n_578), .C1(n_592), .C2(n_616), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_631), .B(n_614), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_629), .B(n_590), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_626), .B(n_583), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_627), .B(n_605), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_622), .Y(n_666) );
AOI222xp33_ASAP7_75t_L g667 ( .A1(n_624), .A2(n_608), .B1(n_603), .B2(n_593), .C1(n_595), .C2(n_615), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_633), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_628), .B(n_594), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_638), .Y(n_670) );
INVxp67_ASAP7_75t_SL g671 ( .A(n_636), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_641), .A2(n_615), .B(n_603), .C(n_609), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_642), .Y(n_673) );
NAND4xp75_ASAP7_75t_L g674 ( .A(n_649), .B(n_609), .C(n_596), .D(n_597), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g675 ( .A(n_644), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_643), .Y(n_676) );
NOR2x1_ASAP7_75t_L g677 ( .A(n_635), .B(n_606), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_641), .A2(n_599), .B(n_606), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g679 ( .A1(n_625), .A2(n_621), .B(n_620), .C(n_319), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g680 ( .A1(n_632), .A2(n_272), .B1(n_623), .B2(n_645), .C(n_646), .Y(n_680) );
INVx3_ASAP7_75t_SL g681 ( .A(n_647), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_681), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_665), .B(n_623), .Y(n_683) );
NAND2x1p5_ASAP7_75t_L g684 ( .A(n_677), .B(n_651), .Y(n_684) );
NAND4xp25_ASAP7_75t_L g685 ( .A(n_672), .B(n_657), .C(n_656), .D(n_653), .Y(n_685) );
NOR3x1_ASAP7_75t_L g686 ( .A(n_671), .B(n_634), .C(n_639), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_666), .Y(n_687) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_678), .B(n_654), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_660), .B(n_652), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_662), .B(n_657), .Y(n_690) );
AOI221xp5_ASAP7_75t_SL g691 ( .A1(n_671), .A2(n_658), .B1(n_655), .B2(n_650), .C(n_648), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_680), .B(n_648), .C(n_674), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_661), .A2(n_669), .B1(n_667), .B2(n_664), .Y(n_693) );
AND3x4_ASAP7_75t_L g694 ( .A(n_675), .B(n_659), .C(n_680), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_668), .Y(n_695) );
INVxp33_ASAP7_75t_L g696 ( .A(n_694), .Y(n_696) );
NOR2xp33_ASAP7_75t_R g697 ( .A(n_682), .B(n_670), .Y(n_697) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_682), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_689), .Y(n_699) );
OAI321xp33_ASAP7_75t_L g700 ( .A1(n_693), .A2(n_663), .A3(n_673), .B1(n_676), .B2(n_679), .C(n_685), .Y(n_700) );
OA22x2_ASAP7_75t_L g701 ( .A1(n_690), .A2(n_679), .B1(n_683), .B2(n_686), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_691), .B(n_692), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_695), .B(n_687), .Y(n_703) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_702), .B(n_688), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_696), .A2(n_684), .B1(n_687), .B2(n_701), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_698), .B(n_701), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_703), .B(n_699), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_707), .Y(n_708) );
XOR2xp5_ASAP7_75t_L g709 ( .A(n_706), .B(n_697), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_704), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_708), .B(n_705), .Y(n_711) );
XOR2x2_ASAP7_75t_L g712 ( .A(n_709), .B(n_700), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_711), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_712), .B(n_710), .Y(n_714) );
endmodule