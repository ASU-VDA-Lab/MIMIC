module fake_netlist_6_4125_n_188 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_188);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_188;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_160;
wire n_90;
wire n_131;
wire n_105;
wire n_54;
wire n_132;
wire n_102;
wire n_186;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

AO21x2_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_53),
.B(n_37),
.Y(n_57)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_2),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_3),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

OR2x6_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_13),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_4),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_38),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

OR2x6_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_42),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_52),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_47),
.B1(n_46),
.B2(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp67_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_50),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_64),
.B1(n_66),
.B2(n_59),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_59),
.B(n_54),
.C(n_56),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

OAI21x1_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_86),
.B(n_54),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_56),
.B(n_54),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_57),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_57),
.Y(n_98)
);

AO32x2_ASAP7_75t_L g99 ( 
.A1(n_78),
.A2(n_62),
.A3(n_57),
.B1(n_68),
.B2(n_54),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_75),
.B(n_63),
.Y(n_100)
);

OAI21x1_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_69),
.B(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_78),
.B(n_68),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

AOI21x1_ASAP7_75t_SL g104 ( 
.A1(n_97),
.A2(n_81),
.B(n_88),
.Y(n_104)
);

O2A1O1Ixp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_54),
.B(n_86),
.C(n_65),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_83),
.Y(n_106)
);

NOR2xp67_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_86),
.Y(n_107)
);

AOI21x1_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_69),
.B(n_57),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_91),
.Y(n_110)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_68),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_106),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_104),
.B(n_95),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_99),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_100),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_115),
.Y(n_126)
);

NAND2x1p5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_102),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_118),
.Y(n_130)
);

NAND4xp25_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_83),
.C(n_39),
.D(n_45),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_118),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_110),
.B(n_37),
.C(n_117),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_58),
.B(n_71),
.Y(n_134)
);

AOI221xp5_ASAP7_75t_L g135 ( 
.A1(n_131),
.A2(n_71),
.B1(n_39),
.B2(n_45),
.C(n_43),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_78),
.B1(n_43),
.B2(n_68),
.Y(n_136)
);

OAI322xp33_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_62),
.A3(n_126),
.B1(n_80),
.B2(n_77),
.C1(n_129),
.C2(n_128),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_78),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_68),
.B(n_62),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_132),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_132),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

AOI221xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_80),
.B1(n_77),
.B2(n_133),
.C(n_36),
.Y(n_148)
);

NAND4xp25_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_70),
.C(n_85),
.D(n_72),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_96),
.B(n_65),
.Y(n_150)
);

OAI322xp33_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_72),
.A3(n_65),
.B1(n_70),
.B2(n_61),
.C1(n_60),
.C2(n_7),
.Y(n_151)
);

AOI221xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_133),
.B1(n_72),
.B2(n_65),
.C(n_101),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_145),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_7),
.Y(n_155)
);

NOR2xp67_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_72),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_72),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_8),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_60),
.C(n_61),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_152),
.B(n_60),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_153),
.Y(n_162)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_60),
.Y(n_164)
);

OAI211xp5_ASAP7_75t_SL g165 ( 
.A1(n_158),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_165)
);

OR2x6_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_101),
.Y(n_166)
);

NAND4xp75_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_10),
.C(n_11),
.D(n_105),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_12),
.Y(n_168)
);

AND2x4_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_15),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_149),
.C(n_111),
.Y(n_170)
);

NOR2x1p5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_61),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_160),
.A3(n_61),
.B1(n_60),
.B2(n_111),
.C1(n_99),
.C2(n_108),
.Y(n_172)
);

OAI211xp5_ASAP7_75t_SL g173 ( 
.A1(n_162),
.A2(n_160),
.B(n_18),
.C(n_19),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_163),
.Y(n_174)
);

AOI221xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_61),
.B1(n_111),
.B2(n_89),
.C(n_91),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_16),
.Y(n_176)
);

NAND4xp25_ASAP7_75t_L g177 ( 
.A(n_170),
.B(n_111),
.C(n_89),
.D(n_91),
.Y(n_177)
);

OAI31xp33_ASAP7_75t_L g178 ( 
.A1(n_171),
.A2(n_164),
.A3(n_163),
.B(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

AOI211xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_177),
.B(n_173),
.C(n_175),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_166),
.B(n_99),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_61),
.B1(n_107),
.B2(n_108),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_20),
.B(n_25),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_29),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_61),
.B1(n_90),
.B2(n_180),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_90),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_178),
.B(n_181),
.Y(n_187)
);

AOI31xp33_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_186),
.A3(n_184),
.B(n_182),
.Y(n_188)
);


endmodule