module real_jpeg_4013_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_0),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_0),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_0),
.A2(n_181),
.B1(n_251),
.B2(n_254),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_0),
.A2(n_84),
.B1(n_86),
.B2(n_181),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_0),
.A2(n_181),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_1),
.A2(n_58),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_1),
.A2(n_58),
.B1(n_360),
.B2(n_381),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_1),
.A2(n_58),
.B1(n_319),
.B2(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_2),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_2),
.Y(n_218)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_2),
.Y(n_228)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_2),
.Y(n_239)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_3),
.Y(n_127)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_3),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_3),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_3),
.Y(n_354)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_3),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_4),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_4),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_88),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_4),
.A2(n_88),
.B1(n_273),
.B2(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_4),
.A2(n_88),
.B1(n_156),
.B2(n_281),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_5),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_5),
.A2(n_51),
.B1(n_184),
.B2(n_307),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_5),
.A2(n_51),
.B1(n_380),
.B2(n_381),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_5),
.A2(n_51),
.B1(n_393),
.B2(n_396),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_6),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_7),
.A2(n_146),
.B1(n_149),
.B2(n_152),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_7),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_7),
.B(n_167),
.C(n_171),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_7),
.B(n_73),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_7),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_7),
.B(n_118),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_7),
.B(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_9),
.Y(n_523)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_10),
.Y(n_103)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_11),
.A2(n_155),
.B1(n_159),
.B2(n_160),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_11),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_159),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_11),
.A2(n_159),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_11),
.A2(n_159),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_12),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_13),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_13),
.A2(n_93),
.B1(n_105),
.B2(n_120),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_93),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_13),
.A2(n_93),
.B1(n_375),
.B2(n_376),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_14),
.Y(n_115)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_14),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_15),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_15),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_15),
.A2(n_120),
.B1(n_272),
.B2(n_360),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_15),
.A2(n_272),
.B1(n_386),
.B2(n_389),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_L g445 ( 
.A1(n_15),
.A2(n_272),
.B1(n_400),
.B2(n_446),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_16),
.A2(n_165),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_16),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_16),
.A2(n_204),
.B1(n_223),
.B2(n_225),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_16),
.A2(n_204),
.B1(n_279),
.B2(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_16),
.A2(n_55),
.B1(n_204),
.B2(n_400),
.Y(n_419)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_521),
.B(n_524),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_135),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_133),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_131),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_131),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_122),
.C(n_128),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_24),
.A2(n_25),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_59),
.C(n_94),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_26),
.B(n_509),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_45),
.B1(n_52),
.B2(n_54),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_27),
.A2(n_52),
.B1(n_54),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_27),
.A2(n_52),
.B1(n_123),
.B2(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_27),
.A2(n_351),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_27),
.A2(n_36),
.B1(n_398),
.B2(n_419),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_27),
.A2(n_45),
.B1(n_52),
.B2(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_28),
.A2(n_349),
.B(n_350),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_28),
.B(n_352),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_36),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_31),
.Y(n_327)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_36),
.B(n_152),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_36)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_37),
.Y(n_329)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_40),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_40),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_40),
.Y(n_388)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_41),
.Y(n_300)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_43),
.Y(n_279)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_43),
.Y(n_391)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_52),
.A2(n_419),
.B(n_447),
.Y(n_457)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_53),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_53),
.B(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_59),
.A2(n_94),
.B1(n_95),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_59),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_83),
.B1(n_89),
.B2(n_90),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_60),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_60),
.A2(n_89),
.B1(n_297),
.B2(n_357),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_60),
.A2(n_89),
.B1(n_385),
.B2(n_392),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_60),
.A2(n_83),
.B1(n_89),
.B2(n_498),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_66),
.Y(n_260)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_72),
.Y(n_265)
);

INVx6_ASAP7_75t_L g433 ( 
.A(n_72),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_73),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_73),
.A2(n_129),
.B1(n_302),
.B2(n_421),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_73),
.A2(n_129),
.B1(n_429),
.B2(n_430),
.Y(n_428)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_79),
.B2(n_82),
.Y(n_73)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_75),
.Y(n_283)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_79),
.Y(n_381)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_81),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_81),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_81),
.Y(n_360)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_SL g257 ( 
.A1(n_86),
.A2(n_152),
.B(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_89),
.B(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_89),
.A2(n_297),
.B(n_301),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_94),
.A2(n_95),
.B1(n_496),
.B2(n_497),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_94),
.B(n_493),
.C(n_496),
.Y(n_504)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_117),
.B(n_119),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_96),
.A2(n_145),
.B(n_153),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_96),
.A2(n_117),
.B1(n_203),
.B2(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_96),
.A2(n_153),
.B(n_250),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_96),
.A2(n_117),
.B1(n_359),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_97),
.B(n_154),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_97),
.A2(n_118),
.B1(n_379),
.B2(n_382),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_97),
.A2(n_118),
.B1(n_382),
.B2(n_407),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_97),
.A2(n_118),
.B1(n_407),
.B2(n_436),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_98)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_99),
.Y(n_380)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_102),
.Y(n_254)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_103),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_106),
.Y(n_158)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_107),
.A2(n_203),
.B(n_208),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_114),
.B2(n_116),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_113),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_113),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_113),
.Y(n_273)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_114),
.Y(n_216)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_115),
.Y(n_342)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_115),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_117),
.A2(n_208),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_118),
.B(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_119),
.Y(n_436)
);

INVx5_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_122),
.B(n_128),
.Y(n_518)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_127),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_129),
.A2(n_257),
.B(n_261),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_129),
.B(n_302),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_129),
.A2(n_261),
.B(n_460),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_515),
.B(n_520),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_486),
.B(n_512),
.Y(n_136)
);

OAI311xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_363),
.A3(n_462),
.B1(n_480),
.C1(n_481),
.Y(n_137)
);

AOI21x1_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_312),
.B(n_362),
.Y(n_138)
);

AO21x1_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_288),
.B(n_311),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_244),
.B(n_287),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_211),
.B(n_243),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_176),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_143),
.B(n_176),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_162),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_144),
.A2(n_162),
.B1(n_163),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_144),
.Y(n_241)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_152),
.A2(n_186),
.B(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_152),
.B(n_331),
.Y(n_330)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_152),
.A2(n_323),
.B(n_330),
.Y(n_349)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_174),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_200),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_177),
.B(n_201),
.C(n_210),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_186),
.B(n_194),
.Y(n_177)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_178),
.Y(n_235)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_186),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_186),
.A2(n_369),
.B1(n_372),
.B2(n_374),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_186),
.A2(n_227),
.B(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_197),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_187),
.A2(n_269),
.B1(n_306),
.B2(n_309),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_187),
.A2(n_337),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_195),
.Y(n_335)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_198),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_209),
.B2(n_210),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_232),
.B(n_242),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_220),
.B(n_231),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_219),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_218),
.Y(n_373)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_218),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_230),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_230),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_229),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_223),
.Y(n_308)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_224),
.Y(n_377)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_227),
.Y(n_309)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_229),
.A2(n_268),
.B(n_274),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_240),
.Y(n_242)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_246),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_266),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_255),
.B2(n_256),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_255),
.C(n_266),
.Y(n_289)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI32xp33_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_278),
.A3(n_280),
.B1(n_282),
.B2(n_284),
.Y(n_277)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_263),
.B(n_329),
.Y(n_328)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_277),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_277),
.Y(n_294)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_283),
.B(n_285),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_289),
.B(n_290),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_310),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_294),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_304),
.C(n_305),
.Y(n_343)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_300),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_300),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_313),
.B(n_314),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_346),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_343),
.B1(n_344),
.B2(n_345),
.Y(n_315)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_316),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_332),
.B2(n_333),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_318),
.B(n_332),
.Y(n_458)
);

OAI32xp33_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_322),
.A3(n_327),
.B1(n_328),
.B2(n_330),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_326),
.Y(n_331)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_343),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_343),
.B(n_344),
.C(n_346),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_355),
.B2(n_361),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_347),
.B(n_356),
.C(n_358),
.Y(n_471)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_355),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_357),
.Y(n_460)
);

NAND2xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_448),
.Y(n_363)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_364),
.A2(n_448),
.B(n_482),
.C(n_485),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_422),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_365),
.B(n_422),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_404),
.C(n_410),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g461 ( 
.A(n_366),
.B(n_404),
.CI(n_410),
.CON(n_461),
.SN(n_461)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_383),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_384),
.C(n_397),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_378),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_368),
.B(n_378),
.Y(n_454)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_369),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_379),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_397),
.Y(n_383)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx4_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_408),
.Y(n_440)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_408),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_409),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_408),
.A2(n_440),
.B(n_443),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.C(n_420),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_411),
.B(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_412),
.B(n_414),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_417),
.A2(n_418),
.B1(n_420),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_420),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_426),
.C(n_438),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_438),
.B2(n_439),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_434),
.B(n_437),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_435),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_430),
.Y(n_498)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_437),
.B(n_489),
.C(n_491),
.Y(n_511)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_461),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_461),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_454),
.C(n_455),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_450),
.A2(n_451),
.B1(n_454),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_454),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_473),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.C(n_459),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_457),
.B1(n_459),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_459),
.Y(n_468)
);

BUFx24_ASAP7_75t_SL g528 ( 
.A(n_461),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_475),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_464),
.A2(n_483),
.B(n_484),
.Y(n_482)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_472),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_472),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.C(n_471),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_466),
.B(n_478),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_469),
.A2(n_470),
.B1(n_471),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_477),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_501),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g487 ( 
.A(n_488),
.B(n_500),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_500),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_490),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_493),
.B1(n_495),
.B2(n_499),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_493),
.B1(n_507),
.B2(n_508),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_503),
.C(n_507),
.Y(n_519)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_495),
.Y(n_499)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_501),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_511),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_511),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_519),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_516),
.B(n_519),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_518),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx13_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx6_ASAP7_75t_L g525 ( 
.A(n_523),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_526),
.Y(n_524)
);


endmodule