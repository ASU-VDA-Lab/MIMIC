module fake_ibex_1132_n_931 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_931);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_931;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_412;
wire n_457;
wire n_357;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_375;
wire n_317;
wire n_340;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_170;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_262;
wire n_439;
wire n_704;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_397;
wire n_366;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_247;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_116),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_20),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_82),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_16),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_45),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_62),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_41),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_65),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_30),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_73),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_67),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_86),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_39),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_85),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_76),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_121),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_38),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_125),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_100),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_24),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_91),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_3),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_58),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_12),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_150),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_117),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_90),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_54),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_139),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_50),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_69),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_4),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_87),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_109),
.Y(n_217)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_84),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_60),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_66),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_140),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_23),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_92),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_107),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_9),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_51),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_23),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_80),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_22),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_103),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_108),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_144),
.B(n_7),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_127),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_37),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_0),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_27),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_43),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_52),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_158),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_49),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_118),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_68),
.Y(n_247)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_15),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_61),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_72),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_17),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_24),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_28),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_137),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_55),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_22),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_79),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_83),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_9),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_29),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_129),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_48),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_46),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_28),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_35),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_165),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_78),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_94),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_102),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_119),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_63),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_133),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_112),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_12),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_89),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_4),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_32),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_21),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_77),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_93),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_42),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_167),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_191),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_193),
.B(n_0),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_167),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_232),
.B(n_191),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_208),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_184),
.B(n_1),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_195),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_2),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_180),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_195),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_230),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_195),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_195),
.Y(n_300)
);

AOI22x1_ASAP7_75t_SL g301 ( 
.A1(n_215),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_222),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

OA21x2_ASAP7_75t_L g305 ( 
.A1(n_209),
.A2(n_96),
.B(n_164),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_216),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_216),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_168),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_220),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_236),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_172),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_228),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_216),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_238),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_242),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_216),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_169),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_211),
.B(n_13),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_255),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_239),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_255),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_208),
.B(n_14),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_170),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_241),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_265),
.B(n_18),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_250),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_171),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_211),
.B(n_19),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_175),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_215),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_275),
.A2(n_101),
.B(n_163),
.Y(n_338)
);

INVx6_ASAP7_75t_L g339 ( 
.A(n_250),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_250),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_265),
.B(n_25),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_241),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_264),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_44),
.Y(n_345)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_177),
.A2(n_104),
.B(n_162),
.Y(n_346)
);

AND2x4_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_26),
.Y(n_347)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_182),
.A2(n_99),
.B(n_161),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_173),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g350 ( 
.A1(n_183),
.A2(n_98),
.B(n_160),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_276),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_196),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_200),
.A2(n_97),
.B(n_157),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_204),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_210),
.Y(n_356)
);

OA21x2_ASAP7_75t_L g357 ( 
.A1(n_212),
.A2(n_95),
.B(n_155),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_213),
.Y(n_358)
);

AND3x2_ASAP7_75t_L g359 ( 
.A(n_351),
.B(n_248),
.C(n_251),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_290),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_339),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_339),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g364 ( 
.A1(n_296),
.A2(n_302),
.B1(n_328),
.B2(n_313),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_343),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_281),
.B1(n_282),
.B2(n_190),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_324),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_192),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_321),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_294),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_312),
.B(n_178),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_321),
.A2(n_276),
.B1(n_282),
.B2(n_268),
.Y(n_374)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_312),
.B(n_186),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_294),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_297),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_297),
.Y(n_379)
);

BUFx8_ASAP7_75t_SL g380 ( 
.A(n_331),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_290),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_333),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_297),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_326),
.B(n_329),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_312),
.B(n_192),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_318),
.B(n_331),
.Y(n_389)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_345),
.Y(n_390)
);

BUFx6f_ASAP7_75t_SL g391 ( 
.A(n_326),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_326),
.B(n_214),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_318),
.B(n_226),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_299),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_299),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_290),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_299),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_299),
.Y(n_400)
);

AND2x6_ASAP7_75t_SL g401 ( 
.A(n_288),
.B(n_185),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_299),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_300),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_318),
.B(n_217),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_300),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_331),
.B(n_271),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_300),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_300),
.Y(n_409)
);

NAND3xp33_ASAP7_75t_L g410 ( 
.A(n_286),
.B(n_189),
.C(n_176),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_300),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_345),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_306),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_306),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_329),
.B(n_221),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_341),
.B(n_271),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_306),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_310),
.A2(n_223),
.B1(n_201),
.B2(n_280),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_306),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_306),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_342),
.B(n_347),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_342),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_307),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_347),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_307),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_347),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_307),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_310),
.B(n_224),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_339),
.A2(n_281),
.B1(n_266),
.B2(n_279),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_341),
.B(n_217),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_341),
.Y(n_434)
);

NAND3xp33_ASAP7_75t_L g435 ( 
.A(n_295),
.B(n_252),
.C(n_227),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_320),
.B(n_261),
.C(n_260),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_320),
.B(n_274),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_285),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_307),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_289),
.Y(n_440)
);

INVx2_ASAP7_75t_SL g441 ( 
.A(n_291),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_327),
.B(n_283),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_304),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_332),
.A2(n_253),
.B1(n_203),
.B2(n_263),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_334),
.B(n_283),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_334),
.B(n_225),
.Y(n_446)
);

AO22x2_ASAP7_75t_L g447 ( 
.A1(n_301),
.A2(n_235),
.B1(n_205),
.B2(n_198),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_355),
.B(n_229),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_355),
.B(n_174),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_308),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_308),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_315),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_301),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_315),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_356),
.A2(n_166),
.B1(n_247),
.B2(n_268),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_311),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_353),
.B(n_267),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_319),
.Y(n_458)
);

BUFx2_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_353),
.B(n_243),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_314),
.Y(n_461)
);

NOR2x1p5_ASAP7_75t_L g462 ( 
.A(n_287),
.B(n_194),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_316),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_319),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_293),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_369),
.A2(n_166),
.B1(n_190),
.B2(n_247),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_375),
.B(n_179),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_365),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_384),
.B(n_316),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_375),
.B(n_181),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_394),
.B(n_317),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_462),
.A2(n_323),
.B1(n_335),
.B2(n_317),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_389),
.B(n_287),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_442),
.B(n_292),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_292),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_369),
.A2(n_325),
.B1(n_335),
.B2(n_323),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_375),
.B(n_187),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_298),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_374),
.B(n_432),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_373),
.B(n_303),
.Y(n_482)
);

BUFx5_ASAP7_75t_L g483 ( 
.A(n_412),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_373),
.B(n_303),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_397),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_423),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_434),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_380),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_459),
.B(n_309),
.Y(n_489)
);

O2A1O1Ixp5_ASAP7_75t_L g490 ( 
.A1(n_387),
.A2(n_218),
.B(n_258),
.C(n_256),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_433),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_412),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_380),
.Y(n_493)
);

AND2x6_ASAP7_75t_SL g494 ( 
.A(n_453),
.B(n_309),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_376),
.B(n_206),
.Y(n_495)
);

NOR3xp33_ASAP7_75t_L g496 ( 
.A(n_366),
.B(n_246),
.C(n_245),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_437),
.B(n_325),
.Y(n_497)
);

BUFx6f_ASAP7_75t_SL g498 ( 
.A(n_367),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_376),
.B(n_188),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_425),
.B(n_340),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_438),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_393),
.B(n_197),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_375),
.B(n_199),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_407),
.B(n_202),
.Y(n_504)
);

OR2x6_ASAP7_75t_L g505 ( 
.A(n_447),
.B(n_348),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_L g506 ( 
.A(n_410),
.B(n_340),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_418),
.B(n_207),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_438),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_360),
.B(n_233),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_457),
.B(n_234),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_362),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_440),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_383),
.B(n_240),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_420),
.B(n_305),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_363),
.Y(n_516)
);

AND2x6_ASAP7_75t_SL g517 ( 
.A(n_447),
.B(n_460),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_427),
.B(n_305),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_429),
.B(n_305),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_432),
.B(n_364),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_449),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_390),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_390),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_447),
.B(n_350),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_383),
.B(n_244),
.Y(n_525)
);

AND2x6_ASAP7_75t_SL g526 ( 
.A(n_460),
.B(n_231),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_440),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_381),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_435),
.B(n_254),
.Y(n_529)
);

BUFx8_ASAP7_75t_L g530 ( 
.A(n_391),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_401),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_436),
.B(n_354),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_392),
.B(n_249),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_406),
.B(n_259),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_416),
.B(n_262),
.Y(n_535)
);

BUFx6f_ASAP7_75t_SL g536 ( 
.A(n_441),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_359),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_416),
.Y(n_539)
);

AND2x6_ASAP7_75t_SL g540 ( 
.A(n_448),
.B(n_231),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_424),
.A2(n_417),
.B1(n_368),
.B2(n_431),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_417),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

O2A1O1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_364),
.A2(n_269),
.B(n_273),
.C(n_277),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_456),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_446),
.B(n_338),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_368),
.A2(n_357),
.B1(n_346),
.B2(n_354),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_461),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_463),
.B(n_346),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_420),
.B(n_357),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_444),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_467),
.B(n_444),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_473),
.B(n_486),
.Y(n_555)
);

BUFx4f_ASAP7_75t_L g556 ( 
.A(n_505),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_548),
.A2(n_464),
.B(n_458),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_547),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g559 ( 
.A(n_549),
.B(n_474),
.C(n_552),
.Y(n_559)
);

NAND2x1p5_ASAP7_75t_L g560 ( 
.A(n_538),
.B(n_330),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_470),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_470),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_518),
.A2(n_454),
.B(n_452),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_491),
.B(n_31),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g565 ( 
.A(n_488),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_539),
.B(n_32),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_530),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_492),
.B(n_322),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_482),
.B(n_33),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_481),
.B(n_33),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_498),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_489),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_553),
.A2(n_322),
.B1(n_337),
.B2(n_344),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_519),
.A2(n_439),
.B(n_430),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_SL g575 ( 
.A1(n_519),
.A2(n_428),
.B(n_426),
.C(n_422),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_472),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_520),
.A2(n_337),
.B1(n_344),
.B2(n_422),
.Y(n_577)
);

AOI21xp33_ASAP7_75t_L g578 ( 
.A1(n_495),
.A2(n_529),
.B(n_521),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_506),
.B(n_34),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

AOI33xp33_ASAP7_75t_L g581 ( 
.A1(n_544),
.A2(n_428),
.A3(n_426),
.B1(n_421),
.B2(n_419),
.B3(n_415),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_496),
.A2(n_337),
.B1(n_344),
.B2(n_415),
.Y(n_582)
);

A2O1A1Ixp33_ASAP7_75t_L g583 ( 
.A1(n_484),
.A2(n_344),
.B(n_411),
.C(n_409),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_541),
.A2(n_414),
.B1(n_411),
.B2(n_409),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_500),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_537),
.B(n_35),
.Y(n_586)
);

BUFx4f_ASAP7_75t_L g587 ( 
.A(n_505),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_499),
.B(n_36),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_487),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_485),
.B(n_36),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_502),
.B(n_37),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_551),
.A2(n_385),
.B(n_405),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_480),
.A2(n_382),
.B1(n_403),
.B2(n_402),
.Y(n_594)
);

AO21x1_ASAP7_75t_L g595 ( 
.A1(n_532),
.A2(n_379),
.B(n_402),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_533),
.B(n_497),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_531),
.A2(n_39),
.B1(n_400),
.B2(n_396),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_492),
.B(n_361),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_515),
.B(n_370),
.Y(n_599)
);

OAI22xp33_ASAP7_75t_L g600 ( 
.A1(n_524),
.A2(n_493),
.B1(n_465),
.B2(n_535),
.Y(n_600)
);

O2A1O1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_475),
.A2(n_476),
.B(n_477),
.C(n_524),
.Y(n_601)
);

BUFx12f_ASAP7_75t_L g602 ( 
.A(n_530),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_466),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g604 ( 
.A1(n_490),
.A2(n_378),
.B(n_371),
.C(n_396),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_532),
.B(n_361),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_543),
.B(n_53),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_534),
.A2(n_386),
.B(n_372),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_L g608 ( 
.A(n_493),
.B(n_386),
.C(n_372),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_545),
.B(n_56),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_524),
.A2(n_408),
.B1(n_398),
.B2(n_395),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_504),
.A2(n_408),
.B(n_398),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_546),
.B(n_57),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_483),
.B(n_507),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_511),
.A2(n_377),
.B(n_361),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_550),
.A2(n_377),
.B1(n_64),
.B2(n_71),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_514),
.A2(n_59),
.B(n_74),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_501),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_512),
.B(n_75),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_468),
.A2(n_479),
.B(n_503),
.Y(n_619)
);

BUFx8_ASAP7_75t_L g620 ( 
.A(n_536),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_152),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_508),
.Y(n_622)
);

CKINVDCx10_ASAP7_75t_R g623 ( 
.A(n_536),
.Y(n_623)
);

BUFx8_ASAP7_75t_L g624 ( 
.A(n_516),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_572),
.B(n_540),
.Y(n_625)
);

CKINVDCx8_ASAP7_75t_R g626 ( 
.A(n_623),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_575),
.A2(n_471),
.B(n_525),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_561),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_562),
.Y(n_629)
);

NAND2x1p5_ASAP7_75t_L g630 ( 
.A(n_567),
.B(n_528),
.Y(n_630)
);

AO31x2_ASAP7_75t_L g631 ( 
.A1(n_595),
.A2(n_527),
.A3(n_513),
.B(n_526),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_618),
.A2(n_523),
.B(n_522),
.Y(n_632)
);

A2O1A1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_576),
.A2(n_523),
.B(n_522),
.C(n_509),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_572),
.B(n_517),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_580),
.A2(n_522),
.B(n_509),
.C(n_483),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_602),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_620),
.Y(n_637)
);

AOI31xp67_ASAP7_75t_L g638 ( 
.A1(n_605),
.A2(n_621),
.A3(n_609),
.B(n_606),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_556),
.Y(n_639)
);

BUFx12f_ASAP7_75t_L g640 ( 
.A(n_620),
.Y(n_640)
);

A2O1A1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_589),
.A2(n_483),
.B(n_494),
.C(n_88),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_603),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_585),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_624),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_554),
.B(n_122),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_SL g646 ( 
.A1(n_613),
.A2(n_124),
.B(n_126),
.C(n_128),
.Y(n_646)
);

BUFx10_ASAP7_75t_L g647 ( 
.A(n_571),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_557),
.A2(n_131),
.B(n_132),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_570),
.B(n_135),
.Y(n_649)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_596),
.A2(n_611),
.B(n_614),
.Y(n_650)
);

BUFx6f_ASAP7_75t_SL g651 ( 
.A(n_618),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_555),
.B(n_142),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_564),
.Y(n_654)
);

A2O1A1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_592),
.A2(n_143),
.B(n_145),
.C(n_149),
.Y(n_655)
);

AOI211x1_ASAP7_75t_L g656 ( 
.A1(n_578),
.A2(n_151),
.B(n_600),
.C(n_569),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_617),
.Y(n_657)
);

BUFx2_ASAP7_75t_L g658 ( 
.A(n_618),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_558),
.B(n_588),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_566),
.B(n_622),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_563),
.A2(n_574),
.B(n_593),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_624),
.B(n_581),
.Y(n_662)
);

INVx4_ASAP7_75t_L g663 ( 
.A(n_560),
.Y(n_663)
);

INVxp67_ASAP7_75t_SL g664 ( 
.A(n_556),
.Y(n_664)
);

BUFx2_ASAP7_75t_L g665 ( 
.A(n_560),
.Y(n_665)
);

CKINVDCx11_ASAP7_75t_R g666 ( 
.A(n_565),
.Y(n_666)
);

AO31x2_ASAP7_75t_L g667 ( 
.A1(n_577),
.A2(n_583),
.A3(n_573),
.B(n_604),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_590),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_587),
.A2(n_612),
.B1(n_582),
.B2(n_579),
.Y(n_669)
);

AO31x2_ASAP7_75t_L g670 ( 
.A1(n_615),
.A2(n_616),
.A3(n_584),
.B(n_594),
.Y(n_670)
);

INVxp67_ASAP7_75t_SL g671 ( 
.A(n_597),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_586),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_599),
.B(n_608),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_619),
.A2(n_598),
.B(n_607),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_599),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_556),
.Y(n_677)
);

OAI22x1_ASAP7_75t_L g678 ( 
.A1(n_567),
.A2(n_467),
.B1(n_374),
.B2(n_469),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_561),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_554),
.B(n_481),
.Y(n_680)
);

BUFx10_ASAP7_75t_L g681 ( 
.A(n_618),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_561),
.A2(n_562),
.B1(n_580),
.B2(n_576),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_572),
.B(n_469),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_572),
.B(n_561),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_SL g685 ( 
.A1(n_572),
.A2(n_455),
.B(n_467),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g686 ( 
.A1(n_575),
.A2(n_519),
.B(n_518),
.Y(n_686)
);

OAI21xp33_ASAP7_75t_L g687 ( 
.A1(n_596),
.A2(n_365),
.B(n_469),
.Y(n_687)
);

AO31x2_ASAP7_75t_L g688 ( 
.A1(n_595),
.A2(n_577),
.A3(n_610),
.B(n_583),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_572),
.B(n_554),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_561),
.B(n_562),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_554),
.B(n_481),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_572),
.B(n_561),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_602),
.B(n_469),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_572),
.B(n_561),
.Y(n_694)
);

A2O1A1Ixp33_ASAP7_75t_L g695 ( 
.A1(n_601),
.A2(n_562),
.B(n_576),
.C(n_561),
.Y(n_695)
);

AO31x2_ASAP7_75t_L g696 ( 
.A1(n_595),
.A2(n_577),
.A3(n_610),
.B(n_583),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_572),
.B(n_561),
.Y(n_697)
);

AO32x2_ASAP7_75t_L g698 ( 
.A1(n_577),
.A2(n_478),
.A3(n_573),
.B1(n_610),
.B2(n_597),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_561),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_554),
.B(n_481),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_572),
.B(n_561),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_572),
.B(n_469),
.Y(n_702)
);

AO31x2_ASAP7_75t_L g703 ( 
.A1(n_595),
.A2(n_577),
.A3(n_610),
.B(n_583),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_570),
.A2(n_455),
.B1(n_478),
.B2(n_520),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_699),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_684),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_692),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_690),
.B(n_694),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_697),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_628),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_661),
.A2(n_650),
.B(n_686),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_644),
.Y(n_712)
);

NAND2x1p5_ASAP7_75t_L g713 ( 
.A(n_639),
.B(n_677),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_701),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_629),
.B(n_679),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_690),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_690),
.B(n_664),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_680),
.B(n_691),
.Y(n_718)
);

AO31x2_ASAP7_75t_L g719 ( 
.A1(n_635),
.A2(n_633),
.A3(n_682),
.B(n_674),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_636),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_642),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_685),
.B(n_625),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_657),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_653),
.A2(n_700),
.B(n_627),
.Y(n_724)
);

AO31x2_ASAP7_75t_L g725 ( 
.A1(n_648),
.A2(n_655),
.A3(n_669),
.B(n_673),
.Y(n_725)
);

OAI21xp5_ASAP7_75t_L g726 ( 
.A1(n_660),
.A2(n_649),
.B(n_654),
.Y(n_726)
);

AO31x2_ASAP7_75t_L g727 ( 
.A1(n_643),
.A2(n_675),
.A3(n_656),
.B(n_641),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_658),
.B(n_681),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_704),
.A2(n_651),
.B1(n_632),
.B2(n_689),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_704),
.A2(n_671),
.B1(n_645),
.B2(n_678),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_659),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_662),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_668),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_683),
.B(n_702),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_687),
.B(n_634),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_681),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_663),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_672),
.B(n_652),
.Y(n_738)
);

NAND2x1p5_ASAP7_75t_L g739 ( 
.A(n_639),
.B(n_677),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_665),
.B(n_630),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_639),
.B(n_677),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_631),
.Y(n_742)
);

INVx6_ASAP7_75t_L g743 ( 
.A(n_636),
.Y(n_743)
);

OA21x2_ASAP7_75t_L g744 ( 
.A1(n_638),
.A2(n_703),
.B(n_688),
.Y(n_744)
);

OR2x6_ASAP7_75t_L g745 ( 
.A(n_640),
.B(n_693),
.Y(n_745)
);

NAND2x1p5_ASAP7_75t_L g746 ( 
.A(n_636),
.B(n_637),
.Y(n_746)
);

AO31x2_ASAP7_75t_L g747 ( 
.A1(n_667),
.A2(n_703),
.A3(n_696),
.B(n_688),
.Y(n_747)
);

NOR2xp67_ASAP7_75t_L g748 ( 
.A(n_626),
.B(n_666),
.Y(n_748)
);

AOI21x1_ASAP7_75t_L g749 ( 
.A1(n_698),
.A2(n_631),
.B(n_670),
.Y(n_749)
);

OA21x2_ASAP7_75t_L g750 ( 
.A1(n_670),
.A2(n_631),
.B(n_698),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_646),
.A2(n_676),
.B(n_647),
.Y(n_751)
);

BUFx12f_ASAP7_75t_L g752 ( 
.A(n_676),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_684),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_695),
.A2(n_559),
.B(n_686),
.Y(n_754)
);

BUFx4f_ASAP7_75t_SL g755 ( 
.A(n_640),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_644),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_682),
.A2(n_704),
.B1(n_587),
.B2(n_556),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_689),
.B(n_572),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_690),
.B(n_684),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_685),
.B(n_520),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_628),
.B(n_561),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_695),
.A2(n_559),
.B(n_686),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_682),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_644),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_644),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_685),
.B(n_520),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_682),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_689),
.B(n_572),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_682),
.A2(n_704),
.B1(n_587),
.B2(n_556),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_695),
.A2(n_559),
.B(n_686),
.Y(n_770)
);

HB1xp67_ASAP7_75t_L g771 ( 
.A(n_682),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_684),
.Y(n_772)
);

NAND2x1p5_ASAP7_75t_L g773 ( 
.A(n_639),
.B(n_677),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_753),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_753),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_706),
.B(n_707),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_760),
.B(n_766),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_716),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_763),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_760),
.B(n_766),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_763),
.A2(n_767),
.B1(n_771),
.B2(n_730),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_743),
.Y(n_782)
);

AO21x2_ASAP7_75t_L g783 ( 
.A1(n_711),
.A2(n_770),
.B(n_754),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_715),
.Y(n_784)
);

INVxp67_ASAP7_75t_L g785 ( 
.A(n_765),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_740),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_709),
.B(n_714),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_708),
.B(n_759),
.Y(n_788)
);

INVx2_ASAP7_75t_SL g789 ( 
.A(n_743),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_742),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_772),
.B(n_758),
.Y(n_791)
);

OA21x2_ASAP7_75t_L g792 ( 
.A1(n_754),
.A2(n_770),
.B(n_762),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_710),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_721),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_768),
.B(n_705),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_761),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_740),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_722),
.A2(n_730),
.B1(n_732),
.B2(n_769),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_723),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_734),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_755),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_724),
.B(n_731),
.Y(n_802)
);

AO31x2_ASAP7_75t_L g803 ( 
.A1(n_757),
.A2(n_769),
.A3(n_722),
.B(n_729),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_743),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_718),
.B(n_735),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_767),
.Y(n_806)
);

INVxp33_ASAP7_75t_SL g807 ( 
.A(n_748),
.Y(n_807)
);

OR2x2_ASAP7_75t_L g808 ( 
.A(n_718),
.B(n_750),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_717),
.B(n_737),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_719),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_726),
.B(n_749),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_737),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_752),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_747),
.B(n_738),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_790),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_777),
.A2(n_729),
.B1(n_738),
.B2(n_728),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_802),
.B(n_747),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_814),
.B(n_744),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_808),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_779),
.Y(n_820)
);

OAI22xp33_ASAP7_75t_L g821 ( 
.A1(n_796),
.A2(n_755),
.B1(n_745),
.B2(n_728),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_780),
.A2(n_798),
.B1(n_805),
.B2(n_781),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_795),
.B(n_725),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_806),
.B(n_736),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_811),
.B(n_725),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_791),
.B(n_719),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_811),
.B(n_792),
.Y(n_827)
);

OAI211xp5_ASAP7_75t_L g828 ( 
.A1(n_812),
.A2(n_720),
.B(n_741),
.C(n_712),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_774),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_775),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_799),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_791),
.B(n_727),
.Y(n_832)
);

NOR2x1_ASAP7_75t_L g833 ( 
.A(n_778),
.B(n_745),
.Y(n_833)
);

INVx3_ASAP7_75t_SL g834 ( 
.A(n_813),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_809),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_785),
.B(n_764),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_803),
.B(n_733),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_831),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_815),
.Y(n_839)
);

AND2x4_ASAP7_75t_SL g840 ( 
.A(n_835),
.B(n_788),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_831),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_826),
.B(n_803),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_826),
.B(n_803),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_822),
.B(n_784),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_836),
.B(n_756),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_827),
.B(n_810),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_820),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_817),
.B(n_783),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_820),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_827),
.B(n_810),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_827),
.B(n_783),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_823),
.B(n_783),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_823),
.B(n_792),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_829),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_829),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_838),
.B(n_830),
.Y(n_856)
);

INVxp67_ASAP7_75t_SL g857 ( 
.A(n_841),
.Y(n_857)
);

OR2x2_ASAP7_75t_L g858 ( 
.A(n_848),
.B(n_819),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_851),
.B(n_853),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_847),
.Y(n_860)
);

OAI21xp5_ASAP7_75t_SL g861 ( 
.A1(n_840),
.A2(n_821),
.B(n_828),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_839),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_851),
.B(n_825),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_853),
.B(n_852),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_852),
.B(n_825),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_839),
.Y(n_866)
);

OAI22xp33_ASAP7_75t_SL g867 ( 
.A1(n_854),
.A2(n_830),
.B1(n_834),
.B2(n_835),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_846),
.B(n_818),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_855),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_859),
.B(n_850),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_869),
.Y(n_871)
);

AND2x4_ASAP7_75t_SL g872 ( 
.A(n_868),
.B(n_835),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_862),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_864),
.B(n_842),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_862),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_856),
.B(n_847),
.C(n_849),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_859),
.B(n_850),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_857),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_864),
.B(n_844),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_865),
.B(n_842),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_866),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_879),
.A2(n_861),
.B1(n_821),
.B2(n_816),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_873),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_879),
.B(n_865),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_875),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_872),
.Y(n_886)
);

AOI21xp33_ASAP7_75t_SL g887 ( 
.A1(n_876),
.A2(n_834),
.B(n_867),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_881),
.Y(n_888)
);

NAND2x1p5_ASAP7_75t_L g889 ( 
.A(n_872),
.B(n_813),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_871),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_878),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_870),
.B(n_863),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_882),
.A2(n_877),
.B1(n_870),
.B2(n_863),
.Y(n_893)
);

OAI22xp33_ASAP7_75t_L g894 ( 
.A1(n_886),
.A2(n_874),
.B1(n_880),
.B2(n_860),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_882),
.A2(n_843),
.B1(n_837),
.B2(n_832),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_889),
.A2(n_877),
.B1(n_840),
.B2(n_843),
.Y(n_896)
);

NAND4xp75_ASAP7_75t_L g897 ( 
.A(n_893),
.B(n_833),
.C(n_891),
.D(n_845),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_894),
.A2(n_887),
.B(n_828),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_896),
.A2(n_884),
.B1(n_892),
.B2(n_890),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_899),
.B(n_895),
.Y(n_900)
);

OAI211xp5_ASAP7_75t_L g901 ( 
.A1(n_898),
.A2(n_801),
.B(n_813),
.C(n_816),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_900),
.Y(n_902)
);

NAND3x1_ASAP7_75t_L g903 ( 
.A(n_901),
.B(n_833),
.C(n_897),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_902),
.Y(n_904)
);

NOR2x1_ASAP7_75t_L g905 ( 
.A(n_903),
.B(n_745),
.Y(n_905)
);

XNOR2xp5_ASAP7_75t_L g906 ( 
.A(n_905),
.B(n_807),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_904),
.B(n_883),
.Y(n_907)
);

OAI21x1_ASAP7_75t_L g908 ( 
.A1(n_906),
.A2(n_746),
.B(n_739),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_907),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_906),
.A2(n_746),
.B(n_813),
.Y(n_910)
);

OAI221xp5_ASAP7_75t_L g911 ( 
.A1(n_910),
.A2(n_813),
.B1(n_782),
.B2(n_789),
.C(n_804),
.Y(n_911)
);

OAI22xp5_ASAP7_75t_L g912 ( 
.A1(n_909),
.A2(n_813),
.B1(n_822),
.B2(n_888),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_908),
.B(n_885),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_L g914 ( 
.A1(n_909),
.A2(n_800),
.B1(n_860),
.B2(n_824),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_909),
.Y(n_915)
);

OAI21x1_ASAP7_75t_SL g916 ( 
.A1(n_913),
.A2(n_789),
.B(n_782),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_SL g917 ( 
.A1(n_915),
.A2(n_713),
.B1(n_773),
.B2(n_739),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_914),
.Y(n_918)
);

OAI22x1_ASAP7_75t_L g919 ( 
.A1(n_911),
.A2(n_713),
.B1(n_773),
.B2(n_804),
.Y(n_919)
);

AO21x2_ASAP7_75t_L g920 ( 
.A1(n_912),
.A2(n_751),
.B(n_797),
.Y(n_920)
);

AOI221xp5_ASAP7_75t_L g921 ( 
.A1(n_915),
.A2(n_786),
.B1(n_793),
.B2(n_794),
.C(n_787),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_915),
.B(n_858),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_921),
.B(n_787),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_918),
.A2(n_837),
.B1(n_809),
.B2(n_794),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_922),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_917),
.Y(n_926)
);

OAI21xp33_ASAP7_75t_L g927 ( 
.A1(n_925),
.A2(n_919),
.B(n_916),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_926),
.B(n_920),
.Y(n_928)
);

OAI21x1_ASAP7_75t_L g929 ( 
.A1(n_923),
.A2(n_751),
.B(n_776),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_928),
.A2(n_924),
.B(n_776),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_930),
.A2(n_927),
.B1(n_929),
.B2(n_778),
.Y(n_931)
);


endmodule