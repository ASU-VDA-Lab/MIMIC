module real_jpeg_17463_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_0),
.Y(n_127)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_0),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_0),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_1),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_2),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g266 ( 
.A1(n_2),
.A2(n_121),
.B1(n_267),
.B2(n_270),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_2),
.A2(n_121),
.B1(n_396),
.B2(n_398),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_2),
.A2(n_121),
.B1(n_361),
.B2(n_463),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_3),
.A2(n_157),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_165),
.B1(n_259),
.B2(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_3),
.A2(n_165),
.B1(n_302),
.B2(n_305),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_3),
.A2(n_165),
.B1(n_386),
.B2(n_390),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_204),
.B1(n_207),
.B2(n_211),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_4),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_4),
.A2(n_211),
.B1(n_442),
.B2(n_445),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g504 ( 
.A1(n_4),
.A2(n_25),
.B1(n_211),
.B2(n_505),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_5),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_5),
.Y(n_202)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_5),
.Y(n_295)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_6),
.A2(n_25),
.A3(n_29),
.B1(n_35),
.B2(n_40),
.Y(n_24)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_39),
.B1(n_150),
.B2(n_156),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_6),
.B(n_188),
.Y(n_187)
);

NAND2xp33_ASAP7_75t_SL g277 ( 
.A(n_6),
.B(n_124),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_6),
.B(n_74),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_6),
.B(n_257),
.Y(n_318)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_6),
.A2(n_349),
.A3(n_352),
.B1(n_356),
.B2(n_360),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_6),
.A2(n_39),
.B1(n_377),
.B2(n_381),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_7),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_7),
.A2(n_67),
.B1(n_174),
.B2(n_178),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_7),
.A2(n_67),
.B1(n_429),
.B2(n_432),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_7),
.A2(n_67),
.B1(n_381),
.B2(n_510),
.Y(n_509)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_8),
.Y(n_97)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_8),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_8),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_8),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_9),
.A2(n_80),
.B1(n_404),
.B2(n_405),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_9),
.A2(n_80),
.B1(n_468),
.B2(n_471),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_10),
.A2(n_106),
.B1(n_112),
.B2(n_113),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_10),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_10),
.A2(n_112),
.B1(n_215),
.B2(n_221),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_10),
.A2(n_112),
.B1(n_283),
.B2(n_286),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_10),
.A2(n_112),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_11),
.A2(n_342),
.B1(n_345),
.B2(n_347),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_11),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_11),
.A2(n_347),
.B1(n_445),
.B2(n_454),
.Y(n_453)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_12),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_12),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_13),
.Y(n_143)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g79 ( 
.A(n_14),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g355 ( 
.A(n_15),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_15),
.Y(n_373)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_15),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_485),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_410),
.B(n_481),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_328),
.B(n_409),
.Y(n_19)
);

AOI21x1_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_227),
.B(n_327),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_167),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_22),
.B(n_167),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_83),
.C(n_122),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_23),
.B(n_324),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_24),
.B(n_50),
.Y(n_169)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g506 ( 
.A(n_27),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_28),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_28),
.Y(n_470)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_28),
.Y(n_475)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_33),
.Y(n_261)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_34),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_34),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_38),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_39),
.B(n_247),
.Y(n_246)
);

OAI21xp33_ASAP7_75t_SL g254 ( 
.A1(n_39),
.A2(n_246),
.B(n_255),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_39),
.A2(n_52),
.B1(n_74),
.B2(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_39),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_45),
.Y(n_193)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_62),
.B(n_71),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_51),
.A2(n_281),
.B1(n_291),
.B2(n_292),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_51),
.A2(n_203),
.B1(n_337),
.B2(n_341),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_51),
.A2(n_71),
.B(n_341),
.Y(n_437)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_52),
.B(n_76),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_52),
.A2(n_266),
.B(n_273),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_52),
.A2(n_282),
.B1(n_301),
.B2(n_316),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_52),
.A2(n_63),
.B(n_493),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_55),
.Y(n_285)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_56),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_57),
.Y(n_290)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_58),
.Y(n_317)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_63),
.B(n_200),
.Y(n_274)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_66),
.Y(n_240)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_66),
.Y(n_304)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_66),
.Y(n_313)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_70),
.Y(n_210)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_70),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_79),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_79),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_82),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_83),
.B(n_122),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_98),
.B1(n_104),
.B2(n_115),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g401 ( 
.A1(n_84),
.A2(n_173),
.B(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_84),
.A2(n_98),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g497 ( 
.A1(n_84),
.A2(n_402),
.B(n_453),
.Y(n_497)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_85),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_85),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_85),
.A2(n_105),
.B1(n_257),
.B2(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_85),
.B(n_403),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_98),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_89),
.B1(n_91),
.B2(n_95),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_87),
.Y(n_248)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

AO22x2_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_125),
.B1(n_128),
.B2(n_131),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_97),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_98),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_98),
.Y(n_257)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_114),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_149),
.B1(n_163),
.B2(n_166),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_123),
.A2(n_163),
.B1(n_166),
.B2(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_123),
.A2(n_166),
.B1(n_214),
.B2(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_123),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_123),
.A2(n_428),
.B(n_466),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_123),
.A2(n_166),
.B1(n_503),
.B2(n_504),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_136),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_124),
.B(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_129),
.Y(n_444)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_130),
.Y(n_456)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_135),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_144),
.B2(n_146),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_142),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_143),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_146),
.Y(n_400)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_155),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_162),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_166),
.B(n_428),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_183),
.B1(n_184),
.B2(n_226),
.Y(n_167)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_169),
.B(n_170),
.C(n_183),
.Y(n_329)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_176),
.Y(n_408)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_213),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_197),
.B2(n_198),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_186),
.B(n_198),
.C(n_213),
.Y(n_333)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OR2x6_ASAP7_75t_SL g368 ( 
.A(n_188),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_188),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_188),
.A2(n_417),
.B1(n_418),
.B2(n_419),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_188),
.B(n_509),
.Y(n_508)
);

AO22x2_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_190),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_SL g196 ( 
.A(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_203),
.B(n_212),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_202),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_212),
.B(n_274),
.Y(n_450)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_220),
.Y(n_431)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_225),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_322),
.B(n_326),
.Y(n_227)
);

AOI21x1_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_278),
.B(n_321),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_264),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_230),
.B(n_264),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_252),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_231),
.A2(n_252),
.B1(n_253),
.B2(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_237),
.A3(n_241),
.B1(n_246),
.B2(n_249),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_257),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_257),
.B(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_265),
.B(n_276),
.C(n_277),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

OAI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_298),
.B(n_320),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_296),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_296),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_314),
.B(n_319),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_308),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_318),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_325),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_329),
.B(n_330),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_366),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_333),
.B(n_334),
.C(n_366),
.Y(n_478)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_348),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_336),
.B(n_348),
.Y(n_434)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_354),
.A2(n_370),
.B1(n_372),
.B2(n_374),
.Y(n_369)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_355),
.Y(n_512)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_393),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_367),
.B(n_394),
.C(n_401),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_376),
.B1(n_385),
.B2(n_392),
.Y(n_367)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_368),
.Y(n_418)
);

OAI22x1_ASAP7_75t_SL g461 ( 
.A1(n_368),
.A2(n_392),
.B1(n_420),
.B2(n_462),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_368),
.A2(n_462),
.B(n_508),
.Y(n_507)
);

INVx6_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_371),
.Y(n_375)
);

BUFx12f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_373),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_373),
.Y(n_423)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx5_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_384),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_395),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_477),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_446),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_413),
.B(n_446),
.C(n_484),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_435),
.C(n_436),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_414),
.B(n_480),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_434),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_424),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_424),
.C(n_434),
.Y(n_447)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B(n_427),
.Y(n_424)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_435),
.B(n_436),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_438),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_438),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_447),
.B(n_476),
.C(n_488),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_457),
.B1(n_458),
.B2(n_476),
.Y(n_448)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_451),
.Y(n_500)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_459),
.B(n_461),
.C(n_465),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_465),
.Y(n_460)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_478),
.B(n_479),
.Y(n_484)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g485 ( 
.A(n_486),
.B(n_516),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_489),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_489),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_490),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_499),
.Y(n_490)
);

OAI22xp33_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

XNOR2x1_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_507),
.Y(n_501)
);

INVx6_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);


endmodule