module fake_jpeg_17319_n_231 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_231);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_38),
.Y(n_43)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_1),
.Y(n_55)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_16),
.B1(n_26),
.B2(n_27),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_33),
.B1(n_42),
.B2(n_34),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_55),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_39),
.A2(n_16),
.B1(n_26),
.B2(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_1),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_25),
.B1(n_20),
.B2(n_15),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_60),
.B1(n_40),
.B2(n_44),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_29),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_28),
.B1(n_24),
.B2(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_33),
.B(n_41),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_80),
.B(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_70),
.C(n_71),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_29),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_3),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_62),
.B1(n_61),
.B2(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_18),
.B(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_44),
.Y(n_79)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_32),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_36),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_85),
.B(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_91),
.A2(n_98),
.B1(n_90),
.B2(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_48),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_93),
.B(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_70),
.B(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_97),
.B(n_107),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_73),
.B(n_4),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_69),
.B(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_103),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_3),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_84),
.Y(n_103)
);

OA21x2_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_73),
.B(n_78),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_78),
.B1(n_80),
.B2(n_73),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_106),
.B1(n_63),
.B2(n_50),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_62),
.B1(n_61),
.B2(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_78),
.B(n_34),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_125),
.B1(n_86),
.B2(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_118),
.B(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_87),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_113),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_80),
.B(n_73),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_115),
.B(n_97),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_120),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_75),
.C(n_67),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_42),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_75),
.B1(n_81),
.B2(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_126),
.B1(n_86),
.B2(n_89),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_34),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_36),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_50),
.B1(n_63),
.B2(n_83),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_57),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_104),
.A2(n_81),
.B1(n_66),
.B2(n_58),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_129),
.A2(n_93),
.B1(n_94),
.B2(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_107),
.B1(n_88),
.B2(n_101),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_135),
.B(n_145),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_95),
.B(n_88),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_147),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_150),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_72),
.B1(n_36),
.B2(n_35),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_146),
.B1(n_149),
.B2(n_68),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_72),
.B(n_5),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_19),
.B1(n_28),
.B2(n_22),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_54),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_122),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_127),
.B1(n_115),
.B2(n_118),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_31),
.B(n_21),
.C(n_19),
.D(n_30),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_123),
.C(n_119),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_154),
.C(n_164),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_117),
.C(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_142),
.B(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_167),
.Y(n_178)
);

BUFx12_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_160),
.Y(n_175)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_117),
.C(n_112),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_126),
.C(n_108),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_31),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_147),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_68),
.C(n_54),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_169),
.A2(n_144),
.B1(n_131),
.B2(n_145),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_171),
.A2(n_174),
.B1(n_168),
.B2(n_161),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_173),
.B(n_184),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_130),
.B1(n_133),
.B2(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_130),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_132),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_151),
.C(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_164),
.B(n_150),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_163),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_194),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_160),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_154),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_192),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_181),
.A2(n_161),
.B(n_169),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_189),
.A2(n_190),
.B(n_172),
.Y(n_201)
);

HAxp5_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_151),
.CON(n_190),
.SN(n_190)
);

AO21x1_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_174),
.B(n_171),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_173),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_196),
.B(n_170),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_SL g198 ( 
.A(n_190),
.B(n_193),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_198),
.A2(n_189),
.B(n_186),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_176),
.B(n_21),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_203),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_195),
.B(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_211),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_188),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_212),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_213),
.B(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_216),
.Y(n_220)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_201),
.B1(n_204),
.B2(n_206),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_218),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_3),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_21),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_6),
.A3(n_7),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_13),
.Y(n_226)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_218),
.A3(n_214),
.B1(n_215),
.B2(n_35),
.C1(n_51),
.C2(n_54),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_225),
.A3(n_226),
.B1(n_222),
.B2(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_227)
);

AOI322xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_228),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_224),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_6),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_14),
.Y(n_231)
);


endmodule