module fake_jpeg_21415_n_135 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_17),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_40),
.B(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_23),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_36),
.C(n_28),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_32),
.B1(n_14),
.B2(n_17),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_30),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_14),
.B1(n_26),
.B2(n_20),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_31),
.A2(n_34),
.B1(n_30),
.B2(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_26),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_53),
.B(n_55),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_63),
.B1(n_73),
.B2(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_40),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_36),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_68),
.C(n_46),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_16),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_69),
.Y(n_80)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_36),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_18),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_83),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_1),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_68),
.B(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_2),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

XOR2x2_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_102),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_62),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_78),
.C(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_63),
.B(n_59),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_103),
.B(n_82),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_59),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

A2O1A1O1Ixp25_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_89),
.B(n_87),
.C(n_91),
.D(n_90),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_112),
.B(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_111),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_76),
.C(n_83),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_54),
.B1(n_81),
.B2(n_88),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_93),
.B(n_98),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_115),
.A2(n_110),
.B(n_95),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_110),
.B1(n_104),
.B2(n_95),
.C(n_79),
.Y(n_124)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_114),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_122),
.A2(n_117),
.B(n_4),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_116),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_126),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_123),
.B1(n_122),
.B2(n_65),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_50),
.A3(n_5),
.B1(n_8),
.B2(n_10),
.C1(n_11),
.C2(n_13),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_128),
.B(n_3),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_130),
.B(n_5),
.Y(n_133)
);

OAI21x1_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_126),
.B(n_8),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_11),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_50),
.Y(n_135)
);


endmodule