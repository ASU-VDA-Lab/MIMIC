module fake_jpeg_6007_n_316 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_23),
.Y(n_68)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_22),
.Y(n_52)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_30),
.B(n_34),
.Y(n_79)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_58),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_18),
.B1(n_29),
.B2(n_24),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_31),
.B1(n_20),
.B2(n_34),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_31),
.B(n_29),
.C(n_27),
.Y(n_75)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_24),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_76),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_25),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_33),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_82),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_18),
.B1(n_34),
.B2(n_25),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_92),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_30),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_43),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_20),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_32),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_62),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_20),
.B1(n_30),
.B2(n_28),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_31),
.B1(n_26),
.B2(n_28),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_94),
.A2(n_59),
.B1(n_46),
.B2(n_63),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_62),
.B1(n_48),
.B2(n_51),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_115),
.B1(n_86),
.B2(n_71),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_101),
.B1(n_103),
.B2(n_107),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_92),
.B1(n_73),
.B2(n_75),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_56),
.B(n_58),
.C(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_119),
.Y(n_144)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_111),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_67),
.C(n_46),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_121),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_75),
.A2(n_59),
.B1(n_47),
.B2(n_54),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_78),
.Y(n_117)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_72),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_118),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_28),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_72),
.B(n_26),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_81),
.B(n_83),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_142),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_117),
.A2(n_84),
.B1(n_87),
.B2(n_93),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_99),
.B1(n_115),
.B2(n_116),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_130),
.A2(n_139),
.B(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_135),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_88),
.B(n_84),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_110),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_88),
.B1(n_80),
.B2(n_85),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_138),
.B1(n_145),
.B2(n_148),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_104),
.B1(n_115),
.B2(n_87),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_69),
.B(n_86),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_141),
.Y(n_160)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_152),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_146),
.B(n_96),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_106),
.A2(n_86),
.B1(n_94),
.B2(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx4_ASAP7_75t_SL g178 ( 
.A(n_149),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_80),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_65),
.A3(n_89),
.B1(n_67),
.B2(n_50),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_114),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_125),
.B1(n_124),
.B2(n_140),
.Y(n_197)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_105),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_139),
.B(n_125),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_156),
.B(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_163),
.B1(n_166),
.B2(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_112),
.C(n_116),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_162),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_112),
.C(n_120),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_100),
.B1(n_101),
.B2(n_103),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_121),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_168),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_103),
.B1(n_113),
.B2(n_119),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_71),
.B1(n_91),
.B2(n_83),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_113),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_174),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_172),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_152),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_175),
.A2(n_133),
.B(n_123),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_131),
.B(n_12),
.Y(n_176)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_129),
.A2(n_50),
.B1(n_67),
.B2(n_54),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_177),
.A2(n_149),
.B1(n_91),
.B2(n_32),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_128),
.B(n_50),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_27),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_135),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_169),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_206),
.C(n_208),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_179),
.B(n_21),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_197),
.B(n_179),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_160),
.B1(n_181),
.B2(n_174),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_0),
.Y(n_200)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_200),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_91),
.B1(n_32),
.B2(n_27),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_177),
.B1(n_163),
.B2(n_166),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_156),
.B(n_27),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_21),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_164),
.B(n_0),
.Y(n_210)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_186),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_229),
.Y(n_246)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_200),
.Y(n_216)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_155),
.B1(n_159),
.B2(n_167),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_235),
.B1(n_193),
.B2(n_203),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_204),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_226),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_153),
.B1(n_161),
.B2(n_162),
.Y(n_220)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_185),
.B1(n_195),
.B2(n_210),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_221),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_223),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_199),
.B(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_171),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_188),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_207),
.B(n_1),
.Y(n_242)
);

NOR4xp25_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_8),
.C(n_15),
.D(n_14),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_8),
.Y(n_253)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_7),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_190),
.A2(n_192),
.B1(n_194),
.B2(n_205),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_186),
.C(n_208),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_244),
.C(n_250),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_237),
.A2(n_235),
.B1(n_215),
.B2(n_228),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_246),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_242),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_220),
.B(n_7),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_231),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_7),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_249),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_0),
.C(n_1),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_8),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_216),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_13),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_266),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_213),
.B1(n_224),
.B2(n_222),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_234),
.B1(n_248),
.B2(n_3),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_262),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_267),
.C(n_236),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_235),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_247),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_237),
.B1(n_245),
.B2(n_240),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_223),
.B1(n_228),
.B2(n_211),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_4),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_255),
.C(n_239),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_275),
.C(n_279),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_259),
.A2(n_252),
.B(n_218),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_5),
.B(n_10),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_258),
.C(n_267),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_256),
.C(n_264),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_256),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_234),
.B(n_253),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_6),
.C(n_12),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_284),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g284 ( 
.A(n_260),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_286),
.A2(n_293),
.B(n_294),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_9),
.B1(n_12),
.B2(n_4),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_275),
.B1(n_16),
.B2(n_2),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_273),
.Y(n_288)
);

XOR2x2_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_295),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_290),
.C(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_6),
.C(n_11),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_5),
.C(n_11),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_277),
.B(n_16),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_295),
.A2(n_283),
.B(n_281),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_302),
.C(n_303),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_288),
.B(n_276),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_301),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_1),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_1),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_285),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_309),
.B(n_2),
.Y(n_311)
);

NOR2x1_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_292),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_2),
.CI(n_304),
.CON(n_312),
.SN(n_312)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_2),
.C(n_299),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_308),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_303),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_310),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_304),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_305),
.Y(n_316)
);


endmodule