module fake_jpeg_10718_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx9p33_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_13),
.B(n_8),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_32),
.Y(n_45)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_13),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_0),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_58),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_21),
.B1(n_23),
.B2(n_15),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_64),
.C(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_68),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_21),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_28),
.A2(n_22),
.B(n_14),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_64)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_33),
.B(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_34),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_73),
.B(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_37),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_9),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_65),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_48),
.B(n_10),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_66),
.C(n_48),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_50),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_92),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_64),
.B1(n_67),
.B2(n_61),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_101),
.B1(n_79),
.B2(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_30),
.B1(n_62),
.B2(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_100),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_62),
.B(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_31),
.B1(n_32),
.B2(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_106),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_84),
.B1(n_71),
.B2(n_70),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_SL g119 ( 
.A1(n_103),
.A2(n_94),
.A3(n_74),
.B1(n_95),
.B2(n_31),
.C1(n_32),
.C2(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_111),
.Y(n_113)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_98),
.B1(n_99),
.B2(n_84),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_100),
.B(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_92),
.C(n_87),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_110),
.C(n_108),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_112),
.B1(n_80),
.B2(n_81),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_125),
.B(n_116),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_111),
.C(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_115),
.A2(n_112),
.B1(n_105),
.B2(n_109),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_114),
.Y(n_130)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_126),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_129),
.B(n_130),
.Y(n_132)
);

AOI21x1_ASAP7_75t_L g131 ( 
.A1(n_128),
.A2(n_121),
.B(n_113),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_113),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_132),
.B(n_120),
.C(n_26),
.D(n_3),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_1),
.C(n_3),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_1),
.Y(n_136)
);


endmodule