module fake_jpeg_23555_n_324 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_15),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_22),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_30),
.A2(n_20),
.B1(n_29),
.B2(n_14),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_58),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_35),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_78),
.C(n_56),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_38),
.B1(n_29),
.B2(n_14),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_72),
.B1(n_30),
.B2(n_34),
.Y(n_92)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_20),
.B1(n_38),
.B2(n_32),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_76),
.B1(n_51),
.B2(n_48),
.Y(n_103)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_50),
.A2(n_14),
.B1(n_29),
.B2(n_20),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_70),
.A2(n_81),
.B1(n_24),
.B2(n_19),
.Y(n_99)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_45),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_22),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_20),
.B1(n_32),
.B2(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_31),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_29),
.B1(n_24),
.B2(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

NAND2xp67_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_15),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_84),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_89),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_88),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_84),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_93),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_97),
.B1(n_67),
.B2(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_94),
.A2(n_102),
.B1(n_108),
.B2(n_71),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_31),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_41),
.B1(n_42),
.B2(n_55),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_83),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g116 ( 
.A1(n_99),
.A2(n_15),
.B(n_28),
.Y(n_116)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_60),
.B1(n_55),
.B2(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_63),
.B1(n_71),
.B2(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_68),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_60),
.B1(n_48),
.B2(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_65),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_105),
.B(n_109),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_72),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_105),
.A2(n_61),
.B1(n_76),
.B2(n_64),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_112),
.B1(n_125),
.B2(n_85),
.Y(n_150)
);

OAI21xp33_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_116),
.B(n_117),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_132),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_109),
.A2(n_80),
.B1(n_77),
.B2(n_63),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_128),
.B1(n_133),
.B2(n_111),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_119),
.A2(n_91),
.B1(n_85),
.B2(n_100),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_80),
.C(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_123),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_75),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_129),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_86),
.A2(n_73),
.B1(n_79),
.B2(n_66),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_73),
.B1(n_67),
.B2(n_79),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_69),
.C(n_15),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_15),
.B1(n_28),
.B2(n_44),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_89),
.B1(n_102),
.B2(n_28),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_87),
.A2(n_24),
.B1(n_19),
.B2(n_15),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_15),
.B1(n_28),
.B2(n_102),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_94),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_138),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_137),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_141),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_152),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_103),
.C(n_107),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_33),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_154),
.B1(n_157),
.B2(n_159),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_160),
.B1(n_148),
.B2(n_153),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_131),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_156),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_122),
.B(n_91),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_94),
.B1(n_89),
.B2(n_93),
.Y(n_157)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_158),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_122),
.B(n_17),
.Y(n_161)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_141),
.A2(n_130),
.B1(n_118),
.B2(n_116),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_162),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_120),
.C(n_129),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_173),
.C(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_183),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_166),
.A2(n_36),
.B1(n_33),
.B2(n_59),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_110),
.B1(n_117),
.B2(n_112),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_175),
.B1(n_160),
.B2(n_36),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_117),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_182),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_142),
.C(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_127),
.B1(n_28),
.B2(n_126),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_127),
.B1(n_126),
.B2(n_28),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_28),
.B1(n_44),
.B2(n_59),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_59),
.B1(n_17),
.B2(n_96),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_96),
.C(n_40),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_16),
.B(n_21),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_180),
.A2(n_186),
.B(n_26),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_88),
.Y(n_197)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_96),
.A3(n_88),
.B1(n_40),
.B2(n_36),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_140),
.B1(n_147),
.B2(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_198),
.B1(n_190),
.B2(n_188),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_152),
.B(n_157),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_212),
.B(n_180),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_145),
.C(n_156),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_196),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_161),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_205),
.C(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_193),
.A2(n_195),
.B1(n_210),
.B2(n_213),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_166),
.A2(n_17),
.B1(n_16),
.B2(n_18),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_200),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_167),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_25),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_209),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_163),
.B(n_88),
.C(n_40),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_179),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_40),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_208),
.C(n_211),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_162),
.B(n_22),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_26),
.C(n_22),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_27),
.B(n_25),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_175),
.B1(n_176),
.B2(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

BUFx12_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_235),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_225),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_222),
.B(n_229),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_188),
.B1(n_174),
.B2(n_167),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_26),
.B1(n_7),
.B2(n_2),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_178),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_R g239 ( 
.A1(n_227),
.A2(n_193),
.B(n_195),
.Y(n_239)
);

NOR4xp25_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_21),
.C(n_18),
.D(n_27),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_201),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_198),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_7),
.B1(n_12),
.B2(n_2),
.Y(n_247)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_201),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_238),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_203),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_223),
.B1(n_220),
.B2(n_227),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_240),
.A2(n_231),
.B(n_215),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_216),
.B(n_212),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_203),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_219),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_207),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_251),
.C(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_247),
.A2(n_215),
.B1(n_218),
.B2(n_229),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_6),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_217),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_8),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_0),
.C(n_1),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_8),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_255),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_272),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_253),
.B1(n_237),
.B2(n_239),
.Y(n_257)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_246),
.B(n_222),
.CI(n_226),
.CON(n_258),
.SN(n_258)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_257),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_235),
.B1(n_230),
.B2(n_214),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_214),
.C(n_232),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_243),
.C(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_224),
.B1(n_234),
.B2(n_228),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_242),
.B1(n_254),
.B2(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_254),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_246),
.B(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_270),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_227),
.B1(n_233),
.B2(n_0),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_285),
.C(n_9),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_276),
.A2(n_279),
.B(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_278),
.B(n_10),
.Y(n_299)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_8),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_2),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_5),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_5),
.B(n_12),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_3),
.B(n_4),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_0),
.C(n_1),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_1),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_286),
.A2(n_272),
.B(n_270),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_262),
.B(n_263),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_288),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_290),
.B(n_293),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_258),
.B1(n_262),
.B2(n_267),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_291),
.A2(n_277),
.B1(n_275),
.B2(n_285),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_287),
.A2(n_258),
.B1(n_268),
.B2(n_4),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_279),
.A2(n_2),
.B(n_3),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_284),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_282),
.B1(n_286),
.B2(n_273),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_3),
.B(n_5),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_10),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_10),
.C(n_11),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_304),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_298),
.C(n_299),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_310),
.C(n_312),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_289),
.C(n_291),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_10),
.B(n_11),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_306),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_316),
.B(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_318),
.B(n_317),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_313),
.C(n_302),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_308),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_12),
.B(n_13),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_13),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_13),
.B(n_295),
.Y(n_324)
);


endmodule