module fake_jpeg_8297_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_17),
.B1(n_19),
.B2(n_24),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_47),
.A2(n_69),
.B1(n_16),
.B2(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_20),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_30),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_56),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_26),
.B1(n_29),
.B2(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_43),
.B1(n_36),
.B2(n_16),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_41),
.B(n_30),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_63)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_24),
.B1(n_17),
.B2(n_19),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_32),
.B1(n_31),
.B2(n_21),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_72),
.A2(n_78),
.B1(n_24),
.B2(n_19),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_32),
.B1(n_21),
.B2(n_43),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_21),
.B(n_18),
.C(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_18),
.Y(n_109)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_86),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_43),
.B1(n_36),
.B2(n_37),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_89),
.A2(n_59),
.B1(n_27),
.B2(n_37),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_43),
.B1(n_36),
.B2(n_16),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_90),
.A2(n_70),
.B1(n_83),
.B2(n_76),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_50),
.B1(n_64),
.B2(n_60),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_66),
.C(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_27),
.C(n_28),
.Y(n_111)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_100),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_69),
.B(n_47),
.C(n_58),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_114),
.B1(n_118),
.B2(n_84),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_89),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_67),
.B1(n_50),
.B2(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_107),
.B1(n_108),
.B2(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_104),
.B(n_106),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_84),
.B1(n_74),
.B2(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_54),
.B1(n_65),
.B2(n_44),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_44),
.B1(n_56),
.B2(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_23),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_61),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_37),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_113),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_44),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_33),
.B(n_27),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_73),
.B(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_42),
.Y(n_144)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_80),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_122),
.Y(n_129)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_133),
.Y(n_149)
);

NOR2x1p5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_59),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_146),
.B(n_115),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_139),
.B1(n_140),
.B2(n_98),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_145),
.B1(n_147),
.B2(n_96),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_135),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_82),
.B1(n_88),
.B2(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_102),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_101),
.Y(n_145)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_82),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_88),
.B1(n_18),
.B2(n_23),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_77),
.Y(n_148)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_114),
.C(n_107),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_151),
.C(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_111),
.C(n_113),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_161),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_113),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_159),
.B(n_33),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_116),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_163),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_140),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_108),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_167),
.C(n_42),
.Y(n_189)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_98),
.B(n_104),
.C(n_99),
.D(n_118),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_132),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_96),
.Y(n_166)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_122),
.C(n_68),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_169),
.B1(n_29),
.B2(n_28),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_123),
.A2(n_42),
.A3(n_29),
.B1(n_68),
.B2(n_61),
.Y(n_170)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_121),
.C(n_103),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_173),
.C(n_33),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_121),
.C(n_103),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_129),
.A2(n_42),
.B1(n_25),
.B2(n_28),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_148),
.B1(n_144),
.B2(n_25),
.Y(n_186)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_135),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_191),
.B(n_158),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_129),
.B1(n_125),
.B2(n_145),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_178),
.A2(n_195),
.B(n_197),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_139),
.B1(n_132),
.B2(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_187),
.B1(n_174),
.B2(n_149),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_180),
.B(n_165),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_33),
.B1(n_51),
.B2(n_45),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_172),
.A2(n_146),
.B1(n_124),
.B2(n_25),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_199),
.C(n_201),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_196),
.B1(n_193),
.B2(n_188),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_0),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_29),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_151),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_42),
.Y(n_193)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_167),
.A2(n_52),
.B1(n_51),
.B2(n_45),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_162),
.B(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_0),
.Y(n_198)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_33),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_2),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_171),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_189),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_192),
.C(n_199),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_201),
.C(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_213),
.Y(n_232)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_211),
.B(n_214),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_212),
.A2(n_221),
.B1(n_225),
.B2(n_194),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_181),
.B(n_158),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_215),
.B(n_222),
.Y(n_242)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_217),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_156),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_175),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_179),
.A2(n_170),
.B1(n_81),
.B2(n_52),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_11),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_223),
.B(n_224),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_195),
.A2(n_2),
.B(n_3),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_228),
.C(n_235),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_183),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_231),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_221),
.A2(n_212),
.B1(n_213),
.B2(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_204),
.C(n_207),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_241),
.C(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_180),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_239),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_200),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_203),
.B(n_176),
.Y(n_240)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_198),
.C(n_185),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_191),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_191),
.C(n_176),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_216),
.C(n_210),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_203),
.B(n_206),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_262),
.B(n_263),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_214),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_251),
.C(n_255),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_206),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_223),
.C(n_224),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_226),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_217),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_258),
.B(n_260),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_253),
.B(n_261),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_11),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_227),
.B1(n_230),
.B2(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_264),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_265),
.A2(n_268),
.B1(n_259),
.B2(n_250),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_270),
.C(n_273),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_227),
.B1(n_244),
.B2(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_3),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_228),
.C(n_81),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_81),
.C(n_45),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_15),
.B(n_14),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_276),
.B(n_12),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_14),
.B(n_13),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_248),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_281),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_13),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_3),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_265),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_288),
.C(n_276),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_267),
.Y(n_287)
);

AOI31xp33_ASAP7_75t_L g295 ( 
.A1(n_287),
.A2(n_275),
.A3(n_264),
.B(n_266),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_4),
.C(n_5),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_291),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_269),
.C(n_273),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_296),
.C(n_288),
.Y(n_300)
);

AOI31xp67_ASAP7_75t_L g303 ( 
.A1(n_295),
.A2(n_6),
.A3(n_7),
.B(n_8),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_4),
.C(n_6),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_286),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_299),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_291),
.C(n_293),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_297),
.A2(n_287),
.B(n_289),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_301),
.A2(n_303),
.B(n_304),
.Y(n_306)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_290),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_7),
.B(n_8),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_7),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g312 ( 
.A1(n_310),
.A2(n_306),
.B(n_8),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_9),
.C(n_311),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_9),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_9),
.Y(n_315)
);


endmodule