module fake_jpeg_13129_n_558 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_558);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_558;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_13),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_60),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_63),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g168 ( 
.A(n_64),
.Y(n_168)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_69),
.Y(n_164)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_72),
.Y(n_167)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_76),
.B(n_91),
.Y(n_141)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_53),
.Y(n_78)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_21),
.B(n_17),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_30),
.Y(n_82)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_83),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_17),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_87),
.B(n_90),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_32),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_17),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_59),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_16),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_98),
.Y(n_152)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_19),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_120),
.Y(n_155)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_32),
.Y(n_103)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx2_ASAP7_75t_R g104 ( 
.A(n_44),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_104),
.B(n_125),
.Y(n_195)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_106),
.Y(n_154)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_113),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_56),
.Y(n_114)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_115),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_33),
.Y(n_118)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_33),
.Y(n_119)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_50),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_46),
.Y(n_158)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_35),
.Y(n_122)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_122),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_35),
.Y(n_123)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_123),
.B(n_124),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_35),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_65),
.A2(n_58),
.B1(n_55),
.B2(n_38),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_126),
.A2(n_133),
.B1(n_113),
.B2(n_71),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_68),
.A2(n_35),
.B1(n_55),
.B2(n_34),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_129),
.A2(n_180),
.B(n_196),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_66),
.A2(n_54),
.B1(n_49),
.B2(n_46),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_146),
.B(n_165),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_64),
.A2(n_29),
.B(n_51),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_147),
.A2(n_176),
.B(n_186),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_81),
.B(n_49),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_162),
.B(n_163),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_45),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_72),
.B(n_45),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_70),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_174),
.B1(n_182),
.B2(n_187),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_89),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_64),
.A2(n_35),
.B1(n_52),
.B2(n_29),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_173),
.A2(n_179),
.B(n_186),
.C(n_197),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_105),
.A2(n_43),
.B1(n_42),
.B2(n_39),
.Y(n_174)
);

AO22x1_ASAP7_75t_SL g179 ( 
.A1(n_71),
.A2(n_52),
.B1(n_51),
.B2(n_47),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_74),
.B(n_20),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_198),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_93),
.A2(n_37),
.B1(n_41),
.B2(n_38),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_97),
.A2(n_41),
.B1(n_34),
.B2(n_27),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_109),
.A2(n_37),
.B1(n_47),
.B2(n_27),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_108),
.B(n_79),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_110),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_101),
.A2(n_26),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_16),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_114),
.A2(n_115),
.B1(n_77),
.B2(n_92),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_204),
.A2(n_83),
.B1(n_116),
.B2(n_118),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_16),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_78),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_206),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_141),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_211),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_156),
.B(n_106),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_208),
.B(n_240),
.Y(n_281)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_209),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx6_ASAP7_75t_L g299 ( 
.A(n_210),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_152),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_155),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_217),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_213),
.Y(n_314)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_214),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_215),
.Y(n_285)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_216),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_184),
.Y(n_218)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_218),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_127),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_219),
.B(n_221),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_222),
.B(n_238),
.Y(n_308)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_224),
.Y(n_317)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_225),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_122),
.B1(n_124),
.B2(n_119),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_226),
.A2(n_243),
.B1(n_271),
.B2(n_257),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_140),
.B(n_128),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_229),
.B(n_233),
.Y(n_279)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_164),
.Y(n_230)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_230),
.Y(n_323)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_231),
.Y(n_325)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_168),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_126),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_234),
.B(n_247),
.Y(n_298)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_149),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_241),
.A2(n_260),
.B1(n_263),
.B2(n_269),
.Y(n_296)
);

INVx3_ASAP7_75t_SL g244 ( 
.A(n_132),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_244),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_170),
.B(n_0),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_255),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_157),
.B(n_13),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_246),
.B(n_250),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_168),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_136),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_248),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_142),
.A2(n_12),
.B(n_5),
.C(n_6),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_262),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_144),
.B(n_12),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_153),
.B(n_0),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_251),
.B(n_254),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_139),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_252),
.A2(n_259),
.B(n_151),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_132),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_257),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_173),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_179),
.A2(n_5),
.B(n_8),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_256),
.B(n_272),
.Y(n_305)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_167),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_150),
.B(n_11),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_258),
.B(n_270),
.Y(n_303)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_167),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_144),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_261),
.B(n_271),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_178),
.B(n_201),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_175),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_139),
.A2(n_191),
.B1(n_134),
.B2(n_136),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_264),
.A2(n_228),
.B1(n_218),
.B2(n_210),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_197),
.A2(n_138),
.B1(n_134),
.B2(n_160),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_138),
.A2(n_130),
.B1(n_137),
.B2(n_135),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_159),
.A2(n_131),
.B1(n_192),
.B2(n_202),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_143),
.B(n_150),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_196),
.C(n_131),
.Y(n_284)
);

INVx8_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_202),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_180),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_189),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_273),
.B(n_245),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_177),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_274),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_242),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_276),
.B(n_295),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_220),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_286),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_318),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_208),
.B(n_177),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_290),
.B(n_216),
.Y(n_356)
);

NAND3xp33_ASAP7_75t_SL g340 ( 
.A(n_292),
.B(n_250),
.C(n_207),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_145),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_234),
.A2(n_145),
.B1(n_171),
.B2(n_265),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_306),
.A2(n_307),
.B1(n_326),
.B2(n_237),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_221),
.A2(n_171),
.B1(n_228),
.B2(n_243),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_311),
.A2(n_312),
.B1(n_316),
.B2(n_328),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_227),
.A2(n_264),
.B1(n_252),
.B2(n_236),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_227),
.A2(n_236),
.B1(n_238),
.B2(n_239),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_268),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_321),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_245),
.B(n_249),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_253),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_208),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_231),
.B(n_227),
.C(n_219),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_324),
.B(n_290),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_227),
.A2(n_245),
.B1(n_273),
.B2(n_230),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_325),
.Y(n_330)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

NOR2x1_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_287),
.Y(n_334)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_334),
.Y(n_372)
);

OA22x2_ASAP7_75t_L g395 ( 
.A1(n_335),
.A2(n_322),
.B1(n_283),
.B2(n_278),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_324),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_355),
.Y(n_384)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_337),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_327),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_339),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_302),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_340),
.A2(n_364),
.B(n_285),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_284),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_275),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_361),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_311),
.A2(n_232),
.B1(n_224),
.B2(n_223),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_344),
.A2(n_348),
.B1(n_352),
.B2(n_309),
.Y(n_390)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_277),
.B(n_211),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g401 ( 
.A(n_346),
.B(n_291),
.C(n_313),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_312),
.A2(n_263),
.B1(n_241),
.B2(n_209),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_326),
.A2(n_213),
.B1(n_225),
.B2(n_269),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_349),
.A2(n_351),
.B1(n_357),
.B2(n_358),
.Y(n_387)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_280),
.Y(n_350)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_350),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_292),
.A2(n_260),
.B1(n_214),
.B2(n_272),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_328),
.A2(n_240),
.B1(n_255),
.B2(n_235),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_212),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_353),
.B(n_304),
.Y(n_396)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_244),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_356),
.B(n_362),
.C(n_313),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_288),
.A2(n_261),
.B1(n_300),
.B2(n_306),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_288),
.A2(n_321),
.B1(n_298),
.B2(n_295),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_360),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_289),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_281),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_286),
.A2(n_319),
.B1(n_320),
.B2(n_297),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_366),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_310),
.A2(n_305),
.B1(n_308),
.B2(n_289),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_310),
.A2(n_318),
.B1(n_309),
.B2(n_314),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_289),
.B(n_303),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_294),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_368),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_301),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_323),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_347),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_379),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_335),
.A2(n_282),
.B1(n_305),
.B2(n_296),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_377),
.A2(n_381),
.B1(n_386),
.B2(n_357),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_378),
.B(n_356),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_281),
.Y(n_380)
);

XNOR2x1_ASAP7_75t_SL g429 ( 
.A(n_380),
.B(n_402),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_360),
.A2(n_293),
.B1(n_281),
.B2(n_279),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_348),
.A2(n_299),
.B1(n_314),
.B2(n_323),
.Y(n_386)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_390),
.Y(n_405)
);

NAND2x1_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_322),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_392),
.A2(n_361),
.B(n_329),
.Y(n_428)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_393),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_394),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_344),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_401),
.Y(n_412)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_350),
.Y(n_399)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_399),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_336),
.C(n_397),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_283),
.Y(n_402)
);

OAI22x1_ASAP7_75t_L g450 ( 
.A1(n_407),
.A2(n_395),
.B1(n_378),
.B2(n_386),
.Y(n_450)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_370),
.Y(n_410)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_411),
.B(n_418),
.C(n_381),
.Y(n_444)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_413),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_339),
.Y(n_414)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_414),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_387),
.A2(n_388),
.B1(n_379),
.B2(n_385),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_362),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_416),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_367),
.Y(n_418)
);

NOR2xp67_ASAP7_75t_R g419 ( 
.A(n_388),
.B(n_355),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_358),
.Y(n_421)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_421),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_377),
.A2(n_341),
.B1(n_349),
.B2(n_342),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_422),
.A2(n_425),
.B1(n_432),
.B2(n_433),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_376),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_423),
.B(n_431),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_424),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_380),
.A2(n_341),
.B1(n_363),
.B2(n_329),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_343),
.Y(n_426)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_426),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_369),
.Y(n_427)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_428),
.A2(n_430),
.B(n_403),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_403),
.A2(n_341),
.B(n_364),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_371),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_387),
.A2(n_333),
.B1(n_366),
.B2(n_367),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_385),
.A2(n_330),
.B1(n_337),
.B2(n_334),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_411),
.B(n_400),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_436),
.B(n_439),
.Y(n_478)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_420),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_440),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_432),
.B(n_384),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_414),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_427),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_442),
.B(n_455),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_446),
.C(n_449),
.Y(n_465)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_405),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_416),
.C(n_425),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_380),
.C(n_392),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_450),
.A2(n_422),
.B1(n_405),
.B2(n_421),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_426),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_456),
.A2(n_428),
.B(n_406),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_395),
.C(n_391),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_449),
.C(n_446),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_407),
.A2(n_395),
.B1(n_399),
.B2(n_398),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_459),
.A2(n_433),
.B1(n_417),
.B2(n_408),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_416),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_466),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_453),
.B(n_412),
.C(n_424),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_462),
.B(n_477),
.Y(n_493)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_463),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_435),
.A2(n_404),
.B1(n_417),
.B2(n_430),
.Y(n_464)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_464),
.Y(n_490)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_467),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_468),
.A2(n_402),
.B(n_372),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_469),
.A2(n_480),
.B1(n_448),
.B2(n_457),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_429),
.C(n_404),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_472),
.C(n_479),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_429),
.C(n_415),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_439),
.B(n_429),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_483),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_412),
.B1(n_413),
.B2(n_409),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_447),
.A2(n_441),
.B1(n_448),
.B2(n_451),
.Y(n_475)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_475),
.Y(n_502)
);

BUFx12f_ASAP7_75t_SL g476 ( 
.A(n_458),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g486 ( 
.A1(n_476),
.A2(n_456),
.B(n_457),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g477 ( 
.A(n_454),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_443),
.B(n_410),
.C(n_409),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_447),
.A2(n_419),
.B1(n_402),
.B2(n_373),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_372),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_484),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_486),
.A2(n_472),
.B(n_479),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_469),
.A2(n_445),
.B1(n_438),
.B2(n_450),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_471),
.B(n_459),
.CI(n_460),
.CON(n_491),
.SN(n_491)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_491),
.B(n_501),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_481),
.B(n_434),
.Y(n_492)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_492),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_437),
.C(n_373),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_497),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_470),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_464),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_480),
.A2(n_398),
.B1(n_389),
.B2(n_331),
.Y(n_499)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_499),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_475),
.B(n_389),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_478),
.C(n_465),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_503),
.B(n_506),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_513),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_465),
.C(n_466),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_493),
.B(n_476),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_507),
.B(n_517),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_496),
.A2(n_487),
.B1(n_492),
.B2(n_502),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_508),
.A2(n_496),
.B1(n_489),
.B2(n_484),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_461),
.C(n_483),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_495),
.C(n_500),
.Y(n_521)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_488),
.B(n_354),
.C(n_473),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_512),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_495),
.B(n_393),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_515),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_518),
.B(n_519),
.Y(n_530)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_514),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_522),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_500),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_487),
.C(n_490),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_524),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_504),
.B(n_486),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_525),
.B(n_526),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_490),
.C(n_502),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_511),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_533),
.B(n_534),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_491),
.Y(n_534)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_529),
.A2(n_509),
.B(n_516),
.Y(n_535)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_535),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_526),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_482),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_521),
.B(n_509),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_537),
.A2(n_522),
.B(n_520),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g538 ( 
.A(n_525),
.B(n_498),
.C(n_501),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_538),
.A2(n_505),
.B(n_491),
.Y(n_542)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_540),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_520),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_541),
.A2(n_544),
.B(n_383),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_542),
.A2(n_546),
.B(n_291),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_532),
.A2(n_513),
.B(n_420),
.Y(n_544)
);

AO221x1_ASAP7_75t_L g547 ( 
.A1(n_543),
.A2(n_539),
.B1(n_535),
.B2(n_530),
.C(n_538),
.Y(n_547)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_547),
.B(n_299),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_499),
.C(n_383),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_548),
.A2(n_550),
.B(n_317),
.Y(n_553)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_541),
.B(n_278),
.Y(n_552)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_552),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_555),
.A2(n_549),
.B(n_554),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_553),
.C(n_317),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_315),
.Y(n_558)
);


endmodule