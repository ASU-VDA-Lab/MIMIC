module real_jpeg_29221_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_299, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_299;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_293;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_242;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_285;
wire n_45;
wire n_160;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_295;
wire n_167;
wire n_179;
wire n_133;
wire n_202;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_0),
.B(n_29),
.Y(n_28)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_1),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g147 ( 
.A1(n_1),
.A2(n_47),
.B(n_51),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_1),
.B(n_49),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_1),
.A2(n_63),
.B(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_1),
.B(n_63),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_1),
.B(n_104),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_1),
.A2(n_27),
.B1(n_35),
.B2(n_225),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_1),
.A2(n_50),
.B(n_241),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_2),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_91)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_4),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_4),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_107),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_107),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_107),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_8),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_66),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_50),
.B1(n_51),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_9),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_88),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_88),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_88),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_10),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_144),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_144),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_144),
.Y(n_225)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_11),
.A2(n_30),
.A3(n_63),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_12),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_133),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_133),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_133),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_13),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_13),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_42),
.Y(n_214)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_16),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_16),
.A2(n_50),
.B1(n_51),
.B2(n_75),
.Y(n_116)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_108),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_22),
.B(n_108),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_78),
.C(n_93),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_23),
.B(n_78),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_23)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_25),
.A2(n_39),
.B(n_57),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_25),
.A2(n_26),
.B1(n_59),
.B2(n_60),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_33),
.B(n_36),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_27),
.A2(n_36),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_27),
.A2(n_97),
.B1(n_98),
.B2(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_27),
.A2(n_33),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_27),
.A2(n_33),
.B1(n_219),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_27),
.A2(n_98),
.B1(n_214),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_28),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_34),
.B1(n_149),
.B2(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_28),
.A2(n_34),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_29),
.A2(n_30),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_29),
.B(n_71),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_29),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_45),
.B1(n_54),
.B2(n_56),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_46),
.B1(n_49),
.B2(n_106),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_43),
.A2(n_53),
.B(n_142),
.C(n_147),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

O2A1O1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_45),
.A2(n_54),
.B1(n_56),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_45),
.A2(n_56),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_46),
.A2(n_49),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_46),
.A2(n_49),
.B1(n_106),
.B2(n_173),
.Y(n_187)
);

AO22x1_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_49)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_81),
.B(n_83),
.C(n_84),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_81),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_50),
.A2(n_64),
.A3(n_81),
.B1(n_242),
.B2(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_51),
.B(n_142),
.Y(n_242)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_67),
.B1(n_73),
.B2(n_76),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_68),
.B1(n_69),
.B2(n_100),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_63),
.B(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_67),
.A2(n_76),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_67),
.A2(n_76),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_68),
.A2(n_69),
.B1(n_74),
.B2(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_68),
.A2(n_69),
.B(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_68),
.A2(n_69),
.B1(n_100),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_68),
.A2(n_69),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_68),
.A2(n_69),
.B1(n_200),
.B2(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_68),
.A2(n_69),
.B1(n_138),
.B2(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_69),
.B(n_142),
.Y(n_226)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_90),
.B(n_92),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_90),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_86),
.B2(n_89),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_80),
.A2(n_84),
.B1(n_131),
.B2(n_134),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_80),
.A2(n_84),
.B1(n_134),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_80),
.A2(n_84),
.B1(n_156),
.B2(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_81),
.Y(n_251)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_109),
.CI(n_121),
.CON(n_108),
.SN(n_108)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_93),
.A2(n_94),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.C(n_105),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_95),
.B(n_101),
.CI(n_105),
.CON(n_279),
.SN(n_279)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_96),
.B(n_99),
.Y(n_183)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_176),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_103),
.A2(n_104),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_104),
.B1(n_132),
.B2(n_155),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g296 ( 
.A(n_108),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_113),
.B2(n_120),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_114),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_117),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_277),
.A3(n_285),
.B1(n_290),
.B2(n_295),
.C(n_299),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_178),
.C(n_190),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_160),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_126),
.B(n_160),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_145),
.C(n_152),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_127),
.B(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_140),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_135),
.B2(n_136),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_136),
.C(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_142),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_145),
.A2(n_152),
.B1(n_153),
.B2(n_275),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_145),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_148),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_151),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_154),
.B(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_157),
.B(n_159),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_158),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_167),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_167),
.C(n_168),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_165),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_177),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_174),
.C(n_177),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g291 ( 
.A1(n_179),
.A2(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_180),
.B(n_181),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_189),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_183),
.B(n_184),
.C(n_189),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_185),
.B(n_187),
.C(n_188),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_271),
.B(n_276),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_257),
.B(n_270),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_235),
.B(n_256),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_215),
.B(n_234),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_195),
.B(n_205),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_199),
.Y(n_203)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_212),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_210),
.C(n_212),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_213),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_222),
.B(n_233),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_227),
.B(n_232),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_226),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_237),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_248),
.B1(n_254),
.B2(n_255),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_243),
.B1(n_246),
.B2(n_247),
.Y(n_238)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_243),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_247),
.C(n_255),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_248),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_252),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_258),
.B(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_264),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_266),
.C(n_268),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_266),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_272),
.B(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_282),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_282),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.C(n_281),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_279),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_286),
.A2(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_287),
.B(n_288),
.Y(n_294)
);


endmodule