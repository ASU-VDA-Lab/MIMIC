module real_jpeg_32025_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_715;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_669;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_719;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_578;
wire n_149;
wire n_620;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_704;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_673;
wire n_175;
wire n_338;
wire n_653;
wire n_718;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_703;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_697;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_716;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_670;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_712;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_714;
wire n_89;
wire n_407;
wire n_693;
wire n_721;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_711;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_635;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_720;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_708;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_457;
wire n_717;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_602;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_636;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_722;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_713;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_0),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_0),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_0),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_1),
.A2(n_69),
.B1(n_176),
.B2(n_179),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_1),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_1),
.A2(n_179),
.B1(n_399),
.B2(n_400),
.Y(n_398)
);

OAI22x1_ASAP7_75t_SL g487 ( 
.A1(n_1),
.A2(n_179),
.B1(n_488),
.B2(n_495),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_1),
.A2(n_179),
.B1(n_578),
.B2(n_580),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_2),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_4),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_4),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_4),
.B(n_26),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g601 ( 
.A1(n_4),
.A2(n_505),
.B1(n_602),
.B2(n_604),
.Y(n_601)
);

OAI21xp33_ASAP7_75t_L g675 ( 
.A1(n_4),
.A2(n_278),
.B(n_626),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_5),
.A2(n_166),
.B1(n_167),
.B2(n_171),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_5),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_5),
.A2(n_166),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_5),
.A2(n_166),
.B1(n_387),
.B2(n_389),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_5),
.A2(n_166),
.B1(n_520),
.B2(n_524),
.Y(n_519)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_6),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_7),
.A2(n_63),
.B1(n_394),
.B2(n_395),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_7),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_7),
.A2(n_394),
.B1(n_480),
.B2(n_484),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_7),
.A2(n_394),
.B1(n_593),
.B2(n_597),
.Y(n_592)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_7),
.A2(n_394),
.B1(n_635),
.B2(n_636),
.Y(n_634)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_8),
.A2(n_67),
.B1(n_68),
.B2(n_72),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_67),
.B1(n_152),
.B2(n_156),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_8),
.A2(n_67),
.B1(n_224),
.B2(n_227),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_8),
.A2(n_67),
.B1(n_273),
.B2(n_276),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_9),
.A2(n_68),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_9),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_9),
.A2(n_184),
.B1(n_249),
.B2(n_253),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_9),
.A2(n_184),
.B1(n_263),
.B2(n_267),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_9),
.A2(n_184),
.B1(n_383),
.B2(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_10),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_10),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_10),
.A2(n_287),
.B1(n_451),
.B2(n_454),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_10),
.A2(n_152),
.B1(n_287),
.B2(n_555),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_10),
.A2(n_287),
.B1(n_621),
.B2(n_624),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_11),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_12),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_13),
.Y(n_99)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_13),
.Y(n_648)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_14),
.Y(n_131)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_14),
.Y(n_135)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_14),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_20),
.B(n_721),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_15),
.B(n_722),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_16),
.A2(n_57),
.B1(n_58),
.B2(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_16),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_16),
.A2(n_57),
.B1(n_101),
.B2(n_105),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_16),
.A2(n_57),
.B1(n_234),
.B2(n_237),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_16),
.A2(n_57),
.B1(n_327),
.B2(n_331),
.Y(n_326)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_17),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_17),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_17),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_18),
.A2(n_112),
.B1(n_118),
.B2(n_119),
.Y(n_111)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_18),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_18),
.A2(n_118),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_18),
.A2(n_118),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_18),
.A2(n_118),
.B1(n_379),
.B2(n_383),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_76),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_65),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_39),
.B(n_56),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_25),
.A2(n_39),
.B1(n_56),
.B2(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_25),
.A2(n_39),
.B1(n_165),
.B2(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_25),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_25),
.A2(n_39),
.B1(n_66),
.B2(n_342),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_26),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_26),
.B(n_175),
.Y(n_283)
);

AO22x1_ASAP7_75t_L g392 ( 
.A1(n_26),
.A2(n_42),
.B1(n_285),
.B2(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_26),
.B(n_393),
.Y(n_413)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_30),
.Y(n_435)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_30),
.Y(n_444)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_32),
.Y(n_606)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_33),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_33),
.Y(n_440)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_36),
.Y(n_211)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_36),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_40),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_316)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_41),
.B(n_501),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_42),
.B(n_175),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_42),
.B(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_51),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_51),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_51),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_51),
.Y(n_290)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_61),
.Y(n_322)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_65),
.B(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_65),
.B(n_338),
.Y(n_720)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_75),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_352),
.B(n_711),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_336),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_309),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_256),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g713 ( 
.A(n_82),
.B(n_256),
.Y(n_713)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_180),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_84),
.B(n_334),
.C(n_335),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_161),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XOR2x2_ASAP7_75t_L g301 ( 
.A(n_86),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_110),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_87),
.B(n_163),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_87),
.A2(n_369),
.B1(n_370),
.B2(n_371),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_87),
.Y(n_369)
);

OA21x2_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_94),
.B(n_100),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_91),
.Y(n_376)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_93),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_94),
.Y(n_278)
);

AO22x1_ASAP7_75t_L g416 ( 
.A1(n_94),
.A2(n_378),
.B1(n_417),
.B2(n_421),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_94),
.B(n_577),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_94),
.A2(n_633),
.B1(n_637),
.B2(n_640),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_95),
.Y(n_280)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx8_ASAP7_75t_L g575 ( 
.A(n_96),
.Y(n_575)
);

INVx8_ASAP7_75t_L g628 ( 
.A(n_96),
.Y(n_628)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_97),
.Y(n_623)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_99),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_99),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_99),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_100),
.B(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_102),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_104),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_104),
.Y(n_526)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_104),
.Y(n_583)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_105),
.Y(n_678)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_108),
.Y(n_523)
);

INVx4_ASAP7_75t_L g579 ( 
.A(n_108),
.Y(n_579)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_109),
.Y(n_625)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_110),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_124),
.B1(n_149),
.B2(n_151),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_111),
.A2(n_124),
.B1(n_149),
.B2(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_115),
.Y(n_155)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_115),
.Y(n_568)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_116),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_117),
.Y(n_236)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_123),
.Y(n_558)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_124),
.A2(n_149),
.B1(n_262),
.B2(n_386),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_SL g553 ( 
.A1(n_124),
.A2(n_554),
.B(n_559),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_124),
.A2(n_149),
.B1(n_554),
.B2(n_592),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_136),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_128),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_135),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_140),
.B1(n_143),
.B2(n_145),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_139),
.Y(n_661)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_142),
.Y(n_599)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_142),
.Y(n_672)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g680 ( 
.A(n_149),
.B(n_505),
.Y(n_680)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_150),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_150),
.B(n_233),
.Y(n_244)
);

AOI22x1_ASAP7_75t_L g486 ( 
.A1(n_150),
.A2(n_232),
.B1(n_487),
.B2(n_498),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_150),
.B(n_487),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_150),
.B(n_615),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_151),
.Y(n_246)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_154),
.Y(n_651)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_160),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_174),
.Y(n_163)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_168),
.Y(n_286)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx4f_ASAP7_75t_SL g186 ( 
.A(n_173),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_174),
.B(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_178),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_241),
.B1(n_254),
.B2(n_255),
.Y(n_180)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_181),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_181),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_182),
.B(n_240),
.C(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_183),
.Y(n_317)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_230),
.B1(n_231),
.B2(n_240),
.Y(n_187)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_212),
.B1(n_220),
.B2(n_223),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_189),
.A2(n_212),
.B1(n_220),
.B2(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_189),
.A2(n_222),
.B1(n_248),
.B2(n_294),
.Y(n_293)
);

AO22x1_ASAP7_75t_L g325 ( 
.A1(n_189),
.A2(n_220),
.B1(n_223),
.B2(n_326),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_R g344 ( 
.A1(n_189),
.A2(n_220),
.B(n_326),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g403 ( 
.A(n_189),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_189),
.B(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_189),
.B(n_398),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_200),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_190),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_195),
.B2(n_197),
.Y(n_190)
);

INVx5_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_194),
.Y(n_573)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_203),
.B1(n_206),
.B2(n_210),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_204),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_205),
.Y(n_402)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_215),
.Y(n_442)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

AOI21x1_ASAP7_75t_L g476 ( 
.A1(n_220),
.A2(n_477),
.B(n_478),
.Y(n_476)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI22x1_ASAP7_75t_L g396 ( 
.A1(n_221),
.A2(n_397),
.B1(n_403),
.B2(n_404),
.Y(n_396)
);

OAI21xp33_ASAP7_75t_SL g515 ( 
.A1(n_221),
.A2(n_516),
.B(n_517),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_221),
.B(n_505),
.Y(n_617)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_222),
.B(n_398),
.Y(n_458)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_229),
.Y(n_332)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_229),
.Y(n_453)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_229),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_230),
.B(n_316),
.C(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_231),
.Y(n_312)
);

XOR2x1_ASAP7_75t_L g324 ( 
.A(n_231),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_232),
.B(n_487),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_232),
.B(n_669),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_236),
.Y(n_239)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_241),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVxp67_ASAP7_75t_SL g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_243),
.B(n_305),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_245),
.C(n_247),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_244),
.Y(n_306)
);

INVxp33_ASAP7_75t_L g307 ( 
.A(n_245),
.Y(n_307)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_247),
.Y(n_308)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_249),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_251),
.Y(n_483)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_251),
.Y(n_603)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_299),
.C(n_303),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g358 ( 
.A(n_258),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_281),
.C(n_291),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_260),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_271),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_261),
.B(n_271),
.Y(n_410)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_265),
.Y(n_388)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_278),
.B(n_279),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_272),
.A2(n_278),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_273),
.Y(n_635)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22x1_ASAP7_75t_L g518 ( 
.A1(n_278),
.A2(n_422),
.B1(n_519),
.B2(n_527),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_278),
.A2(n_620),
.B(n_626),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_282),
.A2(n_292),
.B1(n_293),
.B2(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_283),
.B(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_294),
.Y(n_404)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx5_ASAP7_75t_L g399 ( 
.A(n_298),
.Y(n_399)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_301),
.B(n_360),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B(n_308),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_309),
.A2(n_346),
.B(n_713),
.C(n_714),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_333),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_310),
.B(n_333),
.Y(n_714)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g351 ( 
.A(n_311),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_314),
.B(n_350),
.C(n_351),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

XNOR2x1_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_324),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_319),
.Y(n_342)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx3_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_322),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g711 ( 
.A1(n_337),
.A2(n_712),
.B(n_715),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_337),
.Y(n_718)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.C(n_343),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_339),
.B(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_341),
.B(n_343),
.Y(n_348)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_347),
.B(n_349),
.Y(n_717)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2x1_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_539),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_463),
.B(n_535),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_356),
.B(n_708),
.Y(n_707)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_361),
.B(n_405),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_357),
.B(n_361),
.Y(n_538)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_358),
.B(n_362),
.Y(n_536)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.C(n_372),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_364),
.B(n_460),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_368),
.A2(n_373),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_392),
.C(n_396),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_385),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_375),
.B(n_385),
.Y(n_472)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_386),
.Y(n_498)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_403),
.A2(n_450),
.B(n_458),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_403),
.A2(n_458),
.B(n_601),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_459),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_406),
.B(n_459),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_410),
.C(n_411),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_408),
.B(n_410),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.C(n_448),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_414),
.C(n_448),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_449),
.Y(n_471)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_415),
.B(n_471),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_425),
.Y(n_415)
);

XNOR2x2_ASAP7_75t_SL g512 ( 
.A(n_416),
.B(n_426),
.Y(n_512)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_420),
.Y(n_685)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_426),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_436),
.B1(n_441),
.B2(n_445),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_433),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx4_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_432),
.Y(n_504)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx2_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVxp33_ASAP7_75t_L g506 ( 
.A(n_445),
.Y(n_506)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_451),
.A2(n_562),
.B1(n_565),
.B2(n_569),
.Y(n_561)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_452),
.B(n_570),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_468),
.C(n_507),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g708 ( 
.A1(n_465),
.A2(n_709),
.B(n_710),
.Y(n_708)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_468),
.Y(n_709)
);

MAJx2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.C(n_473),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_470),
.B(n_534),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_472),
.B(n_474),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_485),
.C(n_499),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_486),
.Y(n_511)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx3_ASAP7_75t_SL g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_494),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_494),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_494),
.Y(n_596)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_499),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_502),
.A2(n_505),
.B(n_506),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_505),
.B(n_563),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_505),
.B(n_566),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_505),
.B(n_663),
.Y(n_662)
);

OAI21xp33_ASAP7_75t_SL g669 ( 
.A1(n_505),
.A2(n_662),
.B(n_670),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_505),
.B(n_628),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_533),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_508),
.B(n_533),
.Y(n_710)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_512),
.C(n_513),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_509),
.B(n_544),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g547 ( 
.A(n_509),
.B(n_544),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_511),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_512),
.A2(n_513),
.B1(n_514),
.B2(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_512),
.Y(n_545)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_518),
.C(n_531),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g550 ( 
.A(n_515),
.B(n_551),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_532),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g574 ( 
.A1(n_519),
.A2(n_575),
.B(n_576),
.Y(n_574)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_524),
.Y(n_636)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_536),
.A2(n_537),
.B(n_538),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_707),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_541),
.A2(n_584),
.B(n_705),
.Y(n_540)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_542),
.A2(n_546),
.B(n_548),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_543),
.B(n_547),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_548),
.B(n_706),
.Y(n_705)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_552),
.C(n_560),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_549),
.A2(n_550),
.B1(n_700),
.B2(n_701),
.Y(n_699)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_552),
.A2(n_553),
.B1(n_560),
.B2(n_702),
.Y(n_701)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_558),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_559),
.B(n_668),
.Y(n_667)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_560),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_574),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_561),
.B(n_574),
.Y(n_589)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

OAI21xp33_ASAP7_75t_L g681 ( 
.A1(n_576),
.A2(n_634),
.B(n_682),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_577),
.B(n_627),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

AOI21x1_ASAP7_75t_L g584 ( 
.A1(n_585),
.A2(n_696),
.B(n_703),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_586),
.A2(n_629),
.B(n_694),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_607),
.B(n_609),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_588),
.B(n_608),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_590),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_589),
.B(n_590),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g697 ( 
.A(n_589),
.B(n_591),
.C(n_600),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_SL g590 ( 
.A(n_591),
.B(n_600),
.Y(n_590)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_592),
.Y(n_615)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx3_ASAP7_75t_SL g598 ( 
.A(n_599),
.Y(n_598)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_603),
.Y(n_602)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_609),
.B(n_695),
.Y(n_694)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_610),
.B(n_616),
.C(n_618),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g692 ( 
.A(n_612),
.B(n_617),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_613),
.B(n_614),
.Y(n_612)
);

INVxp33_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_618),
.A2(n_619),
.B1(n_691),
.B2(n_692),
.Y(n_690)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_620),
.Y(n_640)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

AOI21x1_ASAP7_75t_L g629 ( 
.A1(n_630),
.A2(n_688),
.B(n_693),
.Y(n_629)
);

AO21x1_ASAP7_75t_SL g630 ( 
.A1(n_631),
.A2(n_673),
.B(n_687),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_641),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g687 ( 
.A(n_632),
.B(n_641),
.Y(n_687)
);

INVxp33_ASAP7_75t_SL g633 ( 
.A(n_634),
.Y(n_633)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_639),
.Y(n_638)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_642),
.B(n_667),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g689 ( 
.A(n_642),
.B(n_667),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_SL g642 ( 
.A1(n_643),
.A2(n_649),
.B(n_657),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_644),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_645),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_648),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_652),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

AOI21xp33_ASAP7_75t_L g657 ( 
.A1(n_658),
.A2(n_660),
.B(n_662),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_661),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_665),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

BUFx4f_ASAP7_75t_SL g670 ( 
.A(n_671),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_672),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_674),
.A2(n_679),
.B(n_686),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_675),
.B(n_676),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g676 ( 
.A(n_677),
.B(n_678),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_680),
.B(n_681),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_680),
.B(n_681),
.Y(n_686)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_683),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_684),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_685),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_689),
.B(n_690),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_689),
.B(n_690),
.Y(n_693)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_692),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_697),
.B(n_698),
.Y(n_696)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_697),
.Y(n_704)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_699),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g703 ( 
.A(n_699),
.B(n_704),
.Y(n_703)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_701),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_716),
.A2(n_718),
.B(n_719),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_717),
.Y(n_716)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_720),
.Y(n_719)
);


endmodule