module fake_netlist_1_7992_n_719 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_719);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_719;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp67_ASAP7_75t_SL g80 ( .A(n_12), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_29), .Y(n_81) );
BUFx3_ASAP7_75t_L g82 ( .A(n_79), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_40), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_52), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_38), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_51), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_43), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_68), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_50), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_0), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_35), .Y(n_92) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_72), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_30), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx2_ASAP7_75t_SL g96 ( .A(n_6), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_25), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_12), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_61), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_18), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_53), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_47), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_4), .Y(n_103) );
BUFx10_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
INVx1_ASAP7_75t_SL g105 ( .A(n_24), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_64), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_28), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_5), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_49), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_21), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_76), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_46), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_58), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_14), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_54), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_66), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_67), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_5), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_48), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
BUFx10_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_37), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_45), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_57), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_108), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_103), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_93), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_103), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_93), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_93), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_92), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_106), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_92), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_95), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_106), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_95), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_118), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_118), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_85), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_96), .B(n_3), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_87), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_104), .B(n_7), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_82), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_104), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_104), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_85), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_89), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_97), .Y(n_160) );
INVxp33_ASAP7_75t_SL g161 ( .A(n_88), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_125), .B(n_96), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_117), .Y(n_163) );
AND2x4_ASAP7_75t_L g164 ( .A(n_124), .B(n_8), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_99), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_88), .B(n_78), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_124), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_100), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_101), .Y(n_169) );
NOR2x1_ASAP7_75t_L g170 ( .A(n_102), .B(n_8), .Y(n_170) );
HB1xp67_ASAP7_75t_L g171 ( .A(n_98), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_90), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_138), .B(n_143), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_164), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_138), .B(n_115), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_138), .B(n_115), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_138), .B(n_125), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_135), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
OAI22xp5_ASAP7_75t_L g184 ( .A1(n_143), .A2(n_122), .B1(n_113), .B2(n_91), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_161), .B(n_162), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_135), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_162), .B(n_112), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_163), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_172), .B(n_128), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_135), .Y(n_191) );
INVx3_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
BUFx3_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
INVx5_ASAP7_75t_L g194 ( .A(n_164), .Y(n_194) );
INVx1_ASAP7_75t_SL g195 ( .A(n_139), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_171), .B(n_125), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_149), .B(n_112), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_164), .B(n_127), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_145), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_158), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_141), .B(n_94), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_141), .B(n_126), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_153), .B(n_90), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_163), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_148), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_131), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_153), .B(n_94), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_146), .B(n_123), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_140), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_137), .B(n_120), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_131), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_131), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_146), .B(n_121), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_148), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_147), .B(n_107), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_131), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_129), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_131), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_137), .Y(n_220) );
AND2x6_ASAP7_75t_L g221 ( .A(n_170), .B(n_119), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_147), .B(n_114), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_150), .B(n_111), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_133), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_150), .B(n_116), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_133), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_152), .B(n_109), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_152), .B(n_165), .Y(n_228) );
NAND3xp33_ASAP7_75t_L g229 ( .A(n_136), .B(n_80), .C(n_117), .Y(n_229) );
INVxp67_ASAP7_75t_SL g230 ( .A(n_140), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_154), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_159), .B(n_110), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_154), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_159), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_155), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_193), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_198), .A2(n_165), .B1(n_169), .B2(n_168), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_176), .B(n_169), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_177), .B(n_168), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_201), .B(n_160), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_204), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_180), .B(n_160), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
AND2x2_ASAP7_75t_SL g245 ( .A(n_200), .B(n_166), .Y(n_245) );
NOR3xp33_ASAP7_75t_SL g246 ( .A(n_218), .B(n_132), .C(n_130), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_180), .B(n_170), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_188), .B(n_167), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_182), .Y(n_250) );
BUFx12f_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_186), .B(n_151), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_199), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_173), .A2(n_156), .B1(n_167), .B2(n_105), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_187), .Y(n_256) );
AND3x1_ASAP7_75t_L g257 ( .A(n_196), .B(n_9), .C(n_10), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_193), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
BUFx8_ASAP7_75t_L g260 ( .A(n_200), .Y(n_260) );
OR2x2_ASAP7_75t_SL g261 ( .A(n_235), .B(n_117), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_203), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_204), .B(n_167), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_229), .B(n_9), .Y(n_264) );
OAI221xp5_ASAP7_75t_L g265 ( .A1(n_184), .A2(n_117), .B1(n_144), .B2(n_134), .C(n_133), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_196), .B(n_10), .Y(n_266) );
BUFx2_ASAP7_75t_R g267 ( .A(n_235), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_210), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_208), .B(n_157), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_208), .B(n_157), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_194), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_232), .B(n_211), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_173), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_211), .B(n_157), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_194), .B(n_157), .Y(n_275) );
INVx5_ASAP7_75t_L g276 ( .A(n_198), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_198), .Y(n_277) );
AND2x6_ASAP7_75t_SL g278 ( .A(n_190), .B(n_11), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_230), .A2(n_157), .B(n_144), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_211), .B(n_11), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_187), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_191), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_198), .A2(n_157), .B1(n_144), .B2(n_134), .Y(n_283) );
OR2x2_ASAP7_75t_SL g284 ( .A(n_195), .B(n_13), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_211), .B(n_144), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_234), .B(n_144), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_197), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_203), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_234), .B(n_144), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_210), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_198), .Y(n_291) );
INVx5_ASAP7_75t_L g292 ( .A(n_198), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_198), .A2(n_134), .B1(n_133), .B2(n_15), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_206), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_191), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_174), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_194), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_174), .Y(n_298) );
OAI22xp5_ASAP7_75t_SL g299 ( .A1(n_225), .A2(n_13), .B1(n_14), .B2(n_16), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_194), .B(n_134), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_194), .B(n_134), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_228), .B(n_134), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_194), .B(n_133), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_175), .B1(n_192), .B2(n_220), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_260), .Y(n_305) );
AND2x6_ASAP7_75t_L g306 ( .A(n_277), .B(n_175), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_276), .B(n_220), .Y(n_308) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_252), .A2(n_192), .B(n_209), .C(n_202), .Y(n_309) );
BUFx4f_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_248), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_272), .B(n_192), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_260), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_247), .A2(n_221), .B1(n_206), .B2(n_215), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_242), .B(n_227), .Y(n_316) );
AND2x4_ASAP7_75t_L g317 ( .A(n_266), .B(n_222), .Y(n_317) );
BUFx2_ASAP7_75t_R g318 ( .A(n_267), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_269), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_270), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g321 ( .A(n_276), .B(n_233), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_248), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_277), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_277), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_252), .A2(n_221), .B1(n_216), .B2(n_214), .Y(n_325) );
O2A1O1Ixp5_ASAP7_75t_L g326 ( .A1(n_279), .A2(n_223), .B(n_231), .C(n_233), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_238), .A2(n_239), .B(n_241), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_243), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_263), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_254), .Y(n_331) );
O2A1O1Ixp5_ASAP7_75t_L g332 ( .A1(n_249), .A2(n_231), .B(n_215), .C(n_213), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_273), .A2(n_205), .B(n_183), .C(n_185), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_240), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_273), .B(n_221), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_237), .A2(n_178), .B1(n_183), .B2(n_185), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_247), .B(n_221), .Y(n_337) );
INVxp67_ASAP7_75t_SL g338 ( .A(n_291), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_240), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_237), .A2(n_205), .B1(n_178), .B2(n_189), .Y(n_340) );
INVx2_ASAP7_75t_SL g341 ( .A(n_260), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_247), .B(n_221), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_276), .B(n_189), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_255), .A2(n_221), .B1(n_133), .B2(n_213), .C(n_219), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_245), .B(n_221), .Y(n_345) );
AOI21xp33_ASAP7_75t_L g346 ( .A1(n_245), .A2(n_17), .B(n_19), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
INVx1_ASAP7_75t_SL g348 ( .A(n_251), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_259), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_261), .Y(n_350) );
BUFx4_ASAP7_75t_SL g351 ( .A(n_278), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_291), .Y(n_352) );
INVx2_ASAP7_75t_SL g353 ( .A(n_264), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_291), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g355 ( .A1(n_264), .A2(n_219), .B1(n_217), .B2(n_207), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_284), .B(n_20), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_271), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_347), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_347), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_314), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
OAI21x1_ASAP7_75t_SL g362 ( .A1(n_307), .A2(n_293), .B(n_244), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_309), .A2(n_332), .B(n_327), .Y(n_363) );
NAND3xp33_ASAP7_75t_L g364 ( .A(n_309), .B(n_257), .C(n_293), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_349), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_319), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_332), .A2(n_253), .B(n_256), .Y(n_368) );
OAI21x1_ASAP7_75t_SL g369 ( .A1(n_307), .A2(n_253), .B(n_256), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_264), .B1(n_299), .B2(n_287), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_334), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_316), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_323), .Y(n_373) );
OAI21x1_ASAP7_75t_SL g374 ( .A1(n_304), .A2(n_250), .B(n_282), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_326), .A2(n_286), .B(n_289), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_320), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_328), .B(n_288), .Y(n_377) );
CKINVDCx9p33_ASAP7_75t_R g378 ( .A(n_318), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_326), .A2(n_302), .B(n_274), .Y(n_379) );
INVx3_ASAP7_75t_SL g380 ( .A(n_305), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_329), .B(n_262), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_313), .Y(n_384) );
OAI21x1_ASAP7_75t_L g385 ( .A1(n_355), .A2(n_285), .B(n_303), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_341), .B(n_294), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_325), .B(n_282), .Y(n_387) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_355), .A2(n_281), .B(n_250), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_312), .B(n_281), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_337), .B(n_295), .Y(n_390) );
INVx2_ASAP7_75t_SL g391 ( .A(n_306), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_364), .A2(n_356), .B1(n_350), .B2(n_310), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_370), .A2(n_246), .B(n_315), .C(n_346), .Y(n_393) );
INVx6_ASAP7_75t_L g394 ( .A(n_386), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
OAI222xp33_ASAP7_75t_L g397 ( .A1(n_367), .A2(n_344), .B1(n_353), .B2(n_345), .C1(n_315), .C2(n_348), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_377), .A2(n_342), .B1(n_291), .B2(n_317), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_361), .A2(n_317), .B1(n_310), .B2(n_322), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_372), .A2(n_311), .B1(n_306), .B2(n_357), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_384), .B(n_295), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_365), .Y(n_403) );
OA21x2_ASAP7_75t_L g404 ( .A1(n_363), .A2(n_283), .B(n_275), .Y(n_404) );
AOI22xp33_ASAP7_75t_SL g405 ( .A1(n_364), .A2(n_306), .B1(n_265), .B2(n_351), .Y(n_405) );
OAI21xp33_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_336), .B(n_340), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_381), .B(n_357), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_384), .A2(n_306), .B1(n_290), .B2(n_258), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_381), .B(n_296), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_367), .A2(n_306), .B1(n_292), .B2(n_276), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_376), .A2(n_236), .B1(n_258), .B2(n_268), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_376), .A2(n_333), .B1(n_308), .B2(n_321), .C(n_303), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_377), .A2(n_338), .B(n_292), .C(n_236), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_386), .B(n_296), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_360), .A2(n_292), .B1(n_271), .B2(n_338), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_387), .A2(n_292), .B1(n_352), .B2(n_330), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_380), .A2(n_308), .B1(n_321), .B2(n_275), .C(n_301), .Y(n_419) );
OAI22xp33_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_351), .B1(n_324), .B2(n_352), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_392), .A2(n_362), .B1(n_374), .B2(n_380), .Y(n_421) );
INVx4_ASAP7_75t_L g422 ( .A(n_395), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_396), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_402), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_409), .B(n_358), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_403), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_412), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_413), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_401), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_395), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_416), .B(n_359), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_395), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_401), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g434 ( .A1(n_405), .A2(n_358), .B(n_359), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_400), .B(n_391), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_394), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_394), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_398), .B(n_359), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_398), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_393), .B(n_371), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_399), .B(n_371), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_406), .B(n_371), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_420), .B(n_383), .Y(n_444) );
INVx2_ASAP7_75t_R g445 ( .A(n_404), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_404), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_414), .B(n_383), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_417), .B(n_382), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_411), .A2(n_362), .B1(n_374), .B2(n_387), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_418), .Y(n_451) );
INVx4_ASAP7_75t_R g452 ( .A(n_397), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_410), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_408), .B(n_383), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_415), .B(n_389), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_425), .B(n_368), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_421), .A2(n_378), .B1(n_368), .B2(n_382), .C(n_388), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_431), .B(n_388), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_423), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_431), .B(n_385), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_423), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_426), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_425), .B(n_390), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_424), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_426), .B(n_385), .Y(n_466) );
NAND2x1_ASAP7_75t_L g467 ( .A(n_422), .B(n_369), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_427), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_429), .B(n_390), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_427), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_428), .B(n_385), .Y(n_471) );
BUFx2_ASAP7_75t_L g472 ( .A(n_430), .Y(n_472) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_422), .B(n_382), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_428), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_436), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_439), .B(n_389), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_435), .B(n_391), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_439), .B(n_379), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_436), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_443), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_424), .B(n_379), .Y(n_481) );
BUFx2_ASAP7_75t_L g482 ( .A(n_430), .Y(n_482) );
INVx5_ASAP7_75t_L g483 ( .A(n_430), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_437), .Y(n_484) );
OR2x6_ASAP7_75t_L g485 ( .A(n_447), .B(n_369), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_455), .A2(n_382), .B1(n_391), .B2(n_373), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_429), .B(n_379), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_433), .B(n_375), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_455), .A2(n_373), .B1(n_290), .B2(n_268), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_424), .B(n_375), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_436), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_433), .B(n_375), .Y(n_492) );
BUFx2_ASAP7_75t_L g493 ( .A(n_430), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_437), .B(n_301), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_438), .B(n_22), .Y(n_495) );
BUFx2_ASAP7_75t_L g496 ( .A(n_430), .Y(n_496) );
INVx1_ASAP7_75t_SL g497 ( .A(n_438), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_440), .B(n_23), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_446), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_435), .B(n_26), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_438), .Y(n_501) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_446), .A2(n_343), .B(n_300), .Y(n_502) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_446), .A2(n_207), .B(n_217), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_443), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_440), .B(n_442), .Y(n_505) );
OR2x6_ASAP7_75t_L g506 ( .A(n_447), .B(n_354), .Y(n_506) );
NOR2xp67_ASAP7_75t_L g507 ( .A(n_483), .B(n_422), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_458), .B(n_434), .C(n_449), .Y(n_508) );
INVxp67_ASAP7_75t_L g509 ( .A(n_479), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_505), .A2(n_455), .B1(n_456), .B2(n_442), .Y(n_510) );
AOI211xp5_ASAP7_75t_L g511 ( .A1(n_497), .A2(n_434), .B(n_441), .C(n_435), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_505), .B(n_441), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_476), .B(n_444), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_475), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_462), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_465), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_475), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_500), .A2(n_456), .B1(n_453), .B2(n_435), .Y(n_520) );
INVx1_ASAP7_75t_SL g521 ( .A(n_491), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_476), .B(n_432), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_484), .B(n_432), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_463), .B(n_448), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_468), .B(n_444), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_467), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_470), .Y(n_527) );
NOR2xp67_ASAP7_75t_L g528 ( .A(n_483), .B(n_422), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_467), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_474), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_466), .B(n_448), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g532 ( .A(n_500), .B(n_452), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_459), .B(n_432), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_501), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_466), .B(n_447), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_471), .B(n_451), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_471), .B(n_451), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_464), .B(n_451), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_459), .B(n_453), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_477), .B(n_453), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_487), .Y(n_541) );
INVx2_ASAP7_75t_SL g542 ( .A(n_491), .Y(n_542) );
AOI221xp5_ASAP7_75t_L g543 ( .A1(n_480), .A2(n_504), .B1(n_478), .B2(n_461), .C(n_492), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_487), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_488), .Y(n_545) );
AND2x4_ASAP7_75t_SL g546 ( .A(n_500), .B(n_430), .Y(n_546) );
OAI33xp33_ASAP7_75t_L g547 ( .A1(n_480), .A2(n_452), .A3(n_445), .B1(n_450), .B2(n_343), .B3(n_454), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_464), .B(n_454), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_473), .B(n_354), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_488), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_461), .B(n_445), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_492), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_477), .B(n_445), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_504), .B(n_301), .Y(n_554) );
INVx4_ASAP7_75t_SL g555 ( .A(n_485), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_498), .B(n_27), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_457), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_498), .B(n_31), .Y(n_558) );
NAND3xp33_ASAP7_75t_L g559 ( .A(n_495), .B(n_179), .C(n_212), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_477), .B(n_32), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_457), .B(n_33), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_469), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_469), .B(n_34), .Y(n_563) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_486), .B(n_36), .C(n_39), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_481), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g566 ( .A(n_507), .B(n_483), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_513), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_517), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_522), .B(n_478), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_514), .Y(n_570) );
NAND4xp75_ASAP7_75t_L g571 ( .A(n_528), .B(n_481), .C(n_490), .D(n_499), .Y(n_571) );
NAND2x1p5_ASAP7_75t_L g572 ( .A(n_519), .B(n_483), .Y(n_572) );
NAND2x1_ASAP7_75t_L g573 ( .A(n_526), .B(n_485), .Y(n_573) );
AND2x6_ASAP7_75t_L g574 ( .A(n_519), .B(n_490), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_548), .B(n_493), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_527), .Y(n_576) );
OAI21xp33_ASAP7_75t_L g577 ( .A1(n_508), .A2(n_485), .B(n_489), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_562), .B(n_494), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_533), .B(n_472), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_515), .B(n_512), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_516), .B(n_472), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_557), .B(n_524), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_509), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_530), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_524), .B(n_499), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_534), .Y(n_586) );
OAI211xp5_ASAP7_75t_L g587 ( .A1(n_532), .A2(n_494), .B(n_483), .C(n_496), .Y(n_587) );
AND2x4_ASAP7_75t_L g588 ( .A(n_555), .B(n_485), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_521), .B(n_496), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_552), .B(n_493), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_555), .B(n_482), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_542), .B(n_482), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_521), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_559), .A2(n_506), .B(n_502), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_543), .B(n_502), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_555), .B(n_506), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_543), .B(n_502), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_565), .B(n_506), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_526), .B(n_354), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_523), .B(n_506), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_541), .B(n_503), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_518), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_525), .Y(n_603) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_529), .B(n_503), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_544), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_551), .B(n_503), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_545), .B(n_503), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_550), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_41), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_539), .B(n_42), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_531), .B(n_44), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_538), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_531), .Y(n_613) );
INVx3_ASAP7_75t_L g614 ( .A(n_529), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_535), .B(n_55), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_540), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_535), .B(n_300), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_536), .B(n_300), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_613), .B(n_510), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_566), .B(n_511), .Y(n_621) );
NOR2x1_ASAP7_75t_L g622 ( .A(n_571), .B(n_564), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g623 ( .A1(n_566), .A2(n_520), .B1(n_563), .B2(n_561), .Y(n_623) );
AOI222xp33_ASAP7_75t_L g624 ( .A1(n_577), .A2(n_547), .B1(n_537), .B2(n_536), .C1(n_540), .C2(n_560), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_583), .B(n_558), .C(n_556), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_587), .A2(n_546), .B1(n_553), .B2(n_537), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_577), .A2(n_553), .B1(n_564), .B2(n_554), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g628 ( .A1(n_617), .A2(n_549), .B1(n_330), .B2(n_179), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_567), .Y(n_629) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_593), .B(n_549), .C(n_59), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_572), .A2(n_354), .B1(n_323), .B2(n_297), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_574), .B(n_56), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_593), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_572), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_580), .B(n_63), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_618), .B(n_298), .C(n_69), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_576), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_602), .Y(n_641) );
NOR3xp33_ASAP7_75t_L g642 ( .A(n_618), .B(n_298), .C(n_70), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_573), .A2(n_323), .B(n_297), .C(n_74), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_584), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_581), .Y(n_645) );
INVx2_ASAP7_75t_L g646 ( .A(n_606), .Y(n_646) );
OAI322xp33_ASAP7_75t_L g647 ( .A1(n_595), .A2(n_212), .A3(n_226), .B1(n_224), .B2(n_179), .C1(n_65), .C2(n_77), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g648 ( .A1(n_588), .A2(n_71), .A3(n_323), .B(n_297), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_612), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_603), .B(n_179), .Y(n_650) );
AND2x4_ASAP7_75t_L g651 ( .A(n_574), .B(n_179), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_588), .A2(n_297), .B1(n_224), .B2(n_226), .Y(n_652) );
NOR2xp33_ASAP7_75t_SL g653 ( .A(n_574), .B(n_226), .Y(n_653) );
NOR2x1_ASAP7_75t_L g654 ( .A(n_614), .B(n_212), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_582), .B(n_212), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_592), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_605), .B(n_212), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_653), .B(n_591), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_632), .B(n_591), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_620), .B(n_608), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_633), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_644), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_629), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_649), .B(n_569), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_624), .B(n_575), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g666 ( .A(n_632), .B(n_614), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_635), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_646), .B(n_579), .Y(n_668) );
NOR2xp67_ASAP7_75t_SL g669 ( .A(n_625), .B(n_611), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_639), .B(n_595), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_640), .Y(n_671) );
AOI21xp33_ASAP7_75t_L g672 ( .A1(n_622), .A2(n_597), .B(n_615), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_625), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_637), .B(n_597), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_645), .B(n_656), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_641), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_634), .B(n_589), .Y(n_677) );
NOR3x1_ASAP7_75t_L g678 ( .A(n_621), .B(n_590), .C(n_604), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g679 ( .A1(n_648), .A2(n_630), .B(n_627), .C(n_643), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_650), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_626), .A2(n_596), .B1(n_609), .B2(n_610), .Y(n_681) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_679), .B(n_651), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_661), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_676), .Y(n_684) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_679), .A2(n_648), .B(n_642), .Y(n_685) );
OAI21xp5_ASAP7_75t_L g686 ( .A1(n_673), .A2(n_669), .B(n_665), .Y(n_686) );
XOR2x2_ASAP7_75t_L g687 ( .A(n_659), .B(n_623), .Y(n_687) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_681), .A2(n_636), .B(n_651), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_674), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_662), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_663), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_658), .B(n_638), .C(n_594), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_670), .B(n_585), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_675), .B(n_616), .Y(n_694) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_672), .A2(n_578), .A3(n_598), .B1(n_596), .B2(n_600), .C1(n_619), .C2(n_654), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_685), .B(n_647), .C(n_658), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_686), .A2(n_660), .B1(n_667), .B2(n_671), .C(n_680), .Y(n_697) );
OAI21xp5_ASAP7_75t_SL g698 ( .A1(n_682), .A2(n_659), .B(n_666), .Y(n_698) );
A2O1A1Ixp33_ASAP7_75t_L g699 ( .A1(n_695), .A2(n_666), .B(n_661), .C(n_678), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_687), .A2(n_664), .B(n_677), .Y(n_700) );
NAND4xp25_ASAP7_75t_L g701 ( .A(n_692), .B(n_628), .C(n_619), .D(n_655), .Y(n_701) );
AOI211xp5_ASAP7_75t_SL g702 ( .A1(n_688), .A2(n_647), .B(n_652), .C(n_631), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_689), .A2(n_668), .B1(n_657), .B2(n_601), .C(n_607), .Y(n_703) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_698), .B(n_687), .Y(n_704) );
OR5x1_ASAP7_75t_L g705 ( .A(n_699), .B(n_683), .C(n_689), .D(n_694), .E(n_690), .Y(n_705) );
NOR2x1_ASAP7_75t_L g706 ( .A(n_700), .B(n_684), .Y(n_706) );
NAND4xp25_ASAP7_75t_L g707 ( .A(n_696), .B(n_691), .C(n_694), .D(n_693), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_697), .B(n_684), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_706), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_704), .B(n_703), .Y(n_710) );
OR4x2_ASAP7_75t_L g711 ( .A(n_705), .B(n_702), .C(n_701), .D(n_574), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_709), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_710), .B(n_708), .Y(n_713) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_712), .A2(n_711), .B1(n_707), .B2(n_607), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_713), .A2(n_711), .B1(n_668), .B2(n_599), .Y(n_715) );
XOR2xp5_ASAP7_75t_L g716 ( .A(n_714), .B(n_601), .Y(n_716) );
XOR2xp5_ASAP7_75t_L g717 ( .A(n_716), .B(n_715), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_224), .B1(n_226), .B2(n_713), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_224), .B(n_226), .Y(n_719) );
endmodule