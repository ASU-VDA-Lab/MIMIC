module fake_netlist_6_1369_n_2413 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2413);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2413;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_873;
wire n_461;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_1070;
wire n_458;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_235),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_40),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_143),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_36),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_29),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_47),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_49),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_234),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_34),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_142),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_161),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_123),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_33),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_181),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_85),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_162),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_118),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_57),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_81),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_36),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_27),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_62),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_190),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_136),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_150),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_9),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_139),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_70),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_74),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_179),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_66),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_109),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_87),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_54),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_184),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_39),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_26),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_165),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_94),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_73),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_57),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_216),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_200),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_62),
.Y(n_289)
);

INVxp33_ASAP7_75t_R g290 ( 
.A(n_156),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_2),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_85),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_222),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_215),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_41),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_22),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_180),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_19),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_60),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_236),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_229),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_131),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_152),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_186),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_86),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_12),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_127),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_31),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_155),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_105),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_23),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_15),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_82),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_126),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_206),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_99),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_40),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_64),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_50),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_171),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_145),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_31),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_220),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_132),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_27),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_135),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_209),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_10),
.Y(n_329)
);

BUFx10_ASAP7_75t_L g330 ( 
.A(n_232),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_176),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_141),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_55),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_74),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_96),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_230),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_21),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_43),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_0),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_91),
.Y(n_340)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_196),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_61),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_144),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_29),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_43),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_148),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_96),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_199),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_108),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_54),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_140),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_7),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_124),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_100),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_89),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_56),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_170),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_233),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_5),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_18),
.Y(n_360)
);

BUFx10_ASAP7_75t_L g361 ( 
.A(n_63),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_82),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_98),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_84),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_34),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_174),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_41),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_147),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_88),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_97),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_67),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_87),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_114),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_75),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_78),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_192),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_178),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_50),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_42),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_65),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_154),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_117),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_204),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_159),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_33),
.Y(n_385)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_23),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_94),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_104),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_212),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_15),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_207),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_92),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_1),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_104),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_26),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_6),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_2),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_3),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_46),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_198),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_95),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_78),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_86),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_112),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_81),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_191),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_20),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_130),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_21),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_172),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_59),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_107),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_98),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_60),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_91),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_97),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_208),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_80),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_6),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_63),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_47),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_214),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_24),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_202),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_72),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_95),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_115),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_59),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_32),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_7),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_221),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_138),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_163),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_5),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_195),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_37),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_219),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_88),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_1),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_77),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_0),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_164),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_13),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_73),
.Y(n_444)
);

BUFx10_ASAP7_75t_L g445 ( 
.A(n_175),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_167),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_188),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_61),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_185),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_103),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_51),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_75),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_137),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_64),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_146),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_80),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_55),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_46),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_224),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_99),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_44),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_65),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_228),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_111),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_289),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_237),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_289),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_310),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_244),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_289),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_289),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_274),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_305),
.B(n_3),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_289),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_289),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_289),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_246),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_242),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_289),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_247),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_289),
.Y(n_481)
);

CKINVDCx14_ASAP7_75t_R g482 ( 
.A(n_274),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_248),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_305),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_250),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_420),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_327),
.B(n_4),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_409),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_348),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_420),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_251),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_420),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_420),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_411),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_450),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_450),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_254),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_349),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_353),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_327),
.B(n_4),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_450),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_260),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_450),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_411),
.B(n_256),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g509 ( 
.A(n_256),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_263),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_295),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_295),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_357),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_295),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_266),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_456),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_242),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_268),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_R g519 ( 
.A(n_368),
.B(n_106),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_366),
.B(n_8),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_381),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_366),
.B(n_8),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_456),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_282),
.Y(n_525)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_273),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_406),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_408),
.B(n_9),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_240),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_293),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_300),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_424),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_312),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_301),
.Y(n_534)
);

INVxp67_ASAP7_75t_SL g535 ( 
.A(n_408),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_446),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_312),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_455),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_302),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_464),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_313),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_313),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_309),
.B(n_10),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_256),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_273),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_303),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_243),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_307),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_R g549 ( 
.A(n_387),
.B(n_309),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_371),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_371),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_314),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_238),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_389),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_328),
.Y(n_555)
);

CKINVDCx16_ASAP7_75t_R g556 ( 
.A(n_389),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_371),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_431),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_309),
.B(n_11),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_315),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_238),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_241),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_431),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_432),
.Y(n_564)
);

INVxp33_ASAP7_75t_SL g565 ( 
.A(n_245),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_241),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_252),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_252),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_316),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_267),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_267),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_275),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_361),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_321),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_322),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_275),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_249),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_432),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_324),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_447),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_447),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_276),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_276),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_280),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_280),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_331),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_332),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_259),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_453),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_453),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_291),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_291),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_468),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_466),
.B(n_464),
.Y(n_594)
);

NAND2x1_ASAP7_75t_L g595 ( 
.A(n_543),
.B(n_309),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_486),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_469),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_486),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_477),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_480),
.Y(n_601)
);

BUFx3_ASAP7_75t_L g602 ( 
.A(n_540),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_483),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_485),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_493),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_517),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

CKINVDCx16_ASAP7_75t_R g608 ( 
.A(n_478),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_555),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_500),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_558),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_505),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_510),
.B(n_464),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_487),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_482),
.B(n_386),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_515),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_555),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_518),
.Y(n_620)
);

NAND3xp33_ASAP7_75t_L g621 ( 
.A(n_488),
.B(n_306),
.C(n_296),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

CKINVDCx20_ASAP7_75t_R g623 ( 
.A(n_490),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_555),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_525),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_478),
.A2(n_311),
.B1(n_318),
.B2(n_262),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_472),
.A2(n_329),
.B1(n_270),
.B2(n_272),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_474),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_487),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_530),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_491),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_531),
.B(n_271),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_474),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_559),
.A2(n_253),
.B(n_239),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_534),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_539),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_491),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_492),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_492),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_495),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_546),
.B(n_271),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_540),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_495),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_548),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_497),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_497),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_498),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_498),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_501),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_511),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_552),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_565),
.B(n_358),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_499),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_560),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_499),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_521),
.B(n_523),
.C(n_503),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_504),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_504),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_506),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_506),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_465),
.B(n_283),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_569),
.B(n_463),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_507),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_507),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_574),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_511),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_575),
.B(n_343),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_579),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_502),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_586),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_514),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_587),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_513),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_514),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_535),
.B(n_239),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_465),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_467),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_467),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_470),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_561),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_508),
.B(n_346),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_470),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_561),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_562),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_471),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_471),
.B(n_304),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_475),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_562),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_658),
.A2(n_549),
.B1(n_545),
.B2(n_526),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_628),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_680),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_678),
.Y(n_694)
);

OAI21xp33_ASAP7_75t_L g695 ( 
.A1(n_677),
.A2(n_473),
.B(n_528),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_675),
.Y(n_696)
);

AO22x2_ASAP7_75t_L g697 ( 
.A1(n_621),
.A2(n_473),
.B1(n_627),
.B2(n_304),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_644),
.B(n_475),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_632),
.B(n_643),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_602),
.B(n_544),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_679),
.Y(n_701)
);

AND2x6_ASAP7_75t_L g702 ( 
.A(n_688),
.B(n_304),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_602),
.B(n_476),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_602),
.B(n_476),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_679),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_678),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_594),
.B(n_526),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_640),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_613),
.B(n_479),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_683),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_664),
.B(n_669),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_680),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_680),
.Y(n_713)
);

AND2x2_ASAP7_75t_SL g714 ( 
.A(n_634),
.B(n_545),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_640),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_654),
.B(n_556),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_628),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_684),
.Y(n_718)
);

BUFx10_ASAP7_75t_L g719 ( 
.A(n_617),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_597),
.B(n_556),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_628),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_640),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_665),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_684),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_593),
.Y(n_725)
);

NOR3xp33_ASAP7_75t_L g726 ( 
.A(n_626),
.B(n_581),
.C(n_496),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_600),
.B(n_581),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_684),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_678),
.B(n_479),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_687),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_601),
.B(n_603),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_687),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_604),
.B(n_519),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_665),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_628),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_665),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_614),
.A2(n_489),
.B1(n_564),
.B2(n_563),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_682),
.B(n_508),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_605),
.B(n_577),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_628),
.Y(n_740)
);

AO21x2_ASAP7_75t_L g741 ( 
.A1(n_663),
.A2(n_258),
.B(n_253),
.Y(n_741)
);

INVx6_ASAP7_75t_L g742 ( 
.A(n_628),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_623),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_678),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_622),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_687),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_682),
.B(n_544),
.Y(n_747)
);

XNOR2xp5_ASAP7_75t_L g748 ( 
.A(n_626),
.B(n_522),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_663),
.B(n_481),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_621),
.A2(n_400),
.B1(n_384),
.B2(n_306),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_689),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_688),
.B(n_550),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_689),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_633),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_610),
.B(n_573),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_633),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_606),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_612),
.B(n_588),
.Y(n_758)
);

OR2x2_ASAP7_75t_L g759 ( 
.A(n_608),
.B(n_588),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_618),
.B(n_573),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_595),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_633),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_620),
.B(n_578),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_689),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_625),
.B(n_580),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_L g766 ( 
.A(n_679),
.B(n_328),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_630),
.B(n_589),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_679),
.B(n_481),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_679),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_651),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_679),
.Y(n_771)
);

INVx4_ASAP7_75t_L g772 ( 
.A(n_681),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_681),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_681),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_608),
.B(n_496),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_681),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_688),
.B(n_550),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_636),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_685),
.B(n_551),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_646),
.A2(n_257),
.B1(n_405),
.B2(n_261),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_611),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_633),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_596),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_596),
.Y(n_784)
);

INVx6_ASAP7_75t_L g785 ( 
.A(n_633),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_671),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_598),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_598),
.Y(n_788)
);

INVx1_ASAP7_75t_SL g789 ( 
.A(n_611),
.Y(n_789)
);

BUFx10_ASAP7_75t_L g790 ( 
.A(n_653),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_615),
.Y(n_791)
);

AND2x6_ASAP7_75t_L g792 ( 
.A(n_688),
.B(n_384),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_607),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_681),
.B(n_633),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_681),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_648),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_615),
.Y(n_797)
);

AND2x6_ASAP7_75t_L g798 ( 
.A(n_685),
.B(n_384),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_686),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_656),
.B(n_590),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_595),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_667),
.B(n_484),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_670),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_648),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_648),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_607),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_629),
.B(n_551),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_629),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_634),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_672),
.B(n_255),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_686),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_631),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_648),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_631),
.B(n_557),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_690),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_690),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_637),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_637),
.B(n_557),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_638),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_638),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_639),
.B(n_376),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_648),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_634),
.B(n_509),
.Y(n_823)
);

AO22x2_ASAP7_75t_L g824 ( 
.A1(n_634),
.A2(n_400),
.B1(n_319),
.B2(n_326),
.Y(n_824)
);

BUFx4f_ASAP7_75t_L g825 ( 
.A(n_648),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_674),
.Y(n_826)
);

INVxp67_ASAP7_75t_SL g827 ( 
.A(n_624),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_639),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_641),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_641),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_642),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_668),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_642),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_645),
.B(n_377),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_645),
.Y(n_835)
);

AND2x6_ASAP7_75t_L g836 ( 
.A(n_599),
.B(n_400),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_661),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_647),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_647),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_661),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_649),
.Y(n_841)
);

CKINVDCx11_ASAP7_75t_R g842 ( 
.A(n_668),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_649),
.B(n_509),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_650),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_650),
.A2(n_319),
.B1(n_326),
.B2(n_296),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_673),
.Y(n_846)
);

OR2x6_ASAP7_75t_L g847 ( 
.A(n_676),
.B(n_290),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_655),
.B(n_383),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_655),
.B(n_404),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_657),
.B(n_527),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_657),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_659),
.B(n_512),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_710),
.B(n_532),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_699),
.B(n_536),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_716),
.B(n_572),
.C(n_553),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_828),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_710),
.B(n_659),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_709),
.B(n_660),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_828),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_711),
.B(n_660),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_783),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_783),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_829),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_714),
.A2(n_538),
.B1(n_258),
.B2(n_265),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_833),
.B(n_698),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_707),
.B(n_290),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_806),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_829),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_691),
.B(n_695),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_739),
.B(n_269),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_847),
.B(n_264),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_803),
.B(n_372),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_823),
.A2(n_264),
.B1(n_279),
.B2(n_265),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_784),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_830),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_784),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_833),
.B(n_761),
.Y(n_877)
);

CKINVDCx11_ASAP7_75t_R g878 ( 
.A(n_790),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_702),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_757),
.B(n_277),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_761),
.B(n_703),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_704),
.B(n_662),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_696),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_832),
.B(n_410),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_714),
.B(n_412),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_850),
.B(n_417),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_830),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_831),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_823),
.A2(n_697),
.B1(n_777),
.B2(n_752),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_702),
.B(n_341),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_802),
.B(n_278),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_787),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_752),
.B(n_662),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_752),
.B(n_666),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_777),
.B(n_666),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_806),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_697),
.A2(n_435),
.B1(n_437),
.B2(n_427),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_787),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_777),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_799),
.B(n_624),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_831),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_851),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_702),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_811),
.B(n_624),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_738),
.B(n_585),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_697),
.A2(n_449),
.B1(n_459),
.B2(n_442),
.Y(n_906)
);

NOR2x1p5_ASAP7_75t_L g907 ( 
.A(n_775),
.B(n_281),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_758),
.B(n_255),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_735),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_851),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_700),
.B(n_733),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_788),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_815),
.B(n_624),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_809),
.A2(n_340),
.B(n_365),
.C(n_334),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_700),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_816),
.B(n_661),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_801),
.B(n_661),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_801),
.B(n_661),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_755),
.B(n_760),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_852),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_809),
.B(n_279),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_845),
.A2(n_340),
.B1(n_419),
.B2(n_416),
.C(n_415),
.Y(n_922)
);

OR2x2_ASAP7_75t_L g923 ( 
.A(n_775),
.B(n_566),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_846),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_700),
.B(n_661),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_788),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_791),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_738),
.B(n_255),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_843),
.B(n_255),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_747),
.B(n_566),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_824),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_819),
.B(n_599),
.Y(n_932)
);

AND2x6_ASAP7_75t_SL g933 ( 
.A(n_847),
.B(n_334),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_820),
.B(n_599),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_791),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_835),
.B(n_609),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_841),
.B(n_609),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_824),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_794),
.A2(n_616),
.B(n_609),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_797),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_L g941 ( 
.A(n_702),
.B(n_341),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_844),
.B(n_616),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_797),
.Y(n_943)
);

AO22x1_ASAP7_75t_L g944 ( 
.A1(n_798),
.A2(n_288),
.B1(n_294),
.B2(n_287),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_808),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_694),
.B(n_616),
.Y(n_946)
);

BUFx3_ASAP7_75t_L g947 ( 
.A(n_846),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_808),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_697),
.A2(n_288),
.B1(n_294),
.B2(n_287),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_852),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_706),
.B(n_619),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_812),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_727),
.B(n_330),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_702),
.A2(n_325),
.B1(n_336),
.B2(n_297),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_812),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_744),
.B(n_619),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_747),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_827),
.B(n_619),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_817),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_821),
.B(n_673),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_817),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_768),
.A2(n_676),
.B(n_652),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_719),
.B(n_330),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_834),
.B(n_297),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_848),
.B(n_325),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_838),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_719),
.B(n_330),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_750),
.A2(n_336),
.B1(n_373),
.B2(n_351),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_L g969 ( 
.A1(n_750),
.A2(n_351),
.B1(n_382),
.B2(n_373),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_849),
.B(n_382),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_838),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_839),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_SL g973 ( 
.A(n_803),
.B(n_399),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_779),
.B(n_567),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_781),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_SL g976 ( 
.A(n_735),
.B(n_328),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_839),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_750),
.A2(n_391),
.B1(n_422),
.B2(n_433),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_745),
.B(n_810),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_751),
.Y(n_980)
);

O2A1O1Ixp5_ASAP7_75t_L g981 ( 
.A1(n_729),
.A2(n_433),
.B(n_422),
.C(n_391),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_719),
.B(n_330),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_759),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_751),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_779),
.B(n_567),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_764),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_749),
.B(n_652),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_750),
.A2(n_328),
.B1(n_341),
.B2(n_457),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_824),
.A2(n_328),
.B1(n_342),
.B2(n_401),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_692),
.B(n_652),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_692),
.B(n_652),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_790),
.B(n_445),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_692),
.B(n_328),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_759),
.B(n_284),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_702),
.A2(n_402),
.B1(n_423),
.B2(n_452),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_792),
.A2(n_341),
.B1(n_413),
.B2(n_365),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_717),
.B(n_341),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_824),
.B(n_568),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_717),
.B(n_341),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_789),
.B(n_568),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_717),
.B(n_341),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_721),
.B(n_341),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_721),
.B(n_740),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_SL g1004 ( 
.A1(n_748),
.A2(n_847),
.B1(n_725),
.B2(n_770),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_731),
.B(n_285),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_721),
.B(n_341),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_852),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_847),
.B(n_369),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_740),
.B(n_512),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_790),
.B(n_445),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_792),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_741),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_740),
.B(n_516),
.Y(n_1013)
);

NOR2xp67_ASAP7_75t_L g1014 ( 
.A(n_778),
.B(n_110),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_693),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_792),
.A2(n_741),
.B1(n_798),
.B2(n_712),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_793),
.B(n_570),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_764),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_826),
.B(n_780),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_792),
.B(n_570),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_720),
.B(n_286),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_792),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_693),
.Y(n_1023)
);

OR2x6_ASAP7_75t_L g1024 ( 
.A(n_763),
.B(n_369),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_756),
.B(n_516),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_756),
.B(n_520),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_SL g1027 ( 
.A(n_741),
.B(n_374),
.Y(n_1027)
);

NOR3xp33_ASAP7_75t_SL g1028 ( 
.A(n_864),
.B(n_298),
.C(n_292),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1000),
.B(n_826),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_860),
.B(n_792),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_865),
.B(n_712),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_861),
.Y(n_1032)
);

OR2x6_ASAP7_75t_L g1033 ( 
.A(n_924),
.B(n_765),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_883),
.B(n_696),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_915),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_861),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_883),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1007),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_915),
.B(n_1007),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_912),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_854),
.A2(n_767),
.B1(n_800),
.B2(n_726),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_1019),
.B(n_308),
.C(n_299),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_867),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_856),
.B(n_713),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_866),
.B(n_737),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_1000),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_975),
.B(n_905),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_912),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_856),
.B(n_713),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_891),
.B(n_748),
.C(n_842),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_935),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_923),
.B(n_725),
.Y(n_1052)
);

INVx5_ASAP7_75t_L g1053 ( 
.A(n_879),
.Y(n_1053)
);

AOI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_869),
.A2(n_889),
.B1(n_885),
.B2(n_870),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1005),
.B(n_807),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_879),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_935),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_905),
.B(n_743),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_920),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_862),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_899),
.Y(n_1061)
);

BUFx4_ASAP7_75t_SL g1062 ( 
.A(n_933),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_1017),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_920),
.B(n_735),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_896),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_949),
.A2(n_798),
.B1(n_374),
.B2(n_397),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_SL g1067 ( 
.A(n_995),
.B(n_770),
.C(n_743),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_920),
.A2(n_798),
.B1(n_773),
.B2(n_774),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_940),
.Y(n_1069)
);

O2A1O1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_931),
.A2(n_818),
.B(n_814),
.C(n_724),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_940),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_878),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_943),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_SL g1074 ( 
.A(n_853),
.B(n_320),
.C(n_317),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_862),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_957),
.B(n_571),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_859),
.B(n_718),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_983),
.B(n_842),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1017),
.Y(n_1079)
);

INVx5_ASAP7_75t_L g1080 ( 
.A(n_879),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_947),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_855),
.B(n_786),
.C(n_333),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_931),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_943),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_878),
.B(n_786),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_859),
.B(n_718),
.Y(n_1086)
);

INVx2_ASAP7_75t_SL g1087 ( 
.A(n_923),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_950),
.B(n_735),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_945),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_863),
.B(n_724),
.Y(n_1090)
);

INVxp67_ASAP7_75t_SL g1091 ( 
.A(n_950),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_863),
.B(n_728),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_968),
.A2(n_798),
.B1(n_380),
.B2(n_413),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_868),
.B(n_728),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_950),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_897),
.A2(n_798),
.B1(n_776),
.B2(n_795),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_945),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_952),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_947),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_874),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1004),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_L g1102 ( 
.A(n_1024),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_952),
.Y(n_1103)
);

OR2x6_ASAP7_75t_L g1104 ( 
.A(n_924),
.B(n_380),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_874),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_938),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_868),
.B(n_730),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_930),
.B(n_571),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_880),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_879),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_875),
.B(n_887),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_857),
.B(n_771),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_875),
.B(n_730),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_R g1114 ( 
.A(n_872),
.B(n_323),
.Y(n_1114)
);

NAND2x1_ASAP7_75t_L g1115 ( 
.A(n_909),
.B(n_742),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1020),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_887),
.B(n_732),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_930),
.B(n_576),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_972),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_994),
.B(n_756),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_1008),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_974),
.B(n_985),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1011),
.B(n_762),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_974),
.B(n_361),
.Y(n_1124)
);

BUFx12f_ASAP7_75t_L g1125 ( 
.A(n_1008),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_877),
.B(n_762),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_972),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_879),
.B(n_735),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_903),
.B(n_754),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1008),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_1024),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_977),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_985),
.B(n_576),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_1020),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_911),
.B(n_582),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_888),
.B(n_732),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_979),
.B(n_361),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_977),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_876),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1015),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1015),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1023),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_888),
.B(n_762),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_901),
.B(n_746),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_901),
.B(n_753),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_906),
.A2(n_742),
.B1(n_785),
.B2(n_769),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_938),
.Y(n_1147)
);

OR2x6_ASAP7_75t_L g1148 ( 
.A(n_871),
.B(n_397),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_903),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_973),
.B(n_337),
.C(n_335),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_902),
.B(n_796),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1023),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_902),
.B(n_796),
.Y(n_1153)
);

INVx4_ASAP7_75t_L g1154 ( 
.A(n_903),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_910),
.B(n_796),
.Y(n_1155)
);

BUFx4f_ASAP7_75t_L g1156 ( 
.A(n_1024),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_876),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1024),
.Y(n_1158)
);

INVxp33_ASAP7_75t_L g1159 ( 
.A(n_1021),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1020),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_892),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_871),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_881),
.A2(n_825),
.B(n_705),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_910),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_998),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_903),
.Y(n_1166)
);

BUFx4_ASAP7_75t_SL g1167 ( 
.A(n_1008),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_858),
.B(n_805),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_919),
.B(n_361),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_SL g1170 ( 
.A(n_903),
.B(n_754),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_884),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_960),
.B(n_805),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_892),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_898),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_898),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1011),
.B(n_582),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_926),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_964),
.B(n_805),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_R g1179 ( 
.A(n_998),
.B(n_338),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_907),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_SL g1181 ( 
.A(n_871),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_928),
.B(n_583),
.Y(n_1182)
);

OR2x2_ASAP7_75t_L g1183 ( 
.A(n_908),
.B(n_583),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_926),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_922),
.B(n_344),
.C(n_339),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_927),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1022),
.Y(n_1187)
);

BUFx5_ASAP7_75t_L g1188 ( 
.A(n_1022),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_965),
.B(n_813),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_927),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_893),
.A2(n_742),
.B1(n_785),
.B2(n_705),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_886),
.B(n_584),
.Y(n_1192)
);

BUFx3_ASAP7_75t_L g1193 ( 
.A(n_894),
.Y(n_1193)
);

OR2x2_ASAP7_75t_L g1194 ( 
.A(n_929),
.B(n_963),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1022),
.B(n_1014),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1022),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_895),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1027),
.A2(n_970),
.B1(n_1012),
.B2(n_873),
.Y(n_1198)
);

AOI22x1_ASAP7_75t_L g1199 ( 
.A1(n_921),
.A2(n_1012),
.B1(n_948),
.B2(n_959),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1022),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_948),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_R g1202 ( 
.A(n_1027),
.B(n_345),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_955),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_871),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_955),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_909),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_959),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_909),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_961),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_921),
.B(n_961),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_966),
.B(n_813),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_992),
.Y(n_1212)
);

OA22x2_ASAP7_75t_L g1213 ( 
.A1(n_978),
.A2(n_415),
.B1(n_416),
.B2(n_419),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1016),
.B(n_966),
.Y(n_1214)
);

NOR2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1010),
.B(n_347),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_921),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_971),
.B(n_813),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_971),
.B(n_584),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_980),
.Y(n_1219)
);

INVx4_ASAP7_75t_L g1220 ( 
.A(n_980),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_R g1221 ( 
.A(n_890),
.B(n_350),
.Y(n_1221)
);

NOR3xp33_ASAP7_75t_SL g1222 ( 
.A(n_967),
.B(n_354),
.C(n_352),
.Y(n_1222)
);

INVx3_ASAP7_75t_SL g1223 ( 
.A(n_982),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1047),
.B(n_953),
.Y(n_1224)
);

HAxp5_ASAP7_75t_L g1225 ( 
.A(n_1215),
.B(n_355),
.CON(n_1225),
.SN(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1035),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1054),
.B(n_917),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1195),
.A2(n_825),
.B(n_918),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1083),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1214),
.A2(n_925),
.B(n_987),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_1056),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1195),
.A2(n_825),
.B(n_705),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1055),
.B(n_969),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1122),
.B(n_916),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1214),
.A2(n_882),
.B(n_958),
.Y(n_1235)
);

BUFx4f_ASAP7_75t_L g1236 ( 
.A(n_1223),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1055),
.B(n_984),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1199),
.A2(n_1163),
.B(n_1210),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1206),
.Y(n_1239)
);

AOI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1045),
.A2(n_914),
.B(n_989),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1143),
.A2(n_939),
.B(n_1003),
.Y(n_1241)
);

CKINVDCx16_ASAP7_75t_R g1242 ( 
.A(n_1034),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1159),
.B(n_1046),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1111),
.A2(n_999),
.B(n_997),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_SL g1245 ( 
.A(n_1053),
.B(n_984),
.Y(n_1245)
);

AO21x1_ASAP7_75t_L g1246 ( 
.A1(n_1120),
.A2(n_1002),
.B(n_1001),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_1034),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1030),
.A2(n_769),
.B(n_701),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1219),
.Y(n_1249)
);

BUFx6f_ASAP7_75t_L g1250 ( 
.A(n_1056),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1029),
.B(n_988),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1122),
.B(n_986),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1083),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1198),
.A2(n_934),
.B(n_932),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_1056),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1219),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1037),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1151),
.A2(n_1006),
.B(n_993),
.Y(n_1258)
);

OAI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1070),
.A2(n_937),
.B(n_936),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1206),
.A2(n_769),
.B(n_701),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1193),
.B(n_986),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1193),
.B(n_1018),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1153),
.A2(n_951),
.B(n_946),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1206),
.A2(n_772),
.B(n_701),
.Y(n_1264)
);

BUFx4_ASAP7_75t_SL g1265 ( 
.A(n_1162),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1197),
.B(n_1018),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1106),
.Y(n_1267)
);

OR2x2_ASAP7_75t_L g1268 ( 
.A(n_1052),
.B(n_1079),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1206),
.A2(n_1208),
.B(n_1168),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1155),
.A2(n_956),
.B(n_942),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_L g1271 ( 
.A(n_1223),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1120),
.A2(n_981),
.B(n_944),
.C(n_904),
.Y(n_1272)
);

NAND2x1p5_ASAP7_75t_L g1273 ( 
.A(n_1053),
.B(n_772),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1197),
.B(n_1009),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1106),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1108),
.B(n_1013),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1043),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1079),
.B(n_900),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1208),
.A2(n_772),
.B(n_890),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1108),
.B(n_1025),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1118),
.B(n_1026),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1063),
.B(n_913),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1208),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1118),
.B(n_990),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1059),
.B(n_954),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1065),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1045),
.A2(n_941),
.B1(n_996),
.B2(n_742),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1056),
.Y(n_1288)
);

AOI31xp67_ASAP7_75t_L g1289 ( 
.A1(n_1096),
.A2(n_736),
.A3(n_708),
.B(n_715),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1112),
.A2(n_962),
.A3(n_991),
.B(n_715),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1172),
.A2(n_1112),
.B(n_1178),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1208),
.A2(n_941),
.B(n_782),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1085),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1044),
.A2(n_1077),
.B(n_1049),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1128),
.A2(n_782),
.B(n_754),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1194),
.B(n_113),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1147),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1032),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1102),
.A2(n_429),
.B(n_441),
.C(n_457),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1149),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1087),
.B(n_591),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1086),
.A2(n_722),
.B(n_708),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1217),
.A2(n_1115),
.B(n_1088),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1059),
.B(n_754),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1126),
.A2(n_722),
.A3(n_723),
.B(n_734),
.Y(n_1305)
);

BUFx2_ASAP7_75t_SL g1306 ( 
.A(n_1099),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1064),
.A2(n_734),
.B(n_723),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_1081),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1216),
.A2(n_785),
.B1(n_754),
.B2(n_782),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1133),
.B(n_944),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1064),
.A2(n_736),
.B(n_524),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1216),
.A2(n_785),
.B1(n_782),
.B2(n_822),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1159),
.B(n_356),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1147),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1088),
.A2(n_524),
.B(n_520),
.Y(n_1315)
);

NAND2xp33_ASAP7_75t_L g1316 ( 
.A(n_1188),
.B(n_836),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1058),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1090),
.A2(n_592),
.B(n_591),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1110),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1133),
.B(n_782),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1109),
.B(n_822),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_SL g1322 ( 
.A(n_1039),
.B(n_804),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1165),
.B(n_822),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1128),
.A2(n_837),
.B(n_804),
.Y(n_1324)
);

AOI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1092),
.A2(n_976),
.B(n_537),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1094),
.A2(n_592),
.B(n_537),
.Y(n_1326)
);

BUFx6f_ASAP7_75t_L g1327 ( 
.A(n_1149),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1110),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1189),
.A2(n_766),
.B(n_836),
.Y(n_1329)
);

AOI21xp33_ASAP7_75t_L g1330 ( 
.A1(n_1137),
.A2(n_360),
.B(n_359),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1165),
.B(n_804),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1192),
.B(n_804),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1124),
.B(n_804),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1107),
.A2(n_541),
.B(n_533),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1035),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1113),
.A2(n_1136),
.B(n_1117),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1104),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1129),
.A2(n_840),
.B(n_837),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1164),
.B(n_837),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1129),
.A2(n_541),
.B(n_533),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1170),
.A2(n_840),
.B(n_837),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1144),
.A2(n_976),
.B(n_542),
.Y(n_1342)
);

OAI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1169),
.A2(n_363),
.B(n_362),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1031),
.B(n_837),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1091),
.A2(n_840),
.B1(n_428),
.B2(n_426),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1102),
.A2(n_429),
.B(n_441),
.C(n_461),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1170),
.A2(n_840),
.B(n_766),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1145),
.A2(n_542),
.B(n_461),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1053),
.A2(n_840),
.B(n_836),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1135),
.B(n_364),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1135),
.B(n_367),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1032),
.A2(n_836),
.B(n_153),
.Y(n_1352)
);

A2O1A1Ixp33_ASAP7_75t_L g1353 ( 
.A1(n_1156),
.A2(n_375),
.B(n_370),
.C(n_378),
.Y(n_1353)
);

AOI21xp33_ASAP7_75t_L g1354 ( 
.A1(n_1041),
.A2(n_379),
.B(n_385),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1036),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1067),
.B(n_388),
.Y(n_1356)
);

BUFx8_ASAP7_75t_L g1357 ( 
.A(n_1121),
.Y(n_1357)
);

NAND2xp33_ASAP7_75t_SL g1358 ( 
.A(n_1149),
.B(n_390),
.Y(n_1358)
);

AO31x2_ASAP7_75t_L g1359 ( 
.A1(n_1126),
.A2(n_836),
.A3(n_12),
.B(n_13),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1036),
.A2(n_836),
.B(n_133),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1176),
.B(n_392),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1053),
.A2(n_1080),
.B(n_1123),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1060),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1085),
.Y(n_1364)
);

AOI21xp33_ASAP7_75t_L g1365 ( 
.A1(n_1179),
.A2(n_462),
.B(n_460),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1080),
.A2(n_458),
.B1(n_454),
.B2(n_451),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1060),
.A2(n_121),
.B(n_116),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1140),
.A2(n_11),
.A3(n_14),
.B(n_16),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1075),
.A2(n_125),
.B(n_119),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1176),
.B(n_393),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1141),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1076),
.B(n_394),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1068),
.A2(n_448),
.B(n_395),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1080),
.A2(n_120),
.B(n_122),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1066),
.A2(n_430),
.B(n_444),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1218),
.B(n_396),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1066),
.A2(n_425),
.B(n_443),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1075),
.A2(n_1105),
.B(n_1100),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1100),
.A2(n_187),
.B(n_231),
.Y(n_1379)
);

NOR2x1_ASAP7_75t_L g1380 ( 
.A(n_1082),
.B(n_445),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1080),
.A2(n_421),
.B1(n_440),
.B2(n_439),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1218),
.B(n_398),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1123),
.A2(n_201),
.B(n_134),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1154),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1076),
.B(n_403),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1182),
.B(n_407),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1104),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1142),
.A2(n_438),
.B1(n_436),
.B2(n_434),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1105),
.A2(n_1157),
.B(n_1139),
.Y(n_1389)
);

NOR2xp67_ASAP7_75t_L g1390 ( 
.A(n_1171),
.B(n_129),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1149),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1152),
.Y(n_1392)
);

A2O1A1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1233),
.A2(n_1156),
.B(n_1028),
.C(n_1185),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1371),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1251),
.B(n_1182),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1287),
.A2(n_1095),
.B1(n_1061),
.B2(n_1039),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1392),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1231),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1246),
.A2(n_1146),
.B(n_1048),
.Y(n_1399)
);

OAI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1330),
.A2(n_1050),
.B1(n_1042),
.B2(n_1028),
.C(n_1074),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1317),
.A2(n_1131),
.B1(n_1158),
.B2(n_1212),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1229),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1302),
.A2(n_1157),
.B(n_1139),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1354),
.A2(n_1150),
.B1(n_1202),
.B2(n_1033),
.Y(n_1404)
);

INVx8_ASAP7_75t_L g1405 ( 
.A(n_1231),
.Y(n_1405)
);

OAI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1268),
.A2(n_1033),
.B1(n_1104),
.B2(n_1101),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1249),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1286),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1269),
.B(n_1039),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1231),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1302),
.A2(n_1173),
.B(n_1161),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1238),
.A2(n_1173),
.B(n_1161),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1238),
.A2(n_1360),
.B(n_1352),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1249),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1253),
.Y(n_1415)
);

NOR2xp67_ASAP7_75t_L g1416 ( 
.A(n_1257),
.B(n_1180),
.Y(n_1416)
);

INVxp67_ASAP7_75t_SL g1417 ( 
.A(n_1231),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1243),
.B(n_1078),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1348),
.A2(n_1051),
.B(n_1040),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1352),
.A2(n_1201),
.B(n_1174),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1256),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1313),
.A2(n_1114),
.B1(n_1162),
.B2(n_1202),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1240),
.A2(n_1191),
.B(n_1038),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1360),
.A2(n_1174),
.B(n_1201),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_1227),
.B(n_1154),
.Y(n_1425)
);

BUFx2_ASAP7_75t_SL g1426 ( 
.A(n_1247),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1227),
.A2(n_1200),
.B(n_1196),
.Y(n_1427)
);

OAI21xp5_ASAP7_75t_L g1428 ( 
.A1(n_1291),
.A2(n_1185),
.B(n_1132),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1267),
.Y(n_1429)
);

OAI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1242),
.A2(n_1033),
.B1(n_1179),
.B2(n_1183),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1237),
.A2(n_1093),
.B(n_1042),
.C(n_1074),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1275),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1224),
.B(n_1386),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1365),
.A2(n_1114),
.B1(n_1204),
.B2(n_1130),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1297),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1278),
.B(n_1057),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1252),
.B(n_1134),
.Y(n_1437)
);

INVx8_ASAP7_75t_L g1438 ( 
.A(n_1250),
.Y(n_1438)
);

AND2x4_ASAP7_75t_L g1439 ( 
.A(n_1252),
.B(n_1134),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1234),
.B(n_1116),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_1234),
.B(n_1116),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1239),
.B(n_1160),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1314),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1378),
.A2(n_1207),
.B(n_1209),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1250),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1256),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1277),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_1257),
.Y(n_1448)
);

INVx5_ASAP7_75t_L g1449 ( 
.A(n_1250),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1308),
.Y(n_1450)
);

NAND3xp33_ASAP7_75t_L g1451 ( 
.A(n_1313),
.B(n_1222),
.C(n_1078),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1298),
.Y(n_1452)
);

INVx5_ASAP7_75t_L g1453 ( 
.A(n_1250),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1378),
.A2(n_1207),
.B(n_1209),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1298),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1389),
.A2(n_1069),
.B(n_1071),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1355),
.Y(n_1457)
);

NAND2x1p5_ASAP7_75t_L g1458 ( 
.A(n_1389),
.B(n_1166),
.Y(n_1458)
);

CKINVDCx16_ASAP7_75t_R g1459 ( 
.A(n_1247),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1301),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1276),
.B(n_1073),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1355),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_SL g1463 ( 
.A(n_1356),
.B(n_1222),
.C(n_1072),
.Y(n_1463)
);

AO31x2_ASAP7_75t_L g1464 ( 
.A1(n_1299),
.A2(n_1084),
.A3(n_1089),
.B(n_1097),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1274),
.B(n_1098),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1239),
.B(n_1160),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1363),
.Y(n_1467)
);

AO32x2_ASAP7_75t_L g1468 ( 
.A1(n_1289),
.A2(n_1220),
.A3(n_1213),
.B1(n_1221),
.B2(n_1103),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1241),
.A2(n_1119),
.B(n_1127),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1258),
.A2(n_1138),
.B(n_1184),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1343),
.B(n_1181),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1319),
.B(n_1166),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1363),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1258),
.A2(n_1177),
.B(n_1186),
.Y(n_1474)
);

AO31x2_ASAP7_75t_L g1475 ( 
.A1(n_1299),
.A2(n_1175),
.A3(n_1220),
.B(n_1213),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1326),
.A2(n_1190),
.B(n_1205),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1348),
.A2(n_1211),
.B(n_1123),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1346),
.A2(n_1148),
.B(n_1205),
.C(n_1203),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1375),
.A2(n_1221),
.B1(n_1181),
.B2(n_1148),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1315),
.Y(n_1480)
);

AOI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1228),
.A2(n_1211),
.B(n_1148),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1377),
.A2(n_1372),
.B1(n_1385),
.B2(n_1310),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1319),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1265),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1326),
.A2(n_1211),
.B(n_414),
.Y(n_1485)
);

OA21x2_ASAP7_75t_L g1486 ( 
.A1(n_1318),
.A2(n_418),
.B(n_1203),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1280),
.B(n_1190),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1340),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1303),
.A2(n_1188),
.B(n_1196),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1334),
.A2(n_1188),
.B(n_1196),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1334),
.A2(n_1188),
.B(n_1196),
.Y(n_1491)
);

OR2x6_ASAP7_75t_L g1492 ( 
.A(n_1226),
.B(n_1125),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1283),
.B(n_1166),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1281),
.B(n_1166),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1328),
.B(n_1187),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1311),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1284),
.B(n_1187),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1296),
.B(n_1187),
.Y(n_1498)
);

NAND3xp33_ASAP7_75t_L g1499 ( 
.A(n_1353),
.B(n_1187),
.C(n_1167),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1318),
.A2(n_1188),
.B(n_1125),
.Y(n_1500)
);

AO21x2_ASAP7_75t_L g1501 ( 
.A1(n_1254),
.A2(n_1188),
.B(n_445),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1244),
.A2(n_226),
.B(n_225),
.Y(n_1502)
);

AO21x2_ASAP7_75t_L g1503 ( 
.A1(n_1259),
.A2(n_218),
.B(n_217),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1279),
.A2(n_213),
.B(n_211),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1282),
.B(n_14),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1350),
.B(n_16),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1283),
.B(n_210),
.Y(n_1507)
);

NAND2x1p5_ASAP7_75t_L g1508 ( 
.A(n_1328),
.B(n_1384),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1255),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1244),
.A2(n_197),
.B(n_194),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1261),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_1255),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1367),
.A2(n_193),
.B(n_183),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1235),
.A2(n_182),
.B(n_177),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1367),
.A2(n_173),
.B(n_169),
.Y(n_1515)
);

NAND2x1p5_ASAP7_75t_L g1516 ( 
.A(n_1384),
.B(n_168),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1255),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1307),
.Y(n_1518)
);

A2O1A1Ixp33_ASAP7_75t_SL g1519 ( 
.A1(n_1329),
.A2(n_1230),
.B(n_1373),
.C(n_1347),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1369),
.A2(n_166),
.B(n_160),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1262),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1255),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1337),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1305),
.Y(n_1524)
);

AO21x2_ASAP7_75t_L g1525 ( 
.A1(n_1294),
.A2(n_158),
.B(n_149),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1288),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1266),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1305),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1331),
.Y(n_1529)
);

OAI21xp5_ASAP7_75t_L g1530 ( 
.A1(n_1272),
.A2(n_17),
.B(n_18),
.Y(n_1530)
);

AO21x2_ASAP7_75t_L g1531 ( 
.A1(n_1294),
.A2(n_17),
.B(n_19),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1293),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1332),
.B(n_1333),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1380),
.A2(n_1062),
.B1(n_22),
.B2(n_24),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1320),
.B(n_20),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1285),
.A2(n_25),
.B(n_28),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1391),
.B(n_25),
.Y(n_1537)
);

INVx3_ASAP7_75t_L g1538 ( 
.A(n_1288),
.Y(n_1538)
);

INVx1_ASAP7_75t_SL g1539 ( 
.A(n_1265),
.Y(n_1539)
);

OAI211xp5_ASAP7_75t_L g1540 ( 
.A1(n_1351),
.A2(n_28),
.B(n_30),
.C(n_32),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_SL g1541 ( 
.A1(n_1383),
.A2(n_30),
.B(n_35),
.Y(n_1541)
);

AO21x2_ASAP7_75t_L g1542 ( 
.A1(n_1336),
.A2(n_1325),
.B(n_1342),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1369),
.A2(n_35),
.B(n_37),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1379),
.A2(n_38),
.B(n_39),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1288),
.Y(n_1545)
);

INVx2_ASAP7_75t_SL g1546 ( 
.A(n_1226),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1305),
.Y(n_1547)
);

O2A1O1Ixp33_ASAP7_75t_SL g1548 ( 
.A1(n_1346),
.A2(n_38),
.B(n_42),
.C(n_44),
.Y(n_1548)
);

NAND2x1p5_ASAP7_75t_L g1549 ( 
.A(n_1379),
.B(n_45),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1306),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1248),
.A2(n_45),
.B(n_48),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1305),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1323),
.B(n_48),
.Y(n_1553)
);

AO21x2_ASAP7_75t_L g1554 ( 
.A1(n_1336),
.A2(n_51),
.B(n_52),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1236),
.Y(n_1555)
);

OAI21x1_ASAP7_75t_L g1556 ( 
.A1(n_1263),
.A2(n_52),
.B(n_53),
.Y(n_1556)
);

OR2x6_ASAP7_75t_L g1557 ( 
.A(n_1335),
.B(n_53),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1288),
.Y(n_1558)
);

OAI221xp5_ASAP7_75t_L g1559 ( 
.A1(n_1361),
.A2(n_56),
.B1(n_58),
.B2(n_67),
.C(n_68),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1290),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1376),
.B(n_103),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1232),
.A2(n_1341),
.B(n_1285),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1358),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_SL g1564 ( 
.A1(n_1245),
.A2(n_69),
.B(n_70),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1364),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1339),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1300),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_L g1568 ( 
.A(n_1300),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1290),
.Y(n_1569)
);

AOI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1390),
.A2(n_71),
.B1(n_72),
.B2(n_76),
.Y(n_1570)
);

INVx4_ASAP7_75t_L g1571 ( 
.A(n_1300),
.Y(n_1571)
);

OA21x2_ASAP7_75t_L g1572 ( 
.A1(n_1263),
.A2(n_71),
.B(n_76),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1391),
.B(n_77),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1290),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1382),
.Y(n_1575)
);

OAI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1570),
.A2(n_1387),
.B1(n_1271),
.B2(n_1236),
.Y(n_1576)
);

OAI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1418),
.A2(n_1404),
.B1(n_1479),
.B2(n_1482),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1394),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1559),
.A2(n_1358),
.B1(n_1388),
.B2(n_1271),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1395),
.A2(n_1335),
.B1(n_1370),
.B2(n_1353),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1397),
.Y(n_1581)
);

INVx5_ASAP7_75t_L g1582 ( 
.A(n_1557),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1434),
.A2(n_1335),
.B1(n_1364),
.B2(n_1321),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1506),
.A2(n_1381),
.B1(n_1366),
.B2(n_1345),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1433),
.B(n_1225),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1402),
.Y(n_1586)
);

AOI21xp33_ASAP7_75t_L g1587 ( 
.A1(n_1519),
.A2(n_1451),
.B(n_1400),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1536),
.A2(n_1357),
.B1(n_1225),
.B2(n_1374),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1511),
.B(n_1357),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1433),
.B(n_1368),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1447),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1415),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1448),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1563),
.A2(n_1357),
.B1(n_1344),
.B2(n_1322),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1521),
.B(n_1327),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1429),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1432),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1575),
.B(n_1368),
.Y(n_1598)
);

NAND3xp33_ASAP7_75t_SL g1599 ( 
.A(n_1534),
.B(n_1292),
.C(n_1362),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1435),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1530),
.A2(n_1304),
.B1(n_1270),
.B2(n_1316),
.Y(n_1601)
);

AOI221xp5_ASAP7_75t_L g1602 ( 
.A1(n_1430),
.A2(n_1309),
.B1(n_1312),
.B2(n_1304),
.C(n_1316),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1443),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1527),
.B(n_1300),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1422),
.A2(n_1327),
.B1(n_1368),
.B2(n_1338),
.Y(n_1605)
);

NAND2x1_ASAP7_75t_L g1606 ( 
.A(n_1409),
.B(n_1483),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1460),
.A2(n_1327),
.B1(n_1273),
.B2(n_1264),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1398),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1535),
.B(n_1368),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1407),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1461),
.B(n_1327),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1514),
.A2(n_1324),
.B1(n_1295),
.B2(n_1359),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1408),
.B(n_1359),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1436),
.B(n_1359),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1405),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1519),
.A2(n_1260),
.B(n_1273),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1465),
.B(n_1359),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1465),
.B(n_1290),
.Y(n_1618)
);

CKINVDCx20_ASAP7_75t_R g1619 ( 
.A(n_1448),
.Y(n_1619)
);

AOI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1561),
.A2(n_1349),
.B1(n_83),
.B2(n_84),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1413),
.A2(n_79),
.B(n_83),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1452),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_SL g1623 ( 
.A1(n_1393),
.A2(n_79),
.B(n_89),
.C(n_90),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1457),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1535),
.B(n_1487),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1487),
.B(n_90),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1428),
.A2(n_102),
.B1(n_93),
.B2(n_100),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1478),
.A2(n_93),
.B(n_101),
.Y(n_1628)
);

INVx1_ASAP7_75t_SL g1629 ( 
.A(n_1450),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1463),
.A2(n_101),
.B1(n_102),
.B2(n_1557),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1414),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1529),
.B(n_1497),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1523),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1414),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1535),
.B(n_1497),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_SL g1636 ( 
.A(n_1393),
.B(n_1540),
.C(n_1431),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1557),
.A2(n_1406),
.B1(n_1499),
.B2(n_1553),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1498),
.A2(n_1423),
.B(n_1427),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1426),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1505),
.B(n_1553),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1557),
.A2(n_1541),
.B1(n_1533),
.B2(n_1503),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1533),
.B(n_1431),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1550),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1644)
);

CKINVDCx6p67_ASAP7_75t_R g1645 ( 
.A(n_1555),
.Y(n_1645)
);

BUFx10_ASAP7_75t_L g1646 ( 
.A(n_1532),
.Y(n_1646)
);

O2A1O1Ixp33_ASAP7_75t_SL g1647 ( 
.A1(n_1498),
.A2(n_1566),
.B(n_1494),
.C(n_1504),
.Y(n_1647)
);

INVxp67_ASAP7_75t_SL g1648 ( 
.A(n_1483),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1526),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1467),
.Y(n_1651)
);

OAI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1401),
.A2(n_1471),
.B1(n_1492),
.B2(n_1396),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1541),
.A2(n_1503),
.B1(n_1531),
.B2(n_1554),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1493),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1421),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1446),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1437),
.B(n_1439),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1446),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1455),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1455),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1413),
.A2(n_1412),
.B(n_1556),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_SL g1662 ( 
.A1(n_1537),
.A2(n_1573),
.B1(n_1555),
.B2(n_1503),
.Y(n_1662)
);

CKINVDCx8_ASAP7_75t_R g1663 ( 
.A(n_1459),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1462),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1565),
.A2(n_1416),
.B1(n_1440),
.B2(n_1441),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1484),
.B(n_1539),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1442),
.B(n_1466),
.Y(n_1667)
);

AOI221xp5_ASAP7_75t_L g1668 ( 
.A1(n_1548),
.A2(n_1564),
.B1(n_1440),
.B2(n_1441),
.C(n_1565),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1442),
.B(n_1466),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1440),
.A2(n_1532),
.B1(n_1492),
.B2(n_1409),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_L g1671 ( 
.A1(n_1420),
.A2(n_1424),
.B(n_1491),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1507),
.Y(n_1672)
);

OAI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1492),
.A2(n_1409),
.B1(n_1516),
.B2(n_1425),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1405),
.Y(n_1674)
);

INVx6_ASAP7_75t_L g1675 ( 
.A(n_1405),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1473),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1507),
.B(n_1442),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1507),
.B(n_1466),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1538),
.B(n_1545),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1526),
.B(n_1546),
.Y(n_1680)
);

AOI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1564),
.A2(n_1501),
.B1(n_1531),
.B2(n_1554),
.C(n_1574),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1464),
.Y(n_1682)
);

AOI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1481),
.A2(n_1488),
.B(n_1552),
.Y(n_1683)
);

BUFx8_ASAP7_75t_SL g1684 ( 
.A(n_1410),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1546),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1417),
.B(n_1538),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1409),
.A2(n_1508),
.B1(n_1549),
.B2(n_1572),
.Y(n_1687)
);

BUFx2_ASAP7_75t_L g1688 ( 
.A(n_1538),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1545),
.B(n_1464),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1545),
.B(n_1464),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1444),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1464),
.B(n_1475),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1464),
.Y(n_1693)
);

INVx4_ASAP7_75t_L g1694 ( 
.A(n_1405),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1456),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1501),
.A2(n_1562),
.B(n_1399),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1410),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1438),
.Y(n_1698)
);

NAND3xp33_ASAP7_75t_L g1699 ( 
.A(n_1485),
.B(n_1486),
.C(n_1572),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1438),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1475),
.B(n_1398),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1398),
.B(n_1445),
.Y(n_1702)
);

BUFx2_ASAP7_75t_SL g1703 ( 
.A(n_1449),
.Y(n_1703)
);

AOI22xp33_ASAP7_75t_L g1704 ( 
.A1(n_1531),
.A2(n_1554),
.B1(n_1501),
.B2(n_1399),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1456),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1475),
.B(n_1522),
.Y(n_1706)
);

AOI222xp33_ASAP7_75t_L g1707 ( 
.A1(n_1551),
.A2(n_1524),
.B1(n_1528),
.B2(n_1547),
.C1(n_1552),
.C2(n_1574),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1475),
.B(n_1517),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1438),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1425),
.A2(n_1483),
.B1(n_1399),
.B2(n_1562),
.Y(n_1710)
);

NAND3xp33_ASAP7_75t_L g1711 ( 
.A(n_1485),
.B(n_1486),
.C(n_1572),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1551),
.A2(n_1560),
.B1(n_1569),
.B2(n_1525),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1562),
.A2(n_1508),
.B1(n_1517),
.B2(n_1571),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1560),
.A2(n_1569),
.B1(n_1525),
.B2(n_1419),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1438),
.Y(n_1715)
);

INVx5_ASAP7_75t_L g1716 ( 
.A(n_1449),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1475),
.B(n_1571),
.Y(n_1717)
);

OA21x2_ASAP7_75t_L g1718 ( 
.A1(n_1412),
.A2(n_1556),
.B(n_1469),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1449),
.B(n_1453),
.Y(n_1719)
);

CKINVDCx20_ASAP7_75t_R g1720 ( 
.A(n_1445),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1410),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1410),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1509),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1449),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1525),
.A2(n_1419),
.B1(n_1549),
.B2(n_1544),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1449),
.B(n_1453),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1453),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1509),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_1453),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1509),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1509),
.Y(n_1731)
);

AOI21xp33_ASAP7_75t_L g1732 ( 
.A1(n_1419),
.A2(n_1485),
.B(n_1477),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1549),
.A2(n_1480),
.B1(n_1496),
.B2(n_1518),
.C(n_1542),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1454),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1453),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1512),
.Y(n_1736)
);

BUFx4_ASAP7_75t_SL g1737 ( 
.A(n_1445),
.Y(n_1737)
);

BUFx6f_ASAP7_75t_L g1738 ( 
.A(n_1512),
.Y(n_1738)
);

AOI222xp33_ASAP7_75t_L g1739 ( 
.A1(n_1543),
.A2(n_1544),
.B1(n_1571),
.B2(n_1517),
.C1(n_1522),
.C2(n_1558),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1512),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1512),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_R g1742 ( 
.A(n_1512),
.B(n_1568),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1480),
.A2(n_1496),
.B1(n_1518),
.B2(n_1542),
.C(n_1522),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1500),
.B(n_1489),
.Y(n_1744)
);

INVx4_ASAP7_75t_SL g1745 ( 
.A(n_1558),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1472),
.A2(n_1495),
.B1(n_1567),
.B2(n_1558),
.Y(n_1746)
);

NOR2xp67_ASAP7_75t_SL g1747 ( 
.A(n_1558),
.B(n_1568),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1568),
.B(n_1567),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1495),
.A2(n_1458),
.B1(n_1567),
.B2(n_1558),
.Y(n_1749)
);

INVx6_ASAP7_75t_L g1750 ( 
.A(n_1567),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1567),
.B(n_1568),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1568),
.B(n_1477),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_1477),
.B(n_1458),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1500),
.B(n_1470),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1543),
.B(n_1486),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1458),
.Y(n_1756)
);

NAND2x1p5_ASAP7_75t_L g1757 ( 
.A(n_1489),
.B(n_1490),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1474),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1513),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1502),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1474),
.B(n_1468),
.Y(n_1761)
);

INVx4_ASAP7_75t_L g1762 ( 
.A(n_1542),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1502),
.A2(n_1510),
.B1(n_1515),
.B2(n_1513),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_1510),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1403),
.B(n_1411),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_1636),
.Y(n_1766)
);

BUFx4f_ASAP7_75t_SL g1767 ( 
.A(n_1619),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1585),
.B(n_1520),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1613),
.B(n_1403),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1627),
.A2(n_1520),
.B1(n_1515),
.B2(n_1411),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1584),
.A2(n_1468),
.B1(n_1490),
.B2(n_1491),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1720),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1619),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_L g1774 ( 
.A1(n_1630),
.A2(n_1468),
.B1(n_1476),
.B2(n_1420),
.C(n_1424),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1635),
.B(n_1468),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1579),
.B(n_1468),
.C(n_1476),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1640),
.A2(n_1588),
.B1(n_1628),
.B2(n_1620),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1640),
.A2(n_1620),
.B1(n_1579),
.B2(n_1587),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1637),
.A2(n_1594),
.B1(n_1576),
.B2(n_1642),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1623),
.A2(n_1637),
.B(n_1594),
.C(n_1668),
.Y(n_1780)
);

OAI22xp33_ASAP7_75t_L g1781 ( 
.A1(n_1582),
.A2(n_1665),
.B1(n_1670),
.B2(n_1652),
.Y(n_1781)
);

OAI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1623),
.A2(n_1605),
.B(n_1626),
.C(n_1662),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1582),
.A2(n_1589),
.B1(n_1583),
.B2(n_1639),
.Y(n_1783)
);

INVx5_ASAP7_75t_L g1784 ( 
.A(n_1716),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_SL g1785 ( 
.A1(n_1582),
.A2(n_1580),
.B1(n_1672),
.B2(n_1687),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1638),
.A2(n_1647),
.B(n_1673),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1666),
.A2(n_1599),
.B1(n_1677),
.B2(n_1678),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1653),
.A2(n_1641),
.B(n_1605),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1625),
.B(n_1644),
.Y(n_1789)
);

HB1xp67_ASAP7_75t_L g1790 ( 
.A(n_1591),
.Y(n_1790)
);

INVx1_ASAP7_75t_SL g1791 ( 
.A(n_1629),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1632),
.B(n_1611),
.Y(n_1792)
);

CKINVDCx16_ASAP7_75t_R g1793 ( 
.A(n_1646),
.Y(n_1793)
);

AOI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1590),
.A2(n_1598),
.B1(n_1643),
.B2(n_1581),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1586),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1667),
.B(n_1669),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1592),
.A2(n_1600),
.B1(n_1603),
.B2(n_1597),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1641),
.A2(n_1653),
.B1(n_1612),
.B2(n_1647),
.C(n_1633),
.Y(n_1798)
);

AOI22xp33_ASAP7_75t_L g1799 ( 
.A1(n_1596),
.A2(n_1602),
.B1(n_1609),
.B2(n_1614),
.Y(n_1799)
);

AOI222xp33_ASAP7_75t_L g1800 ( 
.A1(n_1677),
.A2(n_1678),
.B1(n_1657),
.B2(n_1650),
.C1(n_1617),
.C2(n_1618),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1645),
.A2(n_1663),
.B1(n_1593),
.B2(n_1672),
.Y(n_1801)
);

AOI22x1_ASAP7_75t_L g1802 ( 
.A1(n_1760),
.A2(n_1764),
.B1(n_1593),
.B2(n_1739),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1677),
.A2(n_1678),
.B1(n_1650),
.B2(n_1657),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_SL g1804 ( 
.A1(n_1704),
.A2(n_1681),
.B1(n_1612),
.B2(n_1725),
.C(n_1763),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1622),
.Y(n_1805)
);

OAI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1645),
.A2(n_1672),
.B1(n_1606),
.B2(n_1720),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1616),
.A2(n_1607),
.B(n_1601),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1709),
.A2(n_1715),
.B1(n_1601),
.B2(n_1650),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1624),
.Y(n_1809)
);

A2O1A1Ixp33_ASAP7_75t_L g1810 ( 
.A1(n_1760),
.A2(n_1764),
.B(n_1710),
.C(n_1704),
.Y(n_1810)
);

OAI22xp5_ASAP7_75t_L g1811 ( 
.A1(n_1709),
.A2(n_1715),
.B1(n_1657),
.B2(n_1685),
.Y(n_1811)
);

AOI222xp33_ASAP7_75t_L g1812 ( 
.A1(n_1651),
.A2(n_1692),
.B1(n_1595),
.B2(n_1604),
.C1(n_1690),
.C2(n_1689),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1659),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1664),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1646),
.A2(n_1621),
.B1(n_1649),
.B2(n_1654),
.Y(n_1815)
);

A2O1A1Ixp33_ASAP7_75t_L g1816 ( 
.A1(n_1696),
.A2(n_1713),
.B(n_1621),
.C(n_1725),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1682),
.A2(n_1693),
.B1(n_1732),
.B2(n_1733),
.C(n_1753),
.Y(n_1817)
);

CKINVDCx11_ASAP7_75t_R g1818 ( 
.A(n_1615),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1676),
.B(n_1748),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1654),
.A2(n_1634),
.B1(n_1610),
.B2(n_1660),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1680),
.B(n_1686),
.Y(n_1821)
);

AOI22xp33_ASAP7_75t_SL g1822 ( 
.A1(n_1742),
.A2(n_1703),
.B1(n_1716),
.B2(n_1740),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1679),
.B(n_1610),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1631),
.A2(n_1658),
.B1(n_1656),
.B2(n_1634),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1746),
.A2(n_1711),
.B1(n_1699),
.B2(n_1743),
.C(n_1712),
.Y(n_1825)
);

AOI221x1_ASAP7_75t_L g1826 ( 
.A1(n_1752),
.A2(n_1749),
.B1(n_1753),
.B2(n_1706),
.C(n_1701),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1712),
.A2(n_1752),
.B1(n_1708),
.B2(n_1717),
.C(n_1705),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1679),
.B(n_1688),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1655),
.B(n_1656),
.Y(n_1829)
);

OAI222xp33_ASAP7_75t_L g1830 ( 
.A1(n_1747),
.A2(n_1719),
.B1(n_1648),
.B2(n_1726),
.C1(n_1727),
.C2(n_1694),
.Y(n_1830)
);

NAND2xp33_ASAP7_75t_SL g1831 ( 
.A(n_1742),
.B(n_1615),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_SL g1832 ( 
.A1(n_1716),
.A2(n_1724),
.B1(n_1735),
.B2(n_1727),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1679),
.A2(n_1759),
.B1(n_1707),
.B2(n_1675),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1751),
.B(n_1697),
.Y(n_1834)
);

AO221x2_ASAP7_75t_L g1835 ( 
.A1(n_1695),
.A2(n_1721),
.B1(n_1741),
.B2(n_1723),
.C(n_1730),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1751),
.B(n_1731),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1759),
.A2(n_1675),
.B1(n_1700),
.B2(n_1694),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1722),
.B(n_1728),
.Y(n_1838)
);

OAI21x1_ASAP7_75t_L g1839 ( 
.A1(n_1671),
.A2(n_1765),
.B(n_1757),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1675),
.A2(n_1716),
.B1(n_1700),
.B2(n_1694),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1759),
.A2(n_1674),
.B1(n_1755),
.B2(n_1702),
.Y(n_1841)
);

AOI221xp5_ASAP7_75t_L g1842 ( 
.A1(n_1714),
.A2(n_1758),
.B1(n_1761),
.B2(n_1759),
.C(n_1762),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1674),
.A2(n_1702),
.B1(n_1615),
.B2(n_1698),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1702),
.B(n_1736),
.Y(n_1844)
);

AOI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1674),
.A2(n_1608),
.B1(n_1719),
.B2(n_1615),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1684),
.Y(n_1846)
);

OAI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1727),
.A2(n_1735),
.B1(n_1724),
.B2(n_1726),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1608),
.A2(n_1684),
.B1(n_1762),
.B2(n_1750),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_L g1849 ( 
.A1(n_1762),
.A2(n_1714),
.B(n_1718),
.Y(n_1849)
);

OAI211xp5_ASAP7_75t_SL g1850 ( 
.A1(n_1756),
.A2(n_1729),
.B(n_1691),
.C(n_1734),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1729),
.A2(n_1756),
.B1(n_1750),
.B2(n_1738),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1729),
.A2(n_1738),
.B1(n_1744),
.B2(n_1754),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1744),
.A2(n_1757),
.B(n_1754),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1734),
.A2(n_1738),
.B1(n_1754),
.B2(n_1718),
.Y(n_1854)
);

AOI22xp33_ASAP7_75t_L g1855 ( 
.A1(n_1738),
.A2(n_1718),
.B1(n_1745),
.B2(n_1661),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1737),
.A2(n_658),
.B1(n_1354),
.B2(n_891),
.C(n_870),
.Y(n_1856)
);

OAI211xp5_ASAP7_75t_L g1857 ( 
.A1(n_1661),
.A2(n_1627),
.B(n_1041),
.C(n_1630),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1745),
.A2(n_1627),
.B1(n_1577),
.B2(n_1630),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1744),
.B(n_1661),
.Y(n_1859)
);

INVxp33_ASAP7_75t_L g1860 ( 
.A(n_1666),
.Y(n_1860)
);

OAI221xp5_ASAP7_75t_L g1861 ( 
.A1(n_1630),
.A2(n_1041),
.B1(n_1045),
.B2(n_716),
.C(n_866),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1591),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1627),
.A2(n_658),
.B1(n_1354),
.B2(n_891),
.C(n_870),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1585),
.B(n_1635),
.Y(n_1865)
);

BUFx4f_ASAP7_75t_SL g1866 ( 
.A(n_1619),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1867)
);

NAND4xp25_ASAP7_75t_L g1868 ( 
.A(n_1640),
.B(n_658),
.C(n_891),
.D(n_1354),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1577),
.A2(n_1045),
.B(n_716),
.C(n_866),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_1404),
.B2(n_866),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1613),
.B(n_1590),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1873)
);

OAI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1630),
.A2(n_1041),
.B1(n_1045),
.B2(n_716),
.C(n_866),
.Y(n_1874)
);

AOI221xp5_ASAP7_75t_L g1875 ( 
.A1(n_1627),
.A2(n_658),
.B1(n_1354),
.B2(n_891),
.C(n_870),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1578),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_973),
.B2(n_872),
.Y(n_1877)
);

OAI21x1_ASAP7_75t_L g1878 ( 
.A1(n_1683),
.A2(n_1413),
.B(n_1671),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1879)
);

OAI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_973),
.B2(n_872),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1577),
.B(n_870),
.C(n_716),
.Y(n_1881)
);

OAI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_1404),
.B2(n_866),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1613),
.B(n_1590),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1884)
);

AOI21xp33_ASAP7_75t_L g1885 ( 
.A1(n_1577),
.A2(n_716),
.B(n_1159),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1886)
);

AOI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1627),
.A2(n_658),
.B1(n_1354),
.B2(n_891),
.C(n_870),
.Y(n_1887)
);

A2O1A1Ixp33_ASAP7_75t_L g1888 ( 
.A1(n_1584),
.A2(n_1041),
.B(n_1159),
.C(n_1451),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1889)
);

AOI22xp33_ASAP7_75t_L g1890 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_1404),
.B2(n_866),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1577),
.A2(n_866),
.B1(n_973),
.B2(n_872),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1578),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_L g1894 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1895)
);

OAI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_973),
.B2(n_872),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1897)
);

AOI221xp5_ASAP7_75t_L g1898 ( 
.A1(n_1627),
.A2(n_658),
.B1(n_1354),
.B2(n_891),
.C(n_870),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1587),
.A2(n_1041),
.B(n_1354),
.C(n_691),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1578),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1578),
.Y(n_1901)
);

AOI222xp33_ASAP7_75t_L g1902 ( 
.A1(n_1627),
.A2(n_626),
.B1(n_866),
.B2(n_1577),
.C1(n_1045),
.C2(n_1506),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1613),
.B(n_1590),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1578),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1907)
);

OAI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1584),
.A2(n_1041),
.B1(n_973),
.B2(n_872),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1909)
);

INVx4_ASAP7_75t_SL g1910 ( 
.A(n_1675),
.Y(n_1910)
);

AOI22xp33_ASAP7_75t_L g1911 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1911)
);

AOI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1577),
.A2(n_1045),
.B1(n_866),
.B2(n_1041),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_SL g1913 ( 
.A1(n_1577),
.A2(n_866),
.B1(n_973),
.B2(n_872),
.Y(n_1913)
);

AOI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1627),
.A2(n_658),
.B1(n_1354),
.B2(n_891),
.C(n_870),
.Y(n_1914)
);

BUFx6f_ASAP7_75t_L g1915 ( 
.A(n_1615),
.Y(n_1915)
);

OR2x6_ASAP7_75t_L g1916 ( 
.A(n_1606),
.B(n_1687),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1578),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1640),
.B(n_1632),
.Y(n_1919)
);

OAI21xp33_ASAP7_75t_L g1920 ( 
.A1(n_1627),
.A2(n_870),
.B(n_716),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1627),
.A2(n_1577),
.B1(n_1630),
.B2(n_658),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1638),
.A2(n_1519),
.B(n_1514),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1684),
.Y(n_1923)
);

AOI222xp33_ASAP7_75t_L g1924 ( 
.A1(n_1627),
.A2(n_626),
.B1(n_866),
.B2(n_1577),
.C1(n_1045),
.C2(n_1506),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1578),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_L g1926 ( 
.A(n_1577),
.B(n_870),
.C(n_716),
.Y(n_1926)
);

NOR2x1_ASAP7_75t_L g1927 ( 
.A(n_1830),
.B(n_1850),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_1839),
.Y(n_1928)
);

HB1xp67_ASAP7_75t_L g1929 ( 
.A(n_1835),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1835),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1871),
.B(n_1883),
.Y(n_1931)
);

OAI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1766),
.A2(n_1905),
.B1(n_1886),
.B2(n_1884),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1805),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1903),
.B(n_1769),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1859),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1853),
.B(n_1916),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1878),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1916),
.B(n_1826),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1799),
.B(n_1812),
.Y(n_1939)
);

AOI22xp33_ASAP7_75t_SL g1940 ( 
.A1(n_1861),
.A2(n_1874),
.B1(n_1870),
.B2(n_1891),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1809),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1835),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1790),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1775),
.B(n_1768),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1916),
.B(n_1854),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1854),
.B(n_1841),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1799),
.B(n_1862),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1827),
.B(n_1865),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1795),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1893),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1900),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1901),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1852),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1904),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1863),
.Y(n_1955)
);

HB1xp67_ASAP7_75t_L g1956 ( 
.A(n_1819),
.Y(n_1956)
);

NAND2x1p5_ASAP7_75t_L g1957 ( 
.A(n_1784),
.B(n_1786),
.Y(n_1957)
);

OR2x6_ASAP7_75t_L g1958 ( 
.A(n_1807),
.B(n_1922),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_SL g1959 ( 
.A1(n_1882),
.A2(n_1857),
.B1(n_1926),
.B2(n_1881),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1917),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_SL g1961 ( 
.A1(n_1780),
.A2(n_1902),
.B1(n_1924),
.B2(n_1782),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1925),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1772),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1813),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1814),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_SL g1966 ( 
.A1(n_1802),
.A2(n_1766),
.B1(n_1783),
.B2(n_1921),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1873),
.B(n_1889),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1876),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1829),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1823),
.Y(n_1970)
);

OA21x2_ASAP7_75t_L g1971 ( 
.A1(n_1816),
.A2(n_1849),
.B(n_1817),
.Y(n_1971)
);

BUFx2_ASAP7_75t_L g1972 ( 
.A(n_1810),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1825),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1774),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1797),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1771),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1794),
.B(n_1788),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1797),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1776),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_L g1980 ( 
.A1(n_1867),
.A2(n_1906),
.B1(n_1921),
.B2(n_1872),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1834),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1897),
.B(n_1919),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1789),
.B(n_1842),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1800),
.B(n_1821),
.Y(n_1984)
);

BUFx3_ASAP7_75t_L g1985 ( 
.A(n_1784),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1836),
.Y(n_1986)
);

OAI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1864),
.A2(n_1898),
.B(n_1875),
.Y(n_1987)
);

INVx2_ASAP7_75t_L g1988 ( 
.A(n_1838),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1804),
.B(n_1792),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1787),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1778),
.B(n_1798),
.Y(n_1991)
);

HB1xp67_ASAP7_75t_L g1992 ( 
.A(n_1828),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1778),
.B(n_1888),
.Y(n_1993)
);

HB1xp67_ASAP7_75t_L g1994 ( 
.A(n_1791),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1777),
.B(n_1824),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1777),
.B(n_1824),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1844),
.Y(n_1997)
);

A2O1A1Ixp33_ASAP7_75t_L g1998 ( 
.A1(n_1920),
.A2(n_1869),
.B(n_1914),
.C(n_1887),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1808),
.Y(n_1999)
);

AOI22xp33_ASAP7_75t_L g2000 ( 
.A1(n_1867),
.A2(n_1884),
.B1(n_1918),
.B2(n_1894),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1855),
.B(n_1803),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1820),
.B(n_1855),
.Y(n_2002)
);

AOI221xp5_ASAP7_75t_L g2003 ( 
.A1(n_1872),
.A2(n_1907),
.B1(n_1906),
.B2(n_1905),
.C(n_1909),
.Y(n_2003)
);

OR2x2_ASAP7_75t_L g2004 ( 
.A(n_1815),
.B(n_1833),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1820),
.B(n_1833),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1785),
.B(n_1860),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1851),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1848),
.B(n_1781),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1847),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1848),
.B(n_1779),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1845),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1779),
.B(n_1796),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1837),
.B(n_1858),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1770),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1910),
.B(n_1915),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1793),
.B(n_1811),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1770),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1840),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1858),
.B(n_1923),
.Y(n_2019)
);

INVxp67_ASAP7_75t_L g2020 ( 
.A(n_1943),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1981),
.B(n_1912),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1944),
.B(n_1832),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1987),
.A2(n_1918),
.B1(n_1911),
.B2(n_1909),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1949),
.Y(n_2024)
);

INVx5_ASAP7_75t_L g2025 ( 
.A(n_1958),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_1987),
.A2(n_1907),
.B1(n_1890),
.B2(n_1911),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1934),
.B(n_1806),
.Y(n_2027)
);

AND2x4_ASAP7_75t_L g2028 ( 
.A(n_1936),
.B(n_1910),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1961),
.A2(n_1879),
.B1(n_1886),
.B2(n_1890),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1981),
.B(n_1885),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1994),
.Y(n_2031)
);

OAI33xp33_ASAP7_75t_L g2032 ( 
.A1(n_1932),
.A2(n_1868),
.A3(n_1896),
.B1(n_1880),
.B2(n_1908),
.B3(n_1877),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1961),
.A2(n_1940),
.B1(n_1932),
.B2(n_2003),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1951),
.Y(n_2034)
);

OAI31xp33_ASAP7_75t_L g2035 ( 
.A1(n_1998),
.A2(n_1899),
.A3(n_1894),
.B(n_1879),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1951),
.Y(n_2036)
);

OAI221xp5_ASAP7_75t_L g2037 ( 
.A1(n_1940),
.A2(n_1913),
.B1(n_1892),
.B2(n_1856),
.C(n_1895),
.Y(n_2037)
);

NOR2xp33_ASAP7_75t_L g2038 ( 
.A(n_1967),
.B(n_1982),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1944),
.B(n_1843),
.Y(n_2039)
);

AOI22xp33_ASAP7_75t_L g2040 ( 
.A1(n_2003),
.A2(n_1972),
.B1(n_1980),
.B2(n_2000),
.Y(n_2040)
);

OR2x6_ASAP7_75t_L g2041 ( 
.A(n_1958),
.B(n_1915),
.Y(n_2041)
);

OAI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1972),
.A2(n_1801),
.B1(n_1767),
.B2(n_1866),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1936),
.B(n_1846),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1935),
.B(n_1843),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1967),
.B(n_1982),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_1943),
.Y(n_2046)
);

AOI22xp5_ASAP7_75t_L g2047 ( 
.A1(n_1959),
.A2(n_1895),
.B1(n_1773),
.B2(n_1831),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1960),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1960),
.Y(n_2049)
);

AND2x6_ASAP7_75t_SL g2050 ( 
.A(n_1993),
.B(n_1767),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1959),
.A2(n_1866),
.B1(n_1818),
.B2(n_1822),
.Y(n_2051)
);

AOI21x1_ASAP7_75t_L g2052 ( 
.A1(n_1973),
.A2(n_1958),
.B(n_1993),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1935),
.B(n_1988),
.Y(n_2053)
);

BUFx6f_ASAP7_75t_L g2054 ( 
.A(n_1985),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1963),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1955),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_1934),
.B(n_1976),
.Y(n_2057)
);

AO21x2_ASAP7_75t_L g2058 ( 
.A1(n_1937),
.A2(n_1979),
.B(n_2014),
.Y(n_2058)
);

BUFx4f_ASAP7_75t_SL g2059 ( 
.A(n_1963),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_1976),
.B(n_1931),
.Y(n_2060)
);

AOI33xp33_ASAP7_75t_L g2061 ( 
.A1(n_1966),
.A2(n_1979),
.A3(n_1977),
.B1(n_2014),
.B2(n_2017),
.B3(n_1974),
.Y(n_2061)
);

OR2x6_ASAP7_75t_L g2062 ( 
.A(n_1958),
.B(n_1957),
.Y(n_2062)
);

NOR2xp33_ASAP7_75t_L g2063 ( 
.A(n_1963),
.B(n_1973),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_1988),
.B(n_1969),
.Y(n_2064)
);

OAI211xp5_ASAP7_75t_SL g2065 ( 
.A1(n_1966),
.A2(n_1939),
.B(n_1991),
.C(n_1989),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_1955),
.B(n_1969),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1964),
.Y(n_2067)
);

OAI221xp5_ASAP7_75t_L g2068 ( 
.A1(n_1958),
.A2(n_1939),
.B1(n_1991),
.B2(n_1947),
.C(n_1989),
.Y(n_2068)
);

AOI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_2010),
.A2(n_1990),
.B1(n_1947),
.B2(n_1938),
.Y(n_2069)
);

AOI221xp5_ASAP7_75t_L g2070 ( 
.A1(n_1977),
.A2(n_2017),
.B1(n_1996),
.B2(n_1995),
.C(n_1999),
.Y(n_2070)
);

BUFx2_ASAP7_75t_L g2071 ( 
.A(n_1936),
.Y(n_2071)
);

OAI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_1995),
.A2(n_1996),
.B1(n_1999),
.B2(n_1990),
.C(n_1971),
.Y(n_2072)
);

BUFx2_ASAP7_75t_L g2073 ( 
.A(n_1929),
.Y(n_2073)
);

AOI31xp33_ASAP7_75t_L g2074 ( 
.A1(n_2016),
.A2(n_1938),
.A3(n_2004),
.B(n_2006),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1990),
.A2(n_2010),
.B1(n_1938),
.B2(n_2006),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1938),
.A2(n_2013),
.B1(n_1984),
.B2(n_2009),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1968),
.Y(n_2077)
);

AOI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2013),
.A2(n_1984),
.B1(n_2009),
.B2(n_2008),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1969),
.B(n_1981),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1986),
.B(n_2002),
.Y(n_2080)
);

INVxp67_ASAP7_75t_L g2081 ( 
.A(n_1992),
.Y(n_2081)
);

AOI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_1974),
.A2(n_1978),
.B1(n_1975),
.B2(n_2012),
.C(n_1948),
.Y(n_2082)
);

NAND4xp25_ASAP7_75t_L g2083 ( 
.A(n_1975),
.B(n_1978),
.C(n_2011),
.D(n_2019),
.Y(n_2083)
);

OAI33xp33_ASAP7_75t_L g2084 ( 
.A1(n_1933),
.A2(n_1950),
.A3(n_1941),
.B1(n_1962),
.B2(n_1954),
.B3(n_1952),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1986),
.B(n_1997),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1965),
.Y(n_2086)
);

OAI221xp5_ASAP7_75t_L g2087 ( 
.A1(n_1971),
.A2(n_2008),
.B1(n_2004),
.B2(n_1974),
.C(n_1927),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2080),
.B(n_1971),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2073),
.Y(n_2089)
);

NAND2x1_ASAP7_75t_SL g2090 ( 
.A(n_2052),
.B(n_1929),
.Y(n_2090)
);

INVx2_ASAP7_75t_SL g2091 ( 
.A(n_2054),
.Y(n_2091)
);

NOR4xp25_ASAP7_75t_SL g2092 ( 
.A(n_2087),
.B(n_1953),
.C(n_2007),
.D(n_2018),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2034),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_2025),
.B(n_2062),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_2053),
.B(n_1971),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2034),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2053),
.B(n_1971),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_2066),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2064),
.B(n_1930),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2046),
.B(n_2085),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2025),
.B(n_1942),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2058),
.B(n_1942),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2058),
.B(n_1956),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_2025),
.B(n_1946),
.Y(n_2104)
);

AND2x2_ASAP7_75t_L g2105 ( 
.A(n_2025),
.B(n_1946),
.Y(n_2105)
);

INVx2_ASAP7_75t_SL g2106 ( 
.A(n_2054),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2025),
.B(n_1946),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2058),
.B(n_1946),
.Y(n_2108)
);

AND2x4_ASAP7_75t_SL g2109 ( 
.A(n_2028),
.B(n_1945),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_2024),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2079),
.B(n_2001),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2079),
.B(n_2001),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2036),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2062),
.B(n_2001),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2036),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2062),
.B(n_2001),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2048),
.Y(n_2117)
);

INVx4_ASAP7_75t_L g2118 ( 
.A(n_2028),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2071),
.B(n_2002),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2049),
.Y(n_2120)
);

CKINVDCx16_ASAP7_75t_R g2121 ( 
.A(n_2028),
.Y(n_2121)
);

INVx4_ASAP7_75t_L g2122 ( 
.A(n_2041),
.Y(n_2122)
);

INVx2_ASAP7_75t_SL g2123 ( 
.A(n_2054),
.Y(n_2123)
);

INVx2_ASAP7_75t_SL g2124 ( 
.A(n_2054),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2049),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2073),
.B(n_1928),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2067),
.Y(n_2127)
);

AND2x2_ASAP7_75t_SL g2128 ( 
.A(n_2029),
.B(n_1945),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2035),
.A2(n_1927),
.B(n_1957),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2024),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2086),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_2056),
.B(n_1970),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2060),
.B(n_1945),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_2066),
.Y(n_2134)
);

CKINVDCx5p33_ASAP7_75t_R g2135 ( 
.A(n_2055),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2096),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2095),
.B(n_2052),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_2090),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2095),
.B(n_2022),
.Y(n_2139)
);

BUFx3_ASAP7_75t_L g2140 ( 
.A(n_2089),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_2088),
.B(n_2038),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2096),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2113),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2110),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2113),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2120),
.Y(n_2146)
);

HB1xp67_ASAP7_75t_L g2147 ( 
.A(n_2115),
.Y(n_2147)
);

BUFx2_ASAP7_75t_L g2148 ( 
.A(n_2090),
.Y(n_2148)
);

AND2x4_ASAP7_75t_L g2149 ( 
.A(n_2094),
.B(n_2041),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2088),
.B(n_2045),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2120),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2095),
.B(n_2097),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2097),
.B(n_2022),
.Y(n_2153)
);

OR2x2_ASAP7_75t_L g2154 ( 
.A(n_2103),
.B(n_2057),
.Y(n_2154)
);

INVxp67_ASAP7_75t_L g2155 ( 
.A(n_2129),
.Y(n_2155)
);

INVx2_ASAP7_75t_SL g2156 ( 
.A(n_2109),
.Y(n_2156)
);

INVx2_ASAP7_75t_SL g2157 ( 
.A(n_2109),
.Y(n_2157)
);

OR2x2_ASAP7_75t_L g2158 ( 
.A(n_2103),
.B(n_2102),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_2097),
.B(n_2044),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_2110),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2094),
.B(n_2041),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2088),
.B(n_2044),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2125),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2125),
.Y(n_2164)
);

OR2x2_ASAP7_75t_L g2165 ( 
.A(n_2103),
.B(n_2077),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2127),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2108),
.B(n_2039),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2127),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_2094),
.B(n_2054),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2119),
.B(n_2020),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2131),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2131),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2090),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2093),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2108),
.B(n_2039),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2093),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2093),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2117),
.Y(n_2178)
);

OAI22xp33_ASAP7_75t_L g2179 ( 
.A1(n_2129),
.A2(n_2033),
.B1(n_2074),
.B2(n_2037),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2108),
.B(n_1953),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_2110),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2110),
.Y(n_2182)
);

INVx2_ASAP7_75t_L g2183 ( 
.A(n_2130),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2119),
.B(n_2069),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2117),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2119),
.B(n_2077),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2117),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_2115),
.Y(n_2188)
);

AOI322xp5_ASAP7_75t_L g2189 ( 
.A1(n_2128),
.A2(n_2040),
.A3(n_2026),
.B1(n_2023),
.B2(n_2078),
.C1(n_2070),
.C2(n_2082),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_2130),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2098),
.B(n_2072),
.Y(n_2191)
);

INVxp67_ASAP7_75t_L g2192 ( 
.A(n_2191),
.Y(n_2192)
);

AOI21xp33_ASAP7_75t_SL g2193 ( 
.A1(n_2179),
.A2(n_2068),
.B(n_2128),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2139),
.B(n_2118),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_2155),
.B(n_2063),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2136),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2136),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2142),
.Y(n_2198)
);

NAND2xp33_ASAP7_75t_R g2199 ( 
.A(n_2138),
.B(n_2092),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2140),
.Y(n_2200)
);

AND2x2_ASAP7_75t_L g2201 ( 
.A(n_2139),
.B(n_2118),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_2155),
.B(n_2111),
.Y(n_2202)
);

NAND3xp33_ASAP7_75t_L g2203 ( 
.A(n_2189),
.B(n_2092),
.C(n_2065),
.Y(n_2203)
);

AND2x2_ASAP7_75t_L g2204 ( 
.A(n_2139),
.B(n_2118),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2153),
.B(n_2167),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_2191),
.B(n_2111),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2142),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2184),
.B(n_2111),
.Y(n_2208)
);

OR2x4_ASAP7_75t_L g2209 ( 
.A(n_2179),
.B(n_2016),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2143),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2184),
.B(n_2112),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2143),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2153),
.B(n_2118),
.Y(n_2213)
);

HB1xp67_ASAP7_75t_L g2214 ( 
.A(n_2140),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2145),
.Y(n_2215)
);

NOR2x1p5_ASAP7_75t_L g2216 ( 
.A(n_2170),
.B(n_2135),
.Y(n_2216)
);

OAI33xp33_ASAP7_75t_L g2217 ( 
.A1(n_2170),
.A2(n_2102),
.A3(n_2081),
.B1(n_2100),
.B2(n_2132),
.B3(n_2030),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2153),
.B(n_2118),
.Y(n_2218)
);

AND2x4_ASAP7_75t_SL g2219 ( 
.A(n_2169),
.B(n_2043),
.Y(n_2219)
);

OR2x2_ASAP7_75t_L g2220 ( 
.A(n_2141),
.B(n_2098),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2141),
.B(n_2134),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_2150),
.B(n_2031),
.Y(n_2222)
);

OAI31xp33_ASAP7_75t_L g2223 ( 
.A1(n_2184),
.A2(n_2042),
.A3(n_2114),
.B(n_2116),
.Y(n_2223)
);

NOR3xp33_ASAP7_75t_L g2224 ( 
.A(n_2173),
.B(n_2032),
.C(n_2061),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_2140),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2145),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_2167),
.B(n_2121),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2156),
.B(n_2094),
.Y(n_2228)
);

NOR2x1_ASAP7_75t_L g2229 ( 
.A(n_2138),
.B(n_2089),
.Y(n_2229)
);

AND2x4_ASAP7_75t_L g2230 ( 
.A(n_2156),
.B(n_2094),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_2146),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2150),
.B(n_2180),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2180),
.B(n_2112),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2146),
.Y(n_2234)
);

NOR2xp33_ASAP7_75t_L g2235 ( 
.A(n_2169),
.B(n_2135),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2167),
.B(n_2121),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2151),
.Y(n_2237)
);

AND2x2_ASAP7_75t_L g2238 ( 
.A(n_2175),
.B(n_2112),
.Y(n_2238)
);

NOR3xp33_ASAP7_75t_L g2239 ( 
.A(n_2173),
.B(n_2083),
.C(n_2047),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2151),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2163),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2163),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2180),
.B(n_2133),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2175),
.B(n_2133),
.Y(n_2244)
);

AND2x4_ASAP7_75t_SL g2245 ( 
.A(n_2169),
.B(n_2043),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2164),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2227),
.B(n_2169),
.Y(n_2247)
);

OAI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2203),
.A2(n_2189),
.B(n_2128),
.Y(n_2248)
);

CKINVDCx20_ASAP7_75t_R g2249 ( 
.A(n_2235),
.Y(n_2249)
);

INVxp67_ASAP7_75t_SL g2250 ( 
.A(n_2229),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2209),
.B(n_2169),
.Y(n_2251)
);

INVx2_ASAP7_75t_SL g2252 ( 
.A(n_2225),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2207),
.Y(n_2253)
);

OR2x2_ASAP7_75t_L g2254 ( 
.A(n_2206),
.B(n_2175),
.Y(n_2254)
);

OAI22xp5_ASAP7_75t_SL g2255 ( 
.A1(n_2209),
.A2(n_2128),
.B1(n_2076),
.B2(n_2051),
.Y(n_2255)
);

AOI222xp33_ASAP7_75t_L g2256 ( 
.A1(n_2192),
.A2(n_2075),
.B1(n_2012),
.B2(n_1948),
.C1(n_2137),
.C2(n_2138),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2207),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2237),
.Y(n_2258)
);

INVx2_ASAP7_75t_SL g2259 ( 
.A(n_2225),
.Y(n_2259)
);

NOR2x1_ASAP7_75t_L g2260 ( 
.A(n_2216),
.B(n_2148),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2239),
.A2(n_2224),
.B1(n_2223),
.B2(n_2217),
.Y(n_2261)
);

INVxp67_ASAP7_75t_SL g2262 ( 
.A(n_2214),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2237),
.Y(n_2263)
);

AOI21xp33_ASAP7_75t_L g2264 ( 
.A1(n_2199),
.A2(n_2148),
.B(n_2140),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2240),
.Y(n_2265)
);

OR2x2_ASAP7_75t_L g2266 ( 
.A(n_2208),
.B(n_2211),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_2202),
.B(n_2159),
.Y(n_2267)
);

A2O1A1Ixp33_ASAP7_75t_L g2268 ( 
.A1(n_2193),
.A2(n_2148),
.B(n_2104),
.C(n_2105),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2195),
.B(n_2159),
.Y(n_2269)
);

OAI21xp33_ASAP7_75t_L g2270 ( 
.A1(n_2232),
.A2(n_2137),
.B(n_2116),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2222),
.B(n_2159),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2240),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2205),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2196),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2209),
.A2(n_2149),
.B1(n_2161),
.B2(n_2114),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2227),
.A2(n_2157),
.B1(n_2156),
.B2(n_2059),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2238),
.B(n_2205),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_SL g2278 ( 
.A(n_2236),
.B(n_2157),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2197),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2198),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_SL g2281 ( 
.A1(n_2236),
.A2(n_2161),
.B(n_2149),
.Y(n_2281)
);

OAI221xp5_ASAP7_75t_SL g2282 ( 
.A1(n_2220),
.A2(n_2137),
.B1(n_2102),
.B2(n_2158),
.C(n_2114),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2238),
.B(n_2162),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2200),
.B(n_2162),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2200),
.B(n_2162),
.Y(n_2285)
);

AOI221xp5_ASAP7_75t_L g2286 ( 
.A1(n_2210),
.A2(n_2149),
.B1(n_2161),
.B2(n_2152),
.C(n_2157),
.Y(n_2286)
);

NOR2x1_ASAP7_75t_SL g2287 ( 
.A(n_2194),
.B(n_2201),
.Y(n_2287)
);

AND2x4_ASAP7_75t_SL g2288 ( 
.A(n_2228),
.B(n_2149),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2248),
.B(n_2233),
.Y(n_2289)
);

AOI221xp5_ASAP7_75t_L g2290 ( 
.A1(n_2261),
.A2(n_2228),
.B1(n_2230),
.B2(n_2246),
.C(n_2215),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2255),
.A2(n_2230),
.B1(n_2228),
.B2(n_2149),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2262),
.Y(n_2292)
);

AOI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2261),
.A2(n_2230),
.B1(n_2161),
.B2(n_2219),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2262),
.Y(n_2294)
);

A2O1A1Ixp33_ASAP7_75t_L g2295 ( 
.A1(n_2268),
.A2(n_2107),
.B(n_2104),
.C(n_2105),
.Y(n_2295)
);

HB1xp67_ASAP7_75t_L g2296 ( 
.A(n_2250),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2250),
.A2(n_2122),
.B1(n_2007),
.B2(n_2021),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2252),
.B(n_2194),
.Y(n_2298)
);

OAI21xp5_ASAP7_75t_L g2299 ( 
.A1(n_2268),
.A2(n_2204),
.B(n_2201),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2253),
.Y(n_2300)
);

OAI221xp5_ASAP7_75t_L g2301 ( 
.A1(n_2260),
.A2(n_2220),
.B1(n_2221),
.B2(n_2244),
.C(n_2218),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2257),
.Y(n_2302)
);

A2O1A1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2275),
.A2(n_2105),
.B(n_2107),
.C(n_2104),
.Y(n_2303)
);

OR2x2_ASAP7_75t_L g2304 ( 
.A(n_2269),
.B(n_2266),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2258),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2259),
.B(n_2204),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2288),
.Y(n_2307)
);

AND2x2_ASAP7_75t_L g2308 ( 
.A(n_2247),
.B(n_2219),
.Y(n_2308)
);

O2A1O1Ixp5_ASAP7_75t_L g2309 ( 
.A1(n_2278),
.A2(n_2213),
.B(n_2218),
.C(n_2161),
.Y(n_2309)
);

OAI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_2264),
.A2(n_2122),
.B1(n_2221),
.B2(n_2055),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2256),
.B(n_2213),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2263),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2249),
.B(n_2251),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2265),
.Y(n_2314)
);

AND2x4_ASAP7_75t_L g2315 ( 
.A(n_2287),
.B(n_2245),
.Y(n_2315)
);

NAND3xp33_ASAP7_75t_L g2316 ( 
.A(n_2251),
.B(n_2278),
.C(n_2286),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2272),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2271),
.B(n_2243),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2288),
.B(n_2245),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2292),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2294),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2290),
.B(n_2273),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_SL g2323 ( 
.A(n_2297),
.B(n_2276),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2296),
.Y(n_2324)
);

XOR2x2_ASAP7_75t_L g2325 ( 
.A(n_2313),
.B(n_2282),
.Y(n_2325)
);

NAND2xp5_ASAP7_75t_SL g2326 ( 
.A(n_2297),
.B(n_2273),
.Y(n_2326)
);

HB1xp67_ASAP7_75t_L g2327 ( 
.A(n_2296),
.Y(n_2327)
);

OR2x2_ASAP7_75t_L g2328 ( 
.A(n_2304),
.B(n_2254),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2300),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2289),
.B(n_2277),
.Y(n_2330)
);

INVxp67_ASAP7_75t_SL g2331 ( 
.A(n_2313),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2293),
.B(n_2274),
.Y(n_2332)
);

OR2x2_ASAP7_75t_L g2333 ( 
.A(n_2318),
.B(n_2285),
.Y(n_2333)
);

XNOR2xp5_ASAP7_75t_L g2334 ( 
.A(n_2291),
.B(n_2043),
.Y(n_2334)
);

AOI31xp33_ASAP7_75t_L g2335 ( 
.A1(n_2316),
.A2(n_2267),
.A3(n_2284),
.B(n_2270),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2307),
.B(n_2279),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2302),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2311),
.B(n_2298),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2305),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2315),
.B(n_2281),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_SL g2341 ( 
.A(n_2310),
.B(n_2280),
.C(n_2283),
.Y(n_2341)
);

INVx2_ASAP7_75t_SL g2342 ( 
.A(n_2315),
.Y(n_2342)
);

NOR2x1_ASAP7_75t_L g2343 ( 
.A(n_2324),
.B(n_2310),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2331),
.B(n_2306),
.Y(n_2344)
);

AOI211xp5_ASAP7_75t_SL g2345 ( 
.A1(n_2327),
.A2(n_2301),
.B(n_2295),
.C(n_2303),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2342),
.B(n_2309),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2342),
.B(n_2308),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_SL g2348 ( 
.A(n_2340),
.B(n_2295),
.Y(n_2348)
);

OA211x2_ASAP7_75t_L g2349 ( 
.A1(n_2323),
.A2(n_2299),
.B(n_2303),
.C(n_2100),
.Y(n_2349)
);

NAND3xp33_ASAP7_75t_L g2350 ( 
.A(n_2341),
.B(n_2314),
.C(n_2312),
.Y(n_2350)
);

NOR3xp33_ASAP7_75t_L g2351 ( 
.A(n_2338),
.B(n_2317),
.C(n_2319),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2325),
.B(n_2212),
.Y(n_2352)
);

OAI32xp33_ASAP7_75t_L g2353 ( 
.A1(n_2322),
.A2(n_2158),
.A3(n_2188),
.B1(n_2147),
.B2(n_2231),
.Y(n_2353)
);

NOR3xp33_ASAP7_75t_L g2354 ( 
.A(n_2332),
.B(n_2122),
.C(n_2226),
.Y(n_2354)
);

OR2x2_ASAP7_75t_L g2355 ( 
.A(n_2328),
.B(n_2154),
.Y(n_2355)
);

NOR2xp67_ASAP7_75t_L g2356 ( 
.A(n_2328),
.B(n_2234),
.Y(n_2356)
);

NOR2x1_ASAP7_75t_L g2357 ( 
.A(n_2320),
.B(n_2241),
.Y(n_2357)
);

AOI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2343),
.A2(n_2325),
.B(n_2323),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2356),
.Y(n_2359)
);

NAND3xp33_ASAP7_75t_L g2360 ( 
.A(n_2345),
.B(n_2321),
.C(n_2326),
.Y(n_2360)
);

NOR4xp25_ASAP7_75t_SL g2361 ( 
.A(n_2346),
.B(n_2348),
.C(n_2326),
.D(n_2339),
.Y(n_2361)
);

AOI221xp5_ASAP7_75t_L g2362 ( 
.A1(n_2350),
.A2(n_2335),
.B1(n_2330),
.B2(n_2336),
.C(n_2329),
.Y(n_2362)
);

O2A1O1Ixp33_ASAP7_75t_L g2363 ( 
.A1(n_2352),
.A2(n_2337),
.B(n_2340),
.C(n_2333),
.Y(n_2363)
);

AOI211xp5_ASAP7_75t_L g2364 ( 
.A1(n_2353),
.A2(n_2334),
.B(n_2333),
.C(n_2158),
.Y(n_2364)
);

OAI211xp5_ASAP7_75t_L g2365 ( 
.A1(n_2345),
.A2(n_2344),
.B(n_2351),
.C(n_2347),
.Y(n_2365)
);

AOI221xp5_ASAP7_75t_L g2366 ( 
.A1(n_2354),
.A2(n_2242),
.B1(n_2089),
.B2(n_2188),
.C(n_2147),
.Y(n_2366)
);

OAI21xp5_ASAP7_75t_L g2367 ( 
.A1(n_2357),
.A2(n_2355),
.B(n_2349),
.Y(n_2367)
);

O2A1O1Ixp33_ASAP7_75t_L g2368 ( 
.A1(n_2348),
.A2(n_2106),
.B(n_2124),
.C(n_2091),
.Y(n_2368)
);

NAND5xp2_ASAP7_75t_L g2369 ( 
.A(n_2345),
.B(n_2019),
.C(n_2107),
.D(n_2116),
.E(n_2101),
.Y(n_2369)
);

AOI221x1_ASAP7_75t_L g2370 ( 
.A1(n_2350),
.A2(n_2176),
.B1(n_2174),
.B2(n_2187),
.C(n_2177),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2347),
.Y(n_2371)
);

NOR2x1_ASAP7_75t_L g2372 ( 
.A(n_2343),
.B(n_2174),
.Y(n_2372)
);

INVx1_ASAP7_75t_SL g2373 ( 
.A(n_2371),
.Y(n_2373)
);

AOI322xp5_ASAP7_75t_L g2374 ( 
.A1(n_2372),
.A2(n_2152),
.A3(n_2005),
.B1(n_2101),
.B2(n_1983),
.C1(n_2126),
.C2(n_2099),
.Y(n_2374)
);

BUFx2_ASAP7_75t_L g2375 ( 
.A(n_2359),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2363),
.Y(n_2376)
);

AOI221xp5_ASAP7_75t_L g2377 ( 
.A1(n_2358),
.A2(n_2360),
.B1(n_2369),
.B2(n_2362),
.C(n_2365),
.Y(n_2377)
);

INVx2_ASAP7_75t_L g2378 ( 
.A(n_2367),
.Y(n_2378)
);

NOR2xp33_ASAP7_75t_R g2379 ( 
.A(n_2361),
.B(n_2050),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2368),
.Y(n_2380)
);

OAI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2364),
.A2(n_2091),
.B1(n_2106),
.B2(n_2124),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2375),
.Y(n_2382)
);

NAND4xp75_ASAP7_75t_L g2383 ( 
.A(n_2377),
.B(n_2370),
.C(n_2366),
.D(n_2101),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2373),
.B(n_2154),
.Y(n_2384)
);

OAI221xp5_ASAP7_75t_L g2385 ( 
.A1(n_2376),
.A2(n_2124),
.B1(n_2123),
.B2(n_2091),
.C(n_2106),
.Y(n_2385)
);

NOR3xp33_ASAP7_75t_SL g2386 ( 
.A(n_2381),
.B(n_2084),
.C(n_2011),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_L g2387 ( 
.A(n_2378),
.B(n_2380),
.C(n_2379),
.Y(n_2387)
);

NOR3xp33_ASAP7_75t_L g2388 ( 
.A(n_2374),
.B(n_2122),
.C(n_2123),
.Y(n_2388)
);

OAI221xp5_ASAP7_75t_SL g2389 ( 
.A1(n_2374),
.A2(n_2123),
.B1(n_2154),
.B2(n_2152),
.C(n_2027),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2382),
.B(n_2164),
.Y(n_2390)
);

AOI21xp5_ASAP7_75t_L g2391 ( 
.A1(n_2387),
.A2(n_2183),
.B(n_2190),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2384),
.Y(n_2392)
);

BUFx2_ASAP7_75t_L g2393 ( 
.A(n_2383),
.Y(n_2393)
);

NAND5xp2_ASAP7_75t_L g2394 ( 
.A(n_2388),
.B(n_2389),
.C(n_2385),
.D(n_2386),
.E(n_1983),
.Y(n_2394)
);

AOI31xp33_ASAP7_75t_L g2395 ( 
.A1(n_2382),
.A2(n_2027),
.A3(n_1957),
.B(n_2015),
.Y(n_2395)
);

OAI211xp5_ASAP7_75t_SL g2396 ( 
.A1(n_2387),
.A2(n_2132),
.B(n_2160),
.C(n_2181),
.Y(n_2396)
);

INVxp67_ASAP7_75t_L g2397 ( 
.A(n_2393),
.Y(n_2397)
);

CKINVDCx20_ASAP7_75t_R g2398 ( 
.A(n_2392),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2390),
.Y(n_2399)
);

CKINVDCx12_ASAP7_75t_R g2400 ( 
.A(n_2396),
.Y(n_2400)
);

AND2x4_ASAP7_75t_L g2401 ( 
.A(n_2391),
.B(n_2186),
.Y(n_2401)
);

AOI22xp5_ASAP7_75t_L g2402 ( 
.A1(n_2398),
.A2(n_2394),
.B1(n_2395),
.B2(n_2122),
.Y(n_2402)
);

INVxp67_ASAP7_75t_SL g2403 ( 
.A(n_2397),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2403),
.A2(n_2400),
.B1(n_2401),
.B2(n_2399),
.Y(n_2404)
);

HB1xp67_ASAP7_75t_L g2405 ( 
.A(n_2404),
.Y(n_2405)
);

INVxp67_ASAP7_75t_L g2406 ( 
.A(n_2404),
.Y(n_2406)
);

OAI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_2406),
.A2(n_2402),
.B1(n_2144),
.B2(n_2190),
.Y(n_2407)
);

AOI221xp5_ASAP7_75t_L g2408 ( 
.A1(n_2405),
.A2(n_2171),
.B1(n_2168),
.B2(n_2172),
.C(n_2166),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2407),
.A2(n_2160),
.B1(n_2190),
.B2(n_2144),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2408),
.Y(n_2410)
);

AOI322xp5_ASAP7_75t_L g2411 ( 
.A1(n_2410),
.A2(n_2126),
.A3(n_2187),
.B1(n_2176),
.B2(n_2185),
.C1(n_2177),
.C2(n_2178),
.Y(n_2411)
);

AOI22xp33_ASAP7_75t_L g2412 ( 
.A1(n_2411),
.A2(n_2409),
.B1(n_2182),
.B2(n_2160),
.Y(n_2412)
);

AOI211xp5_ASAP7_75t_L g2413 ( 
.A1(n_2412),
.A2(n_2165),
.B(n_2172),
.C(n_2171),
.Y(n_2413)
);


endmodule