module fake_netlist_6_3518_n_779 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_779);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_779;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_703;
wire n_578;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_685;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_658;
wire n_616;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx2_ASAP7_75t_SL g154 ( 
.A(n_8),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_19),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_71),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_34),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_52),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_139),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_76),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_1),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_50),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_40),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_152),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_88),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_68),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_102),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_27),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_5),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_70),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_62),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_73),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_28),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_33),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_54),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_119),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_42),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_61),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_19),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_48),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_9),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_59),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_103),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_55),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_149),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_81),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_35),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_32),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_120),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_23),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_156),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_165),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_189),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_187),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_167),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_167),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_0),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_163),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_0),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_169),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_24),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_159),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_175),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_182),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_163),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_179),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_185),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_193),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_170),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_206),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_170),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_154),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_177),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_243),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_226),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_157),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_224),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_232),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_158),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_238),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_192),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_220),
.B(n_164),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_215),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_211),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_217),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_210),
.B(n_161),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_229),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_208),
.A2(n_186),
.B1(n_183),
.B2(n_171),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_240),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_207),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_196),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_208),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_209),
.B(n_198),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_218),
.B(n_199),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_164),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_257),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_277),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_270),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_249),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_260),
.B(n_183),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_160),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_249),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_250),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_282),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_257),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_255),
.B(n_164),
.Y(n_317)
);

INVx8_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_186),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_271),
.B(n_161),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_255),
.A2(n_256),
.B1(n_268),
.B2(n_273),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_164),
.Y(n_325)
);

AND2x4_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_162),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_237),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_281),
.B(n_161),
.Y(n_328)
);

AO21x2_ASAP7_75t_L g329 ( 
.A1(n_253),
.A2(n_172),
.B(n_204),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_273),
.B(n_237),
.Y(n_330)
);

OR2x2_ASAP7_75t_SL g331 ( 
.A(n_290),
.B(n_241),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_256),
.B(n_188),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_280),
.B(n_173),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_261),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_200),
.Y(n_335)
);

NAND2x1p5_ASAP7_75t_L g336 ( 
.A(n_272),
.B(n_197),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_256),
.B(n_202),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_261),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_203),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_281),
.B(n_197),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_275),
.B(n_197),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_2),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_270),
.B(n_272),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_256),
.B(n_25),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_247),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_263),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_247),
.Y(n_350)
);

AND2x4_ASAP7_75t_SL g351 ( 
.A(n_283),
.B(n_241),
.Y(n_351)
);

AND2x6_ASAP7_75t_L g352 ( 
.A(n_272),
.B(n_26),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_265),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_250),
.B(n_29),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_250),
.B(n_151),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_285),
.Y(n_357)
);

AO22x2_ASAP7_75t_L g358 ( 
.A1(n_327),
.A2(n_307),
.B1(n_292),
.B2(n_288),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_250),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_349),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_274),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_250),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_335),
.B(n_264),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_299),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_349),
.A2(n_292),
.B1(n_288),
.B2(n_276),
.Y(n_368)
);

AO22x2_ASAP7_75t_L g369 ( 
.A1(n_330),
.A2(n_293),
.B1(n_289),
.B2(n_284),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_357),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_310),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_274),
.Y(n_372)
);

OAI221xp5_ASAP7_75t_L g373 ( 
.A1(n_309),
.A2(n_269),
.B1(n_252),
.B2(n_254),
.C(n_259),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_348),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_315),
.Y(n_378)
);

AO22x2_ASAP7_75t_L g379 ( 
.A1(n_328),
.A2(n_293),
.B1(n_289),
.B2(n_284),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

AO22x2_ASAP7_75t_L g381 ( 
.A1(n_340),
.A2(n_291),
.B1(n_278),
.B2(n_287),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g382 ( 
.A1(n_322),
.A2(n_286),
.B1(n_269),
.B2(n_267),
.Y(n_382)
);

NAND2x1p5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_283),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_353),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_317),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_343),
.B(n_283),
.Y(n_386)
);

AO22x2_ASAP7_75t_L g387 ( 
.A1(n_326),
.A2(n_267),
.B1(n_3),
.B2(n_4),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

AO22x2_ASAP7_75t_L g391 ( 
.A1(n_326),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_317),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_344),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_337),
.A2(n_283),
.B1(n_265),
.B2(n_254),
.Y(n_394)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_347),
.A2(n_325),
.B(n_336),
.Y(n_395)
);

OAI221xp5_ASAP7_75t_L g396 ( 
.A1(n_309),
.A2(n_259),
.B1(n_252),
.B2(n_265),
.C(n_248),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_339),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_337),
.A2(n_283),
.B1(n_265),
.B2(n_248),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_305),
.Y(n_399)
);

AO22x2_ASAP7_75t_L g400 ( 
.A1(n_333),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_339),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_302),
.B(n_251),
.Y(n_402)
);

OAI221xp5_ASAP7_75t_L g403 ( 
.A1(n_342),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.C(n_10),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_325),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_266),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

OR2x2_ASAP7_75t_SL g407 ( 
.A(n_331),
.B(n_10),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_298),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_329),
.A2(n_266),
.B1(n_89),
.B2(n_90),
.Y(n_409)
);

OAI221xp5_ASAP7_75t_L g410 ( 
.A1(n_323),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_329),
.B(n_266),
.Y(n_411)
);

AO22x2_ASAP7_75t_L g412 ( 
.A1(n_333),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_412)
);

AO22x2_ASAP7_75t_L g413 ( 
.A1(n_347),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_308),
.Y(n_414)
);

AO22x2_ASAP7_75t_L g415 ( 
.A1(n_336),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_316),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_319),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_295),
.A2(n_266),
.B1(n_96),
.B2(n_97),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_298),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_303),
.B(n_30),
.Y(n_420)
);

A2O1A1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_300),
.A2(n_266),
.B(n_20),
.C(n_21),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_298),
.Y(n_423)
);

NAND2x1p5_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_338),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_318),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_SL g427 ( 
.A(n_420),
.B(n_318),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_401),
.B(n_300),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_365),
.B(n_300),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_380),
.B(n_301),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_390),
.B(n_301),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_360),
.B(n_351),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_402),
.B(n_301),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_318),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_295),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_420),
.B(n_362),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g437 ( 
.A(n_361),
.B(n_354),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_385),
.B(n_295),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_378),
.B(n_334),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_371),
.B(n_334),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_371),
.B(n_338),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_367),
.B(n_338),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_372),
.B(n_354),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_372),
.B(n_356),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_394),
.B(n_356),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_398),
.B(n_312),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_370),
.B(n_312),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_SL g448 ( 
.A(n_388),
.B(n_297),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_SL g449 ( 
.A(n_363),
.B(n_297),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_383),
.B(n_314),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_366),
.B(n_314),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_374),
.B(n_297),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_386),
.B(n_352),
.Y(n_453)
);

NAND2xp33_ASAP7_75t_SL g454 ( 
.A(n_411),
.B(n_352),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_395),
.B(n_375),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_376),
.B(n_352),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_377),
.B(n_352),
.Y(n_457)
);

NAND2xp33_ASAP7_75t_SL g458 ( 
.A(n_405),
.B(n_296),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_384),
.B(n_296),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_392),
.B(n_296),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_368),
.B(n_18),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_404),
.B(n_296),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_419),
.B(n_296),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_266),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_359),
.B(n_31),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_364),
.B(n_36),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_368),
.B(n_18),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_408),
.B(n_37),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_408),
.B(n_38),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_409),
.B(n_39),
.Y(n_470)
);

NAND2xp33_ASAP7_75t_SL g471 ( 
.A(n_423),
.B(n_20),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_266),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_382),
.B(n_21),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_389),
.B(n_41),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_382),
.B(n_22),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_369),
.B(n_22),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g477 ( 
.A(n_422),
.B(n_23),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_373),
.B(n_43),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_393),
.B(n_44),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_399),
.B(n_46),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_414),
.B(n_47),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g482 ( 
.A(n_436),
.B(n_403),
.C(n_410),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_432),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_445),
.A2(n_396),
.B(n_416),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_435),
.A2(n_424),
.B(n_417),
.Y(n_485)
);

A2O1A1Ixp33_ASAP7_75t_L g486 ( 
.A1(n_478),
.A2(n_421),
.B(n_418),
.C(n_358),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_438),
.A2(n_379),
.B(n_51),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_379),
.B(n_53),
.Y(n_488)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_461),
.Y(n_489)
);

AO31x2_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_358),
.A3(n_415),
.B(n_413),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_467),
.Y(n_491)
);

BUFx8_ASAP7_75t_L g492 ( 
.A(n_476),
.Y(n_492)
);

AOI221xp5_ASAP7_75t_SL g493 ( 
.A1(n_475),
.A2(n_407),
.B1(n_413),
.B2(n_415),
.C(n_412),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_442),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_443),
.A2(n_381),
.B(n_387),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_427),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_L g497 ( 
.A1(n_434),
.A2(n_381),
.B(n_387),
.Y(n_497)
);

OR2x6_ASAP7_75t_L g498 ( 
.A(n_428),
.B(n_391),
.Y(n_498)
);

OAI22x1_ASAP7_75t_L g499 ( 
.A1(n_439),
.A2(n_412),
.B1(n_400),
.B2(n_391),
.Y(n_499)
);

AOI21x1_ASAP7_75t_SL g500 ( 
.A1(n_426),
.A2(n_400),
.B(n_369),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_437),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_457),
.A2(n_58),
.B(n_60),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_444),
.A2(n_64),
.B(n_65),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

AO21x1_ASAP7_75t_L g505 ( 
.A1(n_454),
.A2(n_66),
.B(n_67),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_441),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_69),
.Y(n_507)
);

O2A1O1Ixp33_ASAP7_75t_L g508 ( 
.A1(n_431),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_477),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_429),
.B(n_77),
.Y(n_510)
);

OAI21x1_ASAP7_75t_SL g511 ( 
.A1(n_464),
.A2(n_78),
.B(n_79),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_455),
.A2(n_82),
.B(n_83),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_472),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_453),
.A2(n_84),
.B(n_85),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_452),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_433),
.B(n_150),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_462),
.A2(n_86),
.B(n_87),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_459),
.Y(n_518)
);

A2O1A1Ixp33_ASAP7_75t_L g519 ( 
.A1(n_470),
.A2(n_92),
.B(n_93),
.C(n_94),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_447),
.B(n_148),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_446),
.A2(n_98),
.B(n_99),
.Y(n_521)
);

NOR2x1p5_ASAP7_75t_L g522 ( 
.A(n_471),
.B(n_100),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_448),
.Y(n_523)
);

AOI221xp5_ASAP7_75t_L g524 ( 
.A1(n_458),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.C(n_106),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_474),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_465),
.A2(n_107),
.B(n_108),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_466),
.A2(n_110),
.B(n_111),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_474),
.B(n_146),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_479),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_485),
.A2(n_481),
.B(n_480),
.Y(n_530)
);

AO21x2_ASAP7_75t_L g531 ( 
.A1(n_487),
.A2(n_481),
.B(n_480),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_490),
.B(n_479),
.Y(n_532)
);

CKINVDCx14_ASAP7_75t_R g533 ( 
.A(n_491),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_488),
.A2(n_469),
.B(n_468),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_490),
.B(n_451),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_483),
.B(n_449),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_490),
.B(n_450),
.Y(n_537)
);

OA21x2_ASAP7_75t_L g538 ( 
.A1(n_484),
.A2(n_460),
.B(n_463),
.Y(n_538)
);

AO21x2_ASAP7_75t_L g539 ( 
.A1(n_486),
.A2(n_112),
.B(n_113),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_518),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_514),
.Y(n_541)
);

OA21x2_ASAP7_75t_L g542 ( 
.A1(n_512),
.A2(n_114),
.B(n_115),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_504),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_489),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_502),
.A2(n_116),
.B(n_118),
.Y(n_546)
);

AOI211xp5_ASAP7_75t_L g547 ( 
.A1(n_497),
.A2(n_122),
.B(n_123),
.C(n_124),
.Y(n_547)
);

AO31x2_ASAP7_75t_L g548 ( 
.A1(n_505),
.A2(n_125),
.A3(n_127),
.B(n_128),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_506),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g550 ( 
.A1(n_517),
.A2(n_129),
.B(n_130),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_131),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_496),
.B(n_132),
.Y(n_552)
);

O2A1O1Ixp33_ASAP7_75t_L g553 ( 
.A1(n_509),
.A2(n_133),
.B(n_135),
.C(n_136),
.Y(n_553)
);

AO21x2_ASAP7_75t_L g554 ( 
.A1(n_495),
.A2(n_137),
.B(n_138),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_507),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_489),
.B(n_144),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_496),
.Y(n_557)
);

OA21x2_ASAP7_75t_L g558 ( 
.A1(n_529),
.A2(n_145),
.B(n_497),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_482),
.B(n_493),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_494),
.B(n_493),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g561 ( 
.A(n_498),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_513),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g563 ( 
.A(n_498),
.Y(n_563)
);

NAND2x1_ASAP7_75t_L g564 ( 
.A(n_511),
.B(n_528),
.Y(n_564)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_526),
.A2(n_527),
.B(n_524),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_515),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_522),
.A2(n_523),
.B1(n_498),
.B2(n_489),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_499),
.B(n_510),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_520),
.B(n_516),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_501),
.A2(n_519),
.B1(n_521),
.B2(n_503),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_540),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_540),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_532),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_530),
.A2(n_501),
.B(n_500),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_532),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_558),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_544),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_558),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_557),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_558),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_539),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_539),
.Y(n_582)
);

AOI21xp33_ASAP7_75t_L g583 ( 
.A1(n_570),
.A2(n_508),
.B(n_492),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_557),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_559),
.B(n_492),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_539),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_557),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_537),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_530),
.A2(n_534),
.B(n_564),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_537),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_565),
.A2(n_569),
.B(n_564),
.Y(n_591)
);

CKINVDCx6p67_ASAP7_75t_R g592 ( 
.A(n_556),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_560),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_531),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_543),
.Y(n_596)
);

OAI21x1_ASAP7_75t_L g597 ( 
.A1(n_534),
.A2(n_550),
.B(n_546),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_531),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_535),
.B(n_568),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_566),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_535),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_549),
.B(n_562),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_531),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_562),
.B(n_547),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_554),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_554),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_554),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_538),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_548),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_548),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_548),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_538),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_R g616 ( 
.A(n_592),
.B(n_533),
.Y(n_616)
);

BUFx10_ASAP7_75t_L g617 ( 
.A(n_577),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_R g618 ( 
.A(n_604),
.B(n_556),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_585),
.B(n_552),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_596),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_594),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_R g622 ( 
.A(n_592),
.B(n_545),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_594),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_R g624 ( 
.A(n_604),
.B(n_536),
.Y(n_624)
);

NAND2xp33_ASAP7_75t_SL g625 ( 
.A(n_585),
.B(n_545),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_602),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_R g627 ( 
.A(n_602),
.B(n_542),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_R g628 ( 
.A(n_592),
.B(n_563),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_R g629 ( 
.A(n_574),
.B(n_542),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_R g630 ( 
.A(n_571),
.B(n_561),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_567),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_R g632 ( 
.A(n_572),
.B(n_584),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_587),
.B(n_552),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_596),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_R g635 ( 
.A(n_572),
.B(n_541),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_600),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_R g637 ( 
.A(n_579),
.B(n_541),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_590),
.B(n_555),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_579),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_590),
.B(n_552),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_R g641 ( 
.A(n_579),
.B(n_551),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_600),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_587),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_579),
.B(n_548),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_599),
.B(n_542),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_584),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_584),
.B(n_587),
.Y(n_647)
);

BUFx10_ASAP7_75t_L g648 ( 
.A(n_588),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_R g649 ( 
.A(n_584),
.B(n_553),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_593),
.B(n_565),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_R g651 ( 
.A(n_599),
.B(n_542),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_588),
.B(n_546),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_610),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_620),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_645),
.B(n_575),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_646),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_636),
.B(n_593),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_640),
.B(n_575),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_626),
.B(n_601),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_623),
.B(n_601),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_650),
.B(n_573),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_573),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_621),
.B(n_591),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_653),
.Y(n_664)
);

INVx1_ASAP7_75t_SL g665 ( 
.A(n_632),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_634),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_652),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_644),
.B(n_615),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_652),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_647),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_635),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_642),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_619),
.B(n_595),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_631),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_638),
.A2(n_565),
.B1(n_631),
.B2(n_619),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_647),
.B(n_591),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_648),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_648),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_651),
.B(n_615),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_639),
.B(n_609),
.Y(n_680)
);

AND2x4_ASAP7_75t_SL g681 ( 
.A(n_674),
.B(n_617),
.Y(n_681)
);

NAND4xp25_ASAP7_75t_L g682 ( 
.A(n_663),
.B(n_624),
.C(n_618),
.D(n_625),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_672),
.B(n_617),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_658),
.B(n_630),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_675),
.B(n_583),
.C(n_627),
.Y(n_685)
);

AOI221xp5_ASAP7_75t_L g686 ( 
.A1(n_675),
.A2(n_583),
.B1(n_612),
.B2(n_614),
.C(n_613),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_654),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_654),
.Y(n_688)
);

OAI221xp5_ASAP7_75t_L g689 ( 
.A1(n_665),
.A2(n_629),
.B1(n_633),
.B2(n_581),
.C(n_607),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_657),
.B(n_609),
.Y(n_690)
);

AO21x2_ASAP7_75t_L g691 ( 
.A1(n_657),
.A2(n_606),
.B(n_605),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_664),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_671),
.A2(n_565),
.B1(n_628),
.B2(n_607),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_658),
.B(n_616),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_664),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_665),
.A2(n_633),
.B1(n_581),
.B2(n_582),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_687),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_684),
.B(n_670),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_683),
.B(n_666),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_690),
.B(n_666),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_688),
.B(n_661),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_692),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_694),
.B(n_670),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_681),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_692),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_695),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_695),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_700),
.B(n_681),
.Y(n_708)
);

OAI221xp5_ASAP7_75t_L g709 ( 
.A1(n_699),
.A2(n_685),
.B1(n_682),
.B2(n_686),
.C(n_693),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_701),
.B(n_693),
.Y(n_710)
);

AO221x2_ASAP7_75t_L g711 ( 
.A1(n_697),
.A2(n_696),
.B1(n_677),
.B2(n_669),
.C(n_667),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_703),
.B(n_667),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_712),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_710),
.B(n_706),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_711),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_708),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_709),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_708),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_713),
.Y(n_719)
);

CKINVDCx8_ASAP7_75t_R g720 ( 
.A(n_717),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_714),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_714),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_721),
.B(n_715),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_722),
.B(n_718),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_719),
.B(n_716),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_719),
.B(n_704),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_725),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_723),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_724),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_726),
.Y(n_730)
);

OAI221xp5_ASAP7_75t_L g731 ( 
.A1(n_729),
.A2(n_720),
.B1(n_689),
.B2(n_656),
.C(n_671),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_730),
.B(n_698),
.Y(n_732)
);

NOR3xp33_ASAP7_75t_L g733 ( 
.A(n_728),
.B(n_656),
.C(n_677),
.Y(n_733)
);

NAND5xp2_ASAP7_75t_L g734 ( 
.A(n_727),
.B(n_679),
.C(n_669),
.D(n_622),
.E(n_662),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_728),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_727),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_SL g737 ( 
.A(n_730),
.B(n_696),
.C(n_660),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_728),
.B(n_678),
.C(n_656),
.Y(n_738)
);

AOI222xp33_ASAP7_75t_L g739 ( 
.A1(n_736),
.A2(n_613),
.B1(n_608),
.B2(n_612),
.C1(n_614),
.C2(n_679),
.Y(n_739)
);

NAND4xp25_ASAP7_75t_L g740 ( 
.A(n_735),
.B(n_659),
.C(n_678),
.D(n_676),
.Y(n_740)
);

AOI211xp5_ASAP7_75t_L g741 ( 
.A1(n_731),
.A2(n_649),
.B(n_641),
.C(n_678),
.Y(n_741)
);

OAI221xp5_ASAP7_75t_SL g742 ( 
.A1(n_733),
.A2(n_673),
.B1(n_667),
.B2(n_661),
.C(n_707),
.Y(n_742)
);

AOI221xp5_ASAP7_75t_L g743 ( 
.A1(n_737),
.A2(n_738),
.B1(n_732),
.B2(n_734),
.C(n_702),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_737),
.A2(n_706),
.B(n_705),
.C(n_702),
.Y(n_744)
);

AOI222xp33_ASAP7_75t_L g745 ( 
.A1(n_736),
.A2(n_608),
.B1(n_606),
.B2(n_605),
.C1(n_586),
.C2(n_582),
.Y(n_745)
);

OAI211xp5_ASAP7_75t_L g746 ( 
.A1(n_735),
.A2(n_637),
.B(n_705),
.C(n_586),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_740),
.Y(n_748)
);

AOI22xp5_ASAP7_75t_L g749 ( 
.A1(n_743),
.A2(n_691),
.B1(n_676),
.B2(n_670),
.Y(n_749)
);

NAND4xp75_ASAP7_75t_L g750 ( 
.A(n_741),
.B(n_746),
.C(n_742),
.D(n_739),
.Y(n_750)
);

INVxp33_ASAP7_75t_L g751 ( 
.A(n_745),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_744),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_744),
.Y(n_753)
);

NAND4xp75_ASAP7_75t_L g754 ( 
.A(n_743),
.B(n_680),
.C(n_538),
.D(n_574),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_747),
.B(n_676),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_R g756 ( 
.A(n_752),
.B(n_670),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_753),
.B(n_673),
.C(n_676),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_R g758 ( 
.A(n_748),
.B(n_643),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_751),
.B(n_691),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_750),
.B(n_643),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_749),
.B(n_680),
.Y(n_761)
);

INVx4_ASAP7_75t_L g762 ( 
.A(n_758),
.Y(n_762)
);

NOR2x1_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_754),
.Y(n_763)
);

OAI211xp5_ASAP7_75t_SL g764 ( 
.A1(n_755),
.A2(n_761),
.B(n_760),
.C(n_756),
.Y(n_764)
);

OAI22xp5_ASAP7_75t_L g765 ( 
.A1(n_759),
.A2(n_664),
.B1(n_586),
.B2(n_582),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_759),
.A2(n_589),
.B(n_597),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_764),
.A2(n_662),
.B1(n_668),
.B2(n_655),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_766),
.A2(n_597),
.B(n_589),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_763),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_762),
.Y(n_770)
);

OAI21xp33_ASAP7_75t_L g771 ( 
.A1(n_769),
.A2(n_765),
.B(n_668),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_770),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_767),
.A2(n_655),
.B1(n_574),
.B2(n_611),
.Y(n_773)
);

AOI31xp33_ASAP7_75t_L g774 ( 
.A1(n_772),
.A2(n_768),
.A3(n_576),
.B(n_578),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_774),
.A2(n_771),
.B(n_773),
.C(n_576),
.Y(n_775)
);

AOI222xp33_ASAP7_75t_L g776 ( 
.A1(n_775),
.A2(n_611),
.B1(n_578),
.B2(n_580),
.C1(n_610),
.C2(n_597),
.Y(n_776)
);

INVxp67_ASAP7_75t_L g777 ( 
.A(n_776),
.Y(n_777)
);

AOI221xp5_ASAP7_75t_L g778 ( 
.A1(n_777),
.A2(n_611),
.B1(n_580),
.B2(n_595),
.C(n_598),
.Y(n_778)
);

AOI211xp5_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_589),
.B(n_603),
.C(n_595),
.Y(n_779)
);


endmodule