module fake_jpeg_12667_n_167 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_7),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_32),
.B(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_16),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_37),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_44),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_15),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_49),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_12),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_21),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_14),
.B1(n_20),
.B2(n_23),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_12),
.B(n_4),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_61),
.B(n_66),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_23),
.B(n_20),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_36),
.B(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_69),
.B(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_78),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_14),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_75),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_34),
.A2(n_29),
.B1(n_6),
.B2(n_10),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_50),
.B1(n_52),
.B2(n_46),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_40),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_58),
.C(n_60),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_89),
.Y(n_110)
);

BUFx16f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_93),
.Y(n_109)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_48),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_90),
.B(n_91),
.Y(n_123)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_100),
.Y(n_114)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_102),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_77),
.B1(n_84),
.B2(n_79),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_103),
.B1(n_107),
.B2(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_70),
.B1(n_82),
.B2(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_58),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_106),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_82),
.B1(n_64),
.B2(n_76),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_82),
.B1(n_70),
.B2(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_68),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_118),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_85),
.A2(n_76),
.B1(n_72),
.B2(n_63),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_103),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_72),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_75),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_122),
.B(n_93),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_86),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_94),
.C(n_99),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_129),
.C(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_115),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_92),
.C(n_106),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_134),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_104),
.C(n_96),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_110),
.B(n_119),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_129),
.A2(n_110),
.B(n_118),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_86),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_126),
.C(n_133),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_110),
.B1(n_124),
.B2(n_128),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_151),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_87),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_117),
.B1(n_113),
.B2(n_121),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_141),
.B(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_156),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_147),
.C(n_145),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_138),
.B(n_113),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_158),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_133),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_116),
.B1(n_152),
.B2(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_160),
.B1(n_157),
.B2(n_131),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.C(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_161),
.B(n_95),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_111),
.C(n_108),
.Y(n_166)
);

AOI221xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_108),
.B1(n_88),
.B2(n_107),
.C(n_75),
.Y(n_167)
);


endmodule