module fake_jpeg_22851_n_41 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_41);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

INVx1_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

HAxp5_ASAP7_75t_SL g22 ( 
.A(n_10),
.B(n_14),
.CON(n_22),
.SN(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_27),
.B(n_3),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_32),
.B1(n_6),
.B2(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_33),
.B(n_22),
.Y(n_34)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_34),
.B(n_36),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_28),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_35),
.B(n_11),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_9),
.C(n_15),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_16),
.B(n_17),
.Y(n_41)
);


endmodule