module fake_jpeg_3425_n_517 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_517);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_10),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g142 ( 
.A(n_57),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_58),
.B(n_62),
.Y(n_133)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_60),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_64),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_67),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_16),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_0),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_68),
.B(n_70),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_69),
.B(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_71),
.Y(n_201)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_72),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_29),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_73),
.B(n_75),
.Y(n_128)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_15),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_79),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_80),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_16),
.C(n_15),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_81),
.B(n_39),
.C(n_23),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_31),
.B(n_12),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_98),
.Y(n_136)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_86),
.Y(n_175)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_88),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_89),
.Y(n_180)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_96),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_97),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_1),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_11),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_100),
.B(n_101),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_21),
.B(n_12),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_26),
.B(n_1),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_103),
.B(n_120),
.Y(n_187)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_104),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_32),
.B(n_1),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_106),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_32),
.B(n_2),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_116),
.Y(n_162)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_43),
.Y(n_109)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_26),
.Y(n_110)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_28),
.Y(n_113)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_28),
.Y(n_114)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_43),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_117),
.B(n_119),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_20),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_121),
.Y(n_176)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_43),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_122),
.B(n_27),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_20),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_78),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_68),
.A2(n_54),
.B1(n_49),
.B2(n_20),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g236 ( 
.A1(n_138),
.A2(n_146),
.B1(n_150),
.B2(n_152),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_143),
.B(n_205),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_68),
.A2(n_54),
.B1(n_41),
.B2(n_38),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_68),
.A2(n_49),
.B1(n_41),
.B2(n_38),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_109),
.A2(n_39),
.B1(n_51),
.B2(n_50),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_151),
.A2(n_156),
.B1(n_166),
.B2(n_167),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_70),
.A2(n_95),
.B1(n_64),
.B2(n_84),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_122),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_154),
.B(n_164),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_64),
.A2(n_49),
.B1(n_38),
.B2(n_41),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_81),
.B(n_37),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_55),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_165),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_98),
.A2(n_37),
.B1(n_51),
.B2(n_50),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_79),
.A2(n_55),
.B1(n_53),
.B2(n_40),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_83),
.A2(n_46),
.B1(n_45),
.B2(n_23),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_170),
.A2(n_178),
.B1(n_146),
.B2(n_156),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_105),
.B(n_53),
.C(n_46),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_171),
.B(n_152),
.C(n_153),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_79),
.A2(n_45),
.B1(n_4),
.B2(n_5),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_172),
.A2(n_191),
.B1(n_204),
.B2(n_206),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_108),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_174),
.A2(n_177),
.B1(n_179),
.B2(n_184),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_88),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_93),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_63),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_71),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_96),
.B(n_72),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_186),
.B(n_192),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_80),
.A2(n_115),
.B1(n_114),
.B2(n_104),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_189),
.A2(n_193),
.B1(n_200),
.B2(n_203),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_84),
.A2(n_66),
.B1(n_60),
.B2(n_107),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_74),
.B(n_76),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_117),
.A2(n_90),
.B1(n_87),
.B2(n_96),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_92),
.B(n_57),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_195),
.B(n_199),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_59),
.B(n_92),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_77),
.A2(n_119),
.B1(n_85),
.B2(n_86),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_119),
.A2(n_91),
.B1(n_57),
.B2(n_97),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_91),
.A2(n_61),
.B1(n_89),
.B2(n_102),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_68),
.A2(n_47),
.B1(n_70),
.B2(n_30),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_58),
.B(n_62),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_197),
.Y(n_247)
);

OR2x2_ASAP7_75t_SL g211 ( 
.A(n_143),
.B(n_171),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_211),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_194),
.B1(n_157),
.B2(n_132),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_214),
.A2(n_222),
.B1(n_243),
.B2(n_248),
.Y(n_308)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_217),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_218),
.B(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_133),
.B(n_128),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_219),
.B(n_224),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_148),
.A2(n_158),
.B1(n_196),
.B2(n_135),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_220),
.A2(n_250),
.B1(n_276),
.B2(n_262),
.Y(n_324)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_132),
.A2(n_180),
.B1(n_209),
.B2(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_139),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_126),
.B(n_182),
.Y(n_224)
);

CKINVDCx12_ASAP7_75t_R g225 ( 
.A(n_142),
.Y(n_225)
);

INVx6_ASAP7_75t_SL g303 ( 
.A(n_225),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_226),
.A2(n_259),
.B1(n_266),
.B2(n_282),
.Y(n_286)
);

AO22x1_ASAP7_75t_SL g227 ( 
.A1(n_205),
.A2(n_139),
.B1(n_198),
.B2(n_150),
.Y(n_227)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_228),
.Y(n_334)
);

BUFx12_ASAP7_75t_L g229 ( 
.A(n_142),
.Y(n_229)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_229),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_176),
.Y(n_230)
);

NAND3xp33_ASAP7_75t_L g312 ( 
.A(n_230),
.B(n_244),
.C(n_247),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_162),
.B(n_124),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_234),
.Y(n_298)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_144),
.Y(n_232)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_232),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_233),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_131),
.B(n_145),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g235 ( 
.A1(n_206),
.A2(n_198),
.B1(n_209),
.B2(n_173),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_235),
.A2(n_278),
.B(n_283),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_141),
.B(n_163),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_237),
.B(n_241),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_125),
.B(n_130),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_239),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_130),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_168),
.Y(n_240)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_138),
.B(n_137),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_134),
.Y(n_242)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_242),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_180),
.A2(n_208),
.B1(n_188),
.B2(n_142),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_190),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_161),
.Y(n_245)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_201),
.Y(n_246)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_188),
.A2(n_208),
.B1(n_204),
.B2(n_160),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_127),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_249),
.B(n_255),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_201),
.A2(n_210),
.B1(n_129),
.B2(n_185),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_252),
.B(n_257),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_183),
.B(n_202),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_153),
.B(n_160),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_129),
.A2(n_185),
.B1(n_149),
.B2(n_191),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_258),
.A2(n_263),
.B(n_275),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_167),
.A2(n_172),
.B1(n_169),
.B2(n_149),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_127),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_261),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_160),
.B(n_140),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_159),
.A2(n_175),
.B1(n_140),
.B2(n_155),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_155),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_265),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_169),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_159),
.A2(n_150),
.B1(n_138),
.B2(n_146),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_176),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_272),
.Y(n_323)
);

BUFx12_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

CKINVDCx10_ASAP7_75t_R g284 ( 
.A(n_270),
.Y(n_284)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_142),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_271),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_176),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_273),
.Y(n_316)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_139),
.B(n_186),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_203),
.A2(n_193),
.B1(n_47),
.B2(n_96),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_163),
.Y(n_277)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_157),
.A2(n_164),
.B1(n_68),
.B2(n_162),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_144),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_279),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g280 ( 
.A1(n_139),
.A2(n_166),
.B(n_170),
.C(n_206),
.Y(n_280)
);

O2A1O1Ixp33_ASAP7_75t_L g320 ( 
.A1(n_280),
.A2(n_252),
.B(n_236),
.C(n_227),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_136),
.B(n_143),
.C(n_131),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g330 ( 
.A(n_281),
.B(n_278),
.CI(n_231),
.CON(n_330),
.SN(n_330)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_286),
.A2(n_299),
.B1(n_325),
.B2(n_331),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_266),
.A2(n_253),
.B1(n_241),
.B2(n_262),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_212),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g368 ( 
.A1(n_302),
.A2(n_304),
.B(n_317),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_215),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_234),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_245),
.Y(n_352)
);

AOI21xp33_ASAP7_75t_L g317 ( 
.A1(n_223),
.A2(n_215),
.B(n_275),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_218),
.B(n_215),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_329),
.Y(n_337)
);

BUFx24_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_275),
.A2(n_213),
.B(n_259),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_322),
.B(n_309),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_324),
.A2(n_314),
.B1(n_289),
.B2(n_322),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_253),
.A2(n_235),
.B1(n_280),
.B2(n_254),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_326),
.B(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_216),
.B(n_237),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_330),
.B(n_230),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_280),
.A2(n_216),
.B1(n_236),
.B2(n_258),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_236),
.A2(n_227),
.B1(n_269),
.B2(n_265),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_333),
.A2(n_335),
.B1(n_257),
.B2(n_244),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_236),
.A2(n_235),
.B1(n_242),
.B2(n_263),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_260),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_340),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_303),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_370),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_294),
.B(n_249),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_341),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_221),
.B1(n_273),
.B2(n_268),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_342),
.A2(n_358),
.B1(n_359),
.B2(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_306),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

OAI22x1_ASAP7_75t_L g398 ( 
.A1(n_346),
.A2(n_347),
.B1(n_293),
.B2(n_301),
.Y(n_398)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_295),
.Y(n_348)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_348),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_319),
.B(n_240),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_321),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_277),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_353),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_352),
.B(n_356),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_292),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_228),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_354),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_286),
.A2(n_217),
.B1(n_274),
.B2(n_256),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_357),
.B1(n_361),
.B2(n_300),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_298),
.B(n_257),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_233),
.B1(n_246),
.B2(n_267),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_325),
.A2(n_279),
.B1(n_232),
.B2(n_251),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_289),
.A2(n_271),
.B1(n_229),
.B2(n_270),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_297),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_326),
.A2(n_311),
.B1(n_328),
.B2(n_320),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_229),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_297),
.Y(n_363)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_304),
.A2(n_270),
.B1(n_302),
.B2(n_308),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_365),
.A2(n_372),
.B(n_321),
.Y(n_389)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_291),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_373),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_298),
.B(n_287),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_367),
.B(n_369),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_290),
.B(n_323),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_312),
.B(n_296),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_309),
.A2(n_305),
.B1(n_330),
.B2(n_332),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_371),
.A2(n_300),
.B1(n_334),
.B2(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_291),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_339),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_381),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g381 ( 
.A(n_361),
.B(n_330),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_332),
.B(n_313),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_382),
.A2(n_383),
.B(n_384),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_372),
.A2(n_313),
.B(n_284),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_336),
.A2(n_284),
.B1(n_327),
.B2(n_285),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_392),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g404 ( 
.A(n_389),
.B(n_395),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_338),
.B(n_306),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_340),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_365),
.A2(n_285),
.B(n_327),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_396),
.A2(n_397),
.B1(n_398),
.B2(n_355),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_346),
.A2(n_310),
.B1(n_295),
.B2(n_301),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_373),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_334),
.C(n_318),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_359),
.C(n_364),
.Y(n_410)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_393),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_403),
.B(n_407),
.Y(n_441)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_396),
.A2(n_374),
.B1(n_398),
.B2(n_342),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_406),
.A2(n_414),
.B1(n_399),
.B2(n_357),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_377),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_408),
.B(n_423),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_400),
.C(n_384),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_344),
.C(n_350),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_424),
.C(n_389),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_379),
.B(n_353),
.Y(n_412)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_412),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_383),
.A2(n_349),
.B(n_368),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_413),
.A2(n_381),
.B(n_349),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_374),
.A2(n_371),
.B1(n_397),
.B2(n_379),
.Y(n_414)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_418),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_395),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_337),
.Y(n_419)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_422),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_375),
.B(n_369),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_421),
.B(n_425),
.Y(n_448)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_337),
.C(n_351),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_376),
.B(n_367),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_391),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_378),
.B(n_360),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_385),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_409),
.A2(n_378),
.B1(n_358),
.B2(n_349),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_429),
.A2(n_440),
.B(n_417),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_434),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_421),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_439),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_435),
.A2(n_445),
.B1(n_403),
.B2(n_402),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_415),
.B(n_382),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_437),
.B(n_413),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_426),
.Y(n_439)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_442),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_401),
.Y(n_443)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_443),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_349),
.B1(n_385),
.B2(n_401),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_426),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_446),
.B(n_345),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_448),
.B(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_461),
.Y(n_470)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_450),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_415),
.C(n_410),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_458),
.C(n_462),
.Y(n_468)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_455),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_467),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_424),
.C(n_411),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_409),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_460),
.B(n_458),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_427),
.C(n_418),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_412),
.C(n_419),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_444),
.C(n_428),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_464),
.A2(n_404),
.B(n_431),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_448),
.B(n_407),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_465),
.B(n_432),
.Y(n_469)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_SL g481 ( 
.A1(n_466),
.A2(n_416),
.B1(n_446),
.B2(n_439),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_444),
.A2(n_404),
.B(n_417),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_469),
.A2(n_481),
.B1(n_455),
.B2(n_467),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_471),
.B(n_472),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_428),
.C(n_440),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_445),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_477),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_475),
.A2(n_443),
.B(n_433),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_451),
.B(n_442),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_478),
.B(n_433),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_470),
.B(n_461),
.Y(n_482)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_482),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_447),
.Y(n_483)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_431),
.B1(n_450),
.B2(n_452),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_486),
.B1(n_487),
.B2(n_438),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_476),
.A2(n_435),
.B1(n_464),
.B2(n_436),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_479),
.A2(n_436),
.B1(n_438),
.B2(n_453),
.Y(n_487)
);

AO21x1_ASAP7_75t_L g488 ( 
.A1(n_475),
.A2(n_460),
.B(n_429),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_488),
.A2(n_492),
.B(n_472),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_490),
.A2(n_491),
.B1(n_471),
.B2(n_474),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_484),
.B(n_416),
.Y(n_493)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_493),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_473),
.Y(n_494)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_499),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_489),
.B(n_477),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_495),
.B(n_496),
.Y(n_507)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_501),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_499),
.B(n_468),
.C(n_454),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_504),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_468),
.C(n_456),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_505),
.A2(n_498),
.B(n_497),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_509),
.B(n_510),
.C(n_511),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_488),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_496),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_502),
.C(n_505),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_511),
.B(n_497),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_514),
.A2(n_515),
.B(n_492),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_512),
.B(n_501),
.C(n_485),
.Y(n_515)
);

FAx1_ASAP7_75t_SL g517 ( 
.A(n_516),
.B(n_462),
.CI(n_487),
.CON(n_517),
.SN(n_517)
);


endmodule